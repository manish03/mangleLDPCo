//`include "GF2_LDPC_fgallag_0x00005_assign_inc.sv"
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00000] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00000] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00001] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00001] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00002] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00003] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00002] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00004] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00005] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00003] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00006] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00007] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00004] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00008] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00009] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00005] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0000a] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0000b] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00006] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0000c] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0000d] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00007] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0000e] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0000f] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00008] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00010] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00011] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00009] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00012] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00013] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0000a] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00014] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00015] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0000b] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00016] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00017] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0000c] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00018] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00019] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0000d] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0001a] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0001b] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0000e] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0001c] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0001d] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0000f] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0001e] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0001f] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00010] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00020] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00021] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00011] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00022] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00023] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00012] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00024] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00025] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00013] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00026] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00027] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00014] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00028] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00029] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00015] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0002a] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0002b] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00016] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0002c] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0002d] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00017] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0002e] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0002f] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00018] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00030] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00031] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00019] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00032] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00033] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0001a] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00034] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00035] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0001b] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00036] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00037] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0001c] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00038] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00039] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0001d] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0003a] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0003b] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0001e] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0003c] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0003d] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0001f] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0003e] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0003f] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00020] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00040] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00041] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00021] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00042] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00043] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00022] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00044] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00045] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00023] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00046] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00047] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00024] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00048] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00049] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00025] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0004a] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0004b] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00026] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0004c] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0004d] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00027] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0004e] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0004f] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00028] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00050] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00051] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00029] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00052] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00053] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0002a] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00054] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00055] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0002b] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00056] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00057] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0002c] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00058] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00059] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0002d] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0005a] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0005b] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0002e] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0005c] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0005d] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0002f] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0005e] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0005f] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00030] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00060] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00061] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00031] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00062] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00063] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00032] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00064] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00065] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00033] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00066] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00067] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00034] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00068] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00069] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00035] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0006a] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0006b] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00036] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0006c] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0006d] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00037] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0006e] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0006f] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00038] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00070] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00071] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00039] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00072] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00073] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0003a] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00074] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00075] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0003b] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00076] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00077] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0003c] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00078] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00079] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0003d] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0007a] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0007b] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0003e] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0007c] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0007d] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0003f] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0007e] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0007f] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00040] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00080] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00081] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00041] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00082] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00083] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00042] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00084] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00085] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00043] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00086] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00087] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00044] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00088] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00089] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00045] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0008a] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0008b] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00046] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0008c] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0008d] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00047] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0008e] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0008f] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00048] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00090] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00091] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00049] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00092] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00093] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0004a] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00094] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00095] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0004b] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00096] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00097] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0004c] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00098] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00099] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0004d] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0009a] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0009b] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0004e] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0009c] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0009d] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0004f] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0009e] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0009f] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00050] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000a0] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000a1] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00051] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000a2] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000a3] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00052] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000a4] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000a5] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00053] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000a6] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000a7] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00054] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000a8] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000a9] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00055] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000aa] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000ab] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00056] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000ac] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000ad] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00057] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000ae] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000af] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00058] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000b0] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000b1] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00059] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000b2] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000b3] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0005a] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000b4] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000b5] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0005b] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000b6] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000b7] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0005c] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000b8] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000b9] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0005d] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000ba] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000bb] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0005e] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000bc] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000bd] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0005f] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000be] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000bf] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00060] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000c0] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000c1] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00061] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000c2] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000c3] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00062] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000c4] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000c5] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00063] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000c6] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000c7] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00064] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000c8] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000c9] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00065] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000ca] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000cb] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00066] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000cc] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000cd] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00067] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000ce] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000cf] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00068] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000d0] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000d1] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00069] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000d2] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000d3] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0006a] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000d4] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000d5] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0006b] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000d6] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000d7] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0006c] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000d8] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000d9] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0006d] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000da] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000db] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0006e] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000dc] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000dd] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0006f] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000de] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000df] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00070] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000e0] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000e1] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00071] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000e2] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000e3] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00072] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000e4] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000e5] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00073] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000e6] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000e7] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00074] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000e8] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000e9] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00075] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000ea] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000eb] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00076] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000ec] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000ed] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00077] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000ee] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000ef] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00078] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000f0] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000f1] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00079] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000f2] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000f3] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0007a] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000f4] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000f5] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0007b] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000f6] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000f7] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0007c] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000f8] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000f9] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0007d] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000fa] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000fb] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0007e] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000fc] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000fd] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0007f] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000fe] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h000ff] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00080] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00100] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00101] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00081] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00102] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00103] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00082] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00104] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00105] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00083] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00106] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00107] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00084] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00108] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00109] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00085] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0010a] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0010b] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00086] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0010c] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0010d] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00087] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0010e] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0010f] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00088] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00110] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00111] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00089] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00112] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00113] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0008a] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00114] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00115] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0008b] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00116] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00117] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0008c] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00118] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00119] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0008d] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0011a] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0011b] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0008e] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0011c] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0011d] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0008f] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0011e] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0011f] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00090] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00120] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00121] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00091] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00122] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00123] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00092] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00124] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00125] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00093] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00126] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00127] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00094] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00128] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00129] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00095] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0012a] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0012b] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00096] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0012c] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0012d] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00097] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0012e] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0012f] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00098] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00130] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00131] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00099] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00132] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00133] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0009a] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00134] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00135] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0009b] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00136] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00137] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0009c] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00138] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00139] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0009d] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0013a] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0013b] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0009e] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0013c] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0013d] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0009f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0013e] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000a0] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00140] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00141] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000a1] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00142] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00143] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000a2] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00144] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00145] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000a3] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00146] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00147] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000a4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00148] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000a5] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0014a] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0014b] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000a6] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0014c] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0014d] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000a7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0014e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000a8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00150] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000a9] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00152] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00153] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000aa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00154] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000ab] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00156] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00157] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000ac] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00158] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00159] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000ad] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0015a] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000ae] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0015c] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0015d] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000af] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0015e] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000b0] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00160] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00161] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000b1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00162] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000b2] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00164] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00165] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000b3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00166] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000b4] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00168] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00169] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000b5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0016a] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000b6] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0016c] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0016d] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000b7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0016e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000b8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00170] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000b9] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00172] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00173] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000ba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00174] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000bb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00176] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000bc] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00178] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00179] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000bd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0017a] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000be] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0017c] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0017d] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000bf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0017e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000c0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00180] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000c1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00182] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000c2] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00184] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00185] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000c3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00186] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000c4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00188] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000c5] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0018a] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0018b] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000c6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0018c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000c7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0018e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000c8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00190] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000c9] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00192] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00193] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000ca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00194] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000cb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00196] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000cc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00198] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000cd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0019a] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000ce] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0019c] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0019d] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000cf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0019e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000d0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000d1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000d2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001a4] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000d3] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001a6] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001a7] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000d4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000d5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000d6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000d7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000d8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000d9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001b2] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000da] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001b4] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001b5] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000db] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000dc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000dd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000de] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000df] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000e0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000e1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001c2] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000e2] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001c4] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001c5] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000e3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000e4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000e5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000e6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000e7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000e8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000e9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000ea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000eb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001d6] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000ec] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001d8] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001d9] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000ed] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000ee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000ef] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000f0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000f1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000f2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000f3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000f4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000f5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000f6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000f7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000f8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000f9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000fa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000fb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000fc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001f8] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000fd] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001fa] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001fb] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000fe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000ff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h001fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00100] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00200] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00101] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00202] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00102] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00204] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00103] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00206] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00104] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00208] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00105] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0020a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00106] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0020c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00107] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0020e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00108] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00210] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00109] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00212] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0010a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00214] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0010b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00216] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0010c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00218] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0010d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0021a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0010e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0021c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0010f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0021e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00110] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00220] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00111] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00222] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00112] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00224] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00113] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00226] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00114] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00228] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00115] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0022a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00116] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0022c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00117] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0022e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00118] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00230] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00119] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00232] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0011a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00234] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0011b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00236] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0011c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00238] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0011d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0023a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0011e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0023c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0011f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0023e] ;
//end
//always_comb begin
              Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00120] = 
          (!fgallag_sel['h00005]) ? 
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00240] : //%
                       Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00241] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00121] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00242] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00122] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00244] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00123] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00246] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00124] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00248] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00125] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0024a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00126] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0024c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00127] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0024e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00128] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00250] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00129] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00252] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0012a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00254] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0012b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00256] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0012c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00258] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0012d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0025a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0012e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0025c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0012f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0025e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00130] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00260] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00131] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00262] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00132] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00264] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00133] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00266] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00134] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00268] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00135] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0026a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00136] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0026c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00137] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0026e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00138] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00270] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00139] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00272] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0013a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00274] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0013b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00276] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0013c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00278] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0013d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0027a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0013e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0027c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0013f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0027e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00140] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00280] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00141] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00282] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00142] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00284] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00143] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00286] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00144] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00288] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00145] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0028a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00146] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0028c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00147] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0028e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00148] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00290] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00149] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00292] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0014a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00294] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0014b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00296] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0014c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00298] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0014d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0029a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0014e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0029c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0014f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0029e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00150] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00151] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00152] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00153] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00154] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00155] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00156] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00157] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00158] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00159] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0015a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0015b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0015c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0015d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0015e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0015f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00160] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00161] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00162] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00163] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00164] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00165] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00166] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00167] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00168] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00169] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0016a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0016b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0016c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0016d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0016e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0016f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00170] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00171] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00172] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00173] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00174] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00175] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00176] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00177] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00178] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00179] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0017a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0017b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0017c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0017d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0017e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0017f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h002fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00180] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00300] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00181] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00302] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00182] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00304] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00183] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00306] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00184] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00308] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00185] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0030a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00186] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0030c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00187] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0030e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00188] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00310] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00189] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00312] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0018a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00314] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0018b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00316] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0018c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00318] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0018d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0031a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0018e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0031c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0018f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0031e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00190] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00320] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00191] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00322] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00192] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00324] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00193] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00326] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00194] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00328] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00195] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0032a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00196] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0032c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00197] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0032e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00198] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00330] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00199] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00332] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0019a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00334] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0019b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00336] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0019c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00338] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0019d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0033a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0019e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0033c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0019f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0033e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001a0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00340] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001a1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00342] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001a2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00344] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001a3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00346] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001a4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00348] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001a5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0034a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001a6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0034c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001a7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0034e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001a8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00350] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001a9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00352] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001aa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00354] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001ab] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00356] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001ac] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00358] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001ad] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0035a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001ae] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0035c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001af] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0035e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001b0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00360] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001b1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00362] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001b2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00364] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001b3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00366] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001b4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00368] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001b5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0036a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001b6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0036c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001b7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0036e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001b8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00370] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001b9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00372] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001ba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00374] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001bb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00376] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001bc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00378] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001bd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0037a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001be] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0037c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001bf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0037e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001c0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00380] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001c1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00382] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001c2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00384] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001c3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00386] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001c4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00388] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001c5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0038a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001c6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0038c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001c7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0038e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001c8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00390] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001c9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00392] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001ca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00394] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001cb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00396] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001cc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00398] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001cd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0039a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001ce] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0039c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001cf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0039e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001d0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001d1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001d2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001d3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001d4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001d5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001d6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001d7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001d8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001d9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001da] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001db] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001dc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001dd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001de] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001df] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001e0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001e1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001e2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001e3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001e4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001e5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001e6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001e7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001e8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001e9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001ea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001eb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001ec] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001ed] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001ee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001ef] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001f0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001f1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001f2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001f3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001f4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001f5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001f6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001f7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001f8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001f9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001fa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001fb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001fc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001fd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001fe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001ff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h003fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00200] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00400] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00201] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00402] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00202] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00404] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00203] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00406] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00204] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00408] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00205] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0040a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00206] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0040c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00207] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0040e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00208] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00410] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00209] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00412] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0020a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00414] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0020b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00416] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0020c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00418] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0020d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0041a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0020e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0041c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0020f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0041e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00210] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00420] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00211] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00422] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00212] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00424] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00213] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00426] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00214] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00428] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00215] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0042a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00216] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0042c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00217] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0042e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00218] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00430] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00219] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00432] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0021a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00434] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0021b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00436] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0021c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00438] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0021d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0043a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0021e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0043c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0021f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0043e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00220] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00440] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00221] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00442] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00222] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00444] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00223] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00446] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00224] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00448] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00225] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0044a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00226] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0044c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00227] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0044e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00228] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00450] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00229] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00452] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0022a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00454] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0022b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00456] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0022c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00458] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0022d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0045a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0022e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0045c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0022f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0045e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00230] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00460] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00231] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00462] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00232] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00464] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00233] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00466] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00234] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00468] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00235] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0046a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00236] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0046c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00237] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0046e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00238] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00470] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00239] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00472] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0023a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00474] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0023b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00476] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0023c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00478] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0023d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0047a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0023e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0047c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0023f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0047e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00240] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00480] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00241] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00482] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00242] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00484] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00243] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00486] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00244] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00488] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00245] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0048a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00246] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0048c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00247] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0048e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00248] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00490] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00249] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00492] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0024a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00494] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0024b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00496] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0024c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00498] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0024d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0049a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0024e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0049c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0024f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0049e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00250] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00251] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00252] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00253] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00254] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00255] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00256] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00257] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00258] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00259] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0025a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0025b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0025c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0025d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0025e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0025f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00260] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00261] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00262] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00263] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00264] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00265] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00266] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00267] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00268] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00269] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0026a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0026b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0026c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0026d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0026e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0026f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00270] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00271] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00272] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00273] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00274] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00275] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00276] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00277] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00278] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00279] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0027a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0027b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0027c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0027d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0027e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0027f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h004fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00280] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00500] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00281] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00502] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00282] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00504] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00283] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00506] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00284] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00508] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00285] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0050a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00286] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0050c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00287] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0050e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00288] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00510] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00289] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00512] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0028a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00514] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0028b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00516] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0028c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00518] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0028d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0051a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0028e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0051c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0028f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0051e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00290] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00520] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00291] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00522] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00292] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00524] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00293] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00526] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00294] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00528] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00295] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0052a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00296] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0052c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00297] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0052e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00298] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00530] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00299] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00532] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0029a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00534] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0029b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00536] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0029c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00538] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0029d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0053a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0029e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0053c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0029f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0053e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002a0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00540] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002a1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00542] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002a2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00544] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002a3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00546] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002a4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00548] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002a5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0054a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002a6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0054c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002a7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0054e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002a8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00550] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002a9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00552] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002aa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00554] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002ab] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00556] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002ac] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00558] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002ad] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0055a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002ae] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0055c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002af] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0055e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002b0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00560] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002b1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00562] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002b2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00564] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002b3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00566] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002b4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00568] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002b5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0056a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002b6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0056c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002b7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0056e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002b8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00570] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002b9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00572] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002ba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00574] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002bb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00576] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002bc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00578] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002bd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0057a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002be] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0057c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002bf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0057e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002c0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00580] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002c1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00582] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002c2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00584] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002c3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00586] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002c4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00588] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002c5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0058a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002c6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0058c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002c7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0058e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002c8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00590] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002c9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00592] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002ca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00594] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002cb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00596] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002cc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00598] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002cd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0059a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002ce] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0059c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002cf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0059e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002d0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002d1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002d2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002d3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002d4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002d5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002d6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002d7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002d8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002d9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002da] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002db] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002dc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002dd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002de] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002df] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002e0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002e1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002e2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002e3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002e4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002e5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002e6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002e7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002e8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002e9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002ea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002eb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002ec] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002ed] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002ee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002ef] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002f0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002f1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002f2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002f3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002f4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002f5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002f6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002f7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002f8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002f9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002fa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002fb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002fc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002fd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002fe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002ff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h005fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00300] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00600] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00301] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00602] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00302] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00604] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00303] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00606] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00304] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00608] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00305] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0060a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00306] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0060c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00307] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0060e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00308] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00610] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00309] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00612] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0030a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00614] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0030b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00616] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0030c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00618] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0030d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0061a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0030e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0061c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0030f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0061e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00310] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00620] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00311] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00622] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00312] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00624] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00313] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00626] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00314] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00628] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00315] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0062a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00316] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0062c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00317] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0062e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00318] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00630] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00319] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00632] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0031a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00634] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0031b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00636] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0031c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00638] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0031d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0063a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0031e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0063c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0031f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0063e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00320] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00640] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00321] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00642] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00322] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00644] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00323] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00646] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00324] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00648] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00325] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0064a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00326] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0064c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00327] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0064e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00328] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00650] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00329] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00652] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0032a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00654] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0032b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00656] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0032c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00658] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0032d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0065a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0032e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0065c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0032f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0065e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00330] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00660] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00331] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00662] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00332] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00664] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00333] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00666] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00334] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00668] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00335] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0066a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00336] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0066c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00337] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0066e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00338] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00670] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00339] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00672] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0033a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00674] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0033b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00676] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0033c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00678] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0033d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0067a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0033e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0067c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0033f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0067e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00340] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00680] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00341] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00682] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00342] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00684] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00343] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00686] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00344] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00688] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00345] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0068a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00346] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0068c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00347] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0068e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00348] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00690] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00349] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00692] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0034a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00694] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0034b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00696] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0034c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00698] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0034d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0069a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0034e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0069c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0034f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0069e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00350] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00351] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00352] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00353] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00354] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00355] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00356] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00357] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00358] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00359] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0035a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0035b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0035c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0035d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0035e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0035f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00360] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00361] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00362] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00363] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00364] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00365] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00366] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00367] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00368] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00369] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0036a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0036b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0036c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0036d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0036e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0036f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00370] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00371] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00372] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00373] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00374] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00375] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00376] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00377] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00378] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00379] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0037a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0037b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0037c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0037d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0037e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0037f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h006fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00380] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00700] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00381] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00702] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00382] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00704] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00383] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00706] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00384] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00708] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00385] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0070a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00386] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0070c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00387] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0070e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00388] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00710] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00389] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00712] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0038a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00714] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0038b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00716] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0038c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00718] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0038d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0071a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0038e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0071c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0038f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0071e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00390] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00720] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00391] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00722] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00392] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00724] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00393] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00726] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00394] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00728] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00395] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0072a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00396] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0072c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00397] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0072e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00398] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00730] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00399] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00732] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0039a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00734] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0039b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00736] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0039c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00738] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0039d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0073a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0039e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0073c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0039f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0073e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003a0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00740] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003a1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00742] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003a2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00744] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003a3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00746] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003a4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00748] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003a5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0074a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003a6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0074c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003a7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0074e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003a8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00750] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003a9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00752] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003aa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00754] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003ab] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00756] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003ac] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00758] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003ad] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0075a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003ae] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0075c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003af] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0075e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003b0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00760] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003b1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00762] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003b2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00764] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003b3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00766] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003b4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00768] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003b5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0076a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003b6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0076c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003b7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0076e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003b8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00770] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003b9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00772] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003ba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00774] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003bb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00776] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003bc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00778] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003bd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0077a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003be] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0077c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003bf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0077e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003c0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00780] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003c1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00782] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003c2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00784] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003c3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00786] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003c4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00788] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003c5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0078a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003c6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0078c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003c7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0078e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003c8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00790] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003c9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00792] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003ca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00794] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003cb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00796] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003cc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00798] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003cd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0079a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003ce] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0079c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003cf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0079e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003d0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003d1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003d2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003d3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003d4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003d5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003d6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003d7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003d8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003d9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003da] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003db] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003dc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003dd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003de] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003df] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003e0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003e1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003e2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003e3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003e4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003e5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003e6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003e7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003e8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003e9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003ea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003eb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003ec] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003ed] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003ee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003ef] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003f0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003f1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003f2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003f3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003f4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003f5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003f6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003f7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003f8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003f9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003fa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003fb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003fc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003fd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003fe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003ff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h007fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00400] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00800] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00401] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00802] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00402] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00804] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00403] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00806] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00404] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00808] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00405] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0080a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00406] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0080c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00407] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0080e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00408] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00810] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00409] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00812] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0040a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00814] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0040b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00816] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0040c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00818] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0040d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0081a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0040e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0081c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0040f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0081e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00410] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00820] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00411] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00822] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00412] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00824] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00413] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00826] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00414] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00828] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00415] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0082a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00416] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0082c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00417] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0082e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00418] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00830] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00419] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00832] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0041a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00834] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0041b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00836] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0041c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00838] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0041d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0083a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0041e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0083c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0041f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0083e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00420] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00840] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00421] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00842] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00422] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00844] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00423] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00846] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00424] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00848] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00425] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0084a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00426] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0084c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00427] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0084e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00428] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00850] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00429] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00852] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0042a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00854] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0042b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00856] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0042c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00858] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0042d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0085a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0042e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0085c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0042f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0085e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00430] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00860] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00431] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00862] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00432] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00864] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00433] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00866] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00434] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00868] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00435] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0086a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00436] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0086c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00437] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0086e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00438] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00870] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00439] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00872] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0043a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00874] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0043b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00876] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0043c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00878] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0043d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0087a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0043e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0087c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0043f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0087e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00440] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00880] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00441] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00882] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00442] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00884] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00443] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00886] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00444] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00888] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00445] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0088a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00446] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0088c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00447] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0088e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00448] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00890] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00449] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00892] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0044a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00894] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0044b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00896] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0044c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00898] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0044d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0089a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0044e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0089c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0044f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0089e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00450] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00451] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00452] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00453] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00454] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00455] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00456] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00457] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00458] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00459] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0045a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0045b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0045c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0045d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0045e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0045f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00460] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00461] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00462] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00463] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00464] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00465] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00466] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00467] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00468] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00469] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0046a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0046b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0046c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0046d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0046e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0046f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00470] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00471] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00472] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00473] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00474] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00475] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00476] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00477] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00478] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00479] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0047a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0047b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0047c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0047d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0047e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0047f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h008fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00480] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00900] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00481] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00902] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00482] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00904] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00483] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00906] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00484] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00908] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00485] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0090a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00486] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0090c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00487] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0090e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00488] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00910] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00489] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00912] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0048a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00914] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0048b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00916] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0048c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00918] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0048d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0091a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0048e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0091c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0048f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0091e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00490] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00920] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00491] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00922] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00492] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00924] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00493] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00926] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00494] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00928] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00495] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0092a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00496] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0092c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00497] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0092e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00498] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00930] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00499] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00932] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0049a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00934] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0049b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00936] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0049c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00938] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0049d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0093a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0049e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0093c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0049f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0093e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004a0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00940] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004a1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00942] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004a2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00944] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004a3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00946] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004a4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00948] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004a5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0094a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004a6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0094c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004a7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0094e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004a8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00950] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004a9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00952] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004aa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00954] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004ab] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00956] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004ac] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00958] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004ad] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0095a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004ae] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0095c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004af] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0095e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004b0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00960] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004b1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00962] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004b2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00964] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004b3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00966] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004b4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00968] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004b5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0096a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004b6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0096c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004b7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0096e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004b8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00970] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004b9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00972] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004ba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00974] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004bb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00976] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004bc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00978] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004bd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0097a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004be] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0097c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004bf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0097e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004c0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00980] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004c1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00982] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004c2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00984] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004c3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00986] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004c4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00988] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004c5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0098a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004c6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0098c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004c7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0098e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004c8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00990] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004c9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00992] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004ca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00994] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004cb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00996] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004cc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00998] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004cd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0099a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004ce] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0099c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004cf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0099e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004d0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004d1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004d2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004d3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004d4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004d5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004d6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004d7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004d8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004d9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004da] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004db] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004dc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004dd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004de] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004df] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004e0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004e1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004e2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004e3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004e4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004e5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004e6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004e7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004e8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004e9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004ea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004eb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004ec] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004ed] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004ee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004ef] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004f0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004f1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004f2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004f3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004f4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004f5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004f6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004f7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004f8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004f9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004fa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004fb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004fc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004fd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004fe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004ff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h009fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00500] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a00] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00501] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a02] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00502] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a04] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00503] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a06] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00504] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a08] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00505] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a0a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00506] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a0c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00507] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a0e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00508] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a10] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00509] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a12] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0050a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a14] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0050b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a16] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0050c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a18] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0050d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a1a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0050e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a1c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0050f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a1e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00510] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a20] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00511] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a22] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00512] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a24] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00513] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a26] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00514] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a28] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00515] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a2a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00516] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a2c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00517] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a2e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00518] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a30] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00519] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a32] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0051a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a34] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0051b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a36] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0051c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a38] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0051d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a3a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0051e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a3c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0051f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a3e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00520] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a40] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00521] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a42] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00522] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a44] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00523] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a46] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00524] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a48] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00525] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a4a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00526] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a4c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00527] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a4e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00528] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a50] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00529] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a52] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0052a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a54] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0052b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a56] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0052c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a58] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0052d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a5a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0052e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a5c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0052f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a5e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00530] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a60] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00531] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a62] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00532] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a64] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00533] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a66] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00534] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a68] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00535] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a6a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00536] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a6c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00537] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a6e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00538] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a70] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00539] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a72] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0053a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a74] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0053b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a76] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0053c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a78] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0053d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a7a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0053e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a7c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0053f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a7e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00540] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a80] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00541] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a82] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00542] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a84] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00543] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a86] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00544] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a88] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00545] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a8a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00546] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a8c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00547] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a8e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00548] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a90] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00549] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a92] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0054a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a94] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0054b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a96] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0054c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a98] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0054d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a9a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0054e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a9c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0054f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00a9e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00550] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aa0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00551] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aa2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00552] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aa4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00553] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aa6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00554] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aa8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00555] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aaa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00556] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00557] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00558] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ab0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00559] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ab2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0055a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ab4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0055b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ab6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0055c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ab8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0055d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0055e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00abc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0055f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00abe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00560] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ac0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00561] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ac2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00562] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ac4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00563] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ac6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00564] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ac8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00565] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00566] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00acc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00567] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ace] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00568] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ad0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00569] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ad2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0056a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ad4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0056b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ad6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0056c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ad8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0056d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ada] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0056e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00adc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0056f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ade] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00570] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ae0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00571] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ae2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00572] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ae4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00573] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ae6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00574] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ae8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00575] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00576] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00577] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00aee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00578] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00af0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00579] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00af2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0057a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00af4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0057b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00af6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0057c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00af8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0057d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00afa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0057e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00afc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0057f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00afe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00580] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b00] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00581] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b02] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00582] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b04] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00583] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b06] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00584] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b08] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00585] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b0a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00586] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b0c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00587] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b0e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00588] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b10] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00589] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b12] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0058a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b14] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0058b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b16] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0058c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b18] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0058d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b1a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0058e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b1c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0058f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b1e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00590] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b20] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00591] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b22] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00592] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b24] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00593] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b26] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00594] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b28] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00595] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b2a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00596] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b2c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00597] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b2e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00598] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b30] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00599] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b32] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0059a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b34] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0059b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b36] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0059c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b38] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0059d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b3a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0059e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b3c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0059f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b3e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005a0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b40] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005a1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b42] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005a2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b44] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005a3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b46] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005a4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b48] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005a5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b4a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005a6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b4c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005a7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b4e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005a8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b50] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005a9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b52] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005aa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b54] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005ab] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b56] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005ac] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b58] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005ad] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b5a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005ae] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b5c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005af] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b5e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005b0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b60] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005b1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b62] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005b2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b64] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005b3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b66] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005b4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b68] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005b5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b6a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005b6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b6c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005b7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b6e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005b8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b70] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005b9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b72] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005ba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b74] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005bb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b76] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005bc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b78] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005bd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b7a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005be] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b7c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005bf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b7e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005c0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b80] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005c1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b82] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005c2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b84] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005c3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b86] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005c4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b88] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005c5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b8a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005c6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b8c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005c7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b8e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005c8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b90] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005c9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b92] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005ca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b94] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005cb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b96] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005cc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b98] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005cd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b9a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005ce] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b9c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005cf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00b9e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005d0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ba0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005d1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ba2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005d2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ba4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005d3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ba6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005d4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ba8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005d5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00baa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005d6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005d7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005d8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bb0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005d9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bb2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005da] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bb4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005db] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bb6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005dc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bb8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005dd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005de] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bbc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005df] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bbe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005e0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bc0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005e1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bc2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005e2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bc4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005e3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bc6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005e4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bc8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005e5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005e6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bcc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005e7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005e8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bd0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005e9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bd2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005ea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bd4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005eb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bd6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005ec] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bd8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005ed] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bda] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005ee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bdc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005ef] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bde] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005f0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00be0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005f1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00be2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005f2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00be4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005f3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00be6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005f4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00be8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005f5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005f6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005f7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005f8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bf0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005f9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bf2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005fa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bf4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005fb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bf6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005fc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bf8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005fd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bfa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005fe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bfc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005ff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00bfe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00600] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c00] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00601] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c02] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00602] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c04] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00603] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c06] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00604] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c08] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00605] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c0a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00606] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c0c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00607] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c0e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00608] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c10] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00609] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c12] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0060a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c14] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0060b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c16] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0060c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c18] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0060d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c1a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0060e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c1c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0060f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c1e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00610] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c20] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00611] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c22] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00612] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c24] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00613] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c26] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00614] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c28] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00615] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c2a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00616] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c2c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00617] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c2e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00618] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c30] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00619] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c32] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0061a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c34] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0061b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c36] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0061c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c38] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0061d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c3a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0061e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c3c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0061f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c3e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00620] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c40] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00621] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c42] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00622] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c44] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00623] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c46] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00624] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c48] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00625] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c4a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00626] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c4c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00627] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c4e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00628] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c50] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00629] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c52] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0062a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c54] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0062b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c56] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0062c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c58] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0062d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c5a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0062e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c5c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0062f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c5e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00630] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c60] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00631] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c62] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00632] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c64] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00633] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c66] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00634] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c68] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00635] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c6a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00636] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c6c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00637] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c6e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00638] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c70] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00639] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c72] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0063a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c74] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0063b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c76] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0063c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c78] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0063d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c7a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0063e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c7c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0063f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c7e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00640] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c80] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00641] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c82] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00642] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c84] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00643] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c86] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00644] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c88] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00645] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c8a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00646] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c8c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00647] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c8e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00648] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c90] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00649] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c92] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0064a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c94] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0064b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c96] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0064c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c98] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0064d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c9a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0064e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c9c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0064f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00c9e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00650] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ca0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00651] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ca2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00652] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ca4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00653] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ca6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00654] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ca8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00655] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00caa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00656] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00657] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00658] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cb0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00659] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cb2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0065a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cb4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0065b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cb6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0065c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cb8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0065d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0065e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cbc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0065f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cbe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00660] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cc0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00661] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cc2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00662] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cc4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00663] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cc6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00664] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cc8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00665] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00666] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ccc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00667] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00668] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cd0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00669] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cd2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0066a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cd4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0066b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cd6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0066c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cd8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0066d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cda] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0066e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cdc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0066f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cde] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00670] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ce0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00671] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ce2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00672] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ce4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00673] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ce6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00674] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ce8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00675] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00676] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00677] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00678] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cf0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00679] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cf2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0067a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cf4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0067b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cf6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0067c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cf8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0067d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cfa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0067e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cfc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0067f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00cfe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00680] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d00] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00681] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d02] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00682] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d04] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00683] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d06] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00684] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d08] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00685] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d0a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00686] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d0c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00687] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d0e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00688] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d10] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00689] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d12] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0068a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d14] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0068b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d16] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0068c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d18] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0068d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d1a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0068e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d1c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0068f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d1e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00690] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d20] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00691] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d22] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00692] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d24] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00693] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d26] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00694] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d28] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00695] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d2a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00696] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d2c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00697] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d2e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00698] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d30] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00699] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d32] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0069a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d34] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0069b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d36] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0069c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d38] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0069d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d3a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0069e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d3c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0069f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d3e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006a0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d40] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006a1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d42] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006a2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d44] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006a3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d46] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006a4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d48] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006a5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d4a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006a6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d4c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006a7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d4e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006a8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d50] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006a9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d52] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006aa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d54] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006ab] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d56] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006ac] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d58] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006ad] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d5a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006ae] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d5c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006af] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d5e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006b0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d60] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006b1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d62] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006b2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d64] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006b3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d66] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006b4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d68] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006b5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d6a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006b6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d6c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006b7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d6e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006b8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d70] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006b9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d72] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006ba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d74] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006bb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d76] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006bc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d78] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006bd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d7a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006be] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d7c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006bf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d7e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006c0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d80] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006c1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d82] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006c2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d84] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006c3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d86] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006c4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d88] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006c5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d8a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006c6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d8c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006c7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d8e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006c8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d90] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006c9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d92] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006ca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d94] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006cb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d96] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006cc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d98] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006cd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d9a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006ce] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d9c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006cf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00d9e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006d0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00da0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006d1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00da2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006d2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00da4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006d3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00da6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006d4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00da8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006d5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00daa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006d6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006d7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006d8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00db0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006d9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00db2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006da] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00db4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006db] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00db6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006dc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00db8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006dd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006de] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dbc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006df] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dbe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006e0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dc0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006e1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dc2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006e2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dc4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006e3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dc6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006e4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dc8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006e5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006e6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dcc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006e7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006e8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dd0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006e9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dd2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006ea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dd4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006eb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dd6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006ec] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dd8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006ed] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dda] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006ee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ddc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006ef] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dde] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006f0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00de0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006f1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00de2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006f2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00de4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006f3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00de6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006f4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00de8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006f5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006f6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006f7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006f8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00df0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006f9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00df2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006fa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00df4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006fb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00df6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006fc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00df8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006fd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dfa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006fe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dfc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006ff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00dfe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00700] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e00] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00701] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e02] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00702] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e04] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00703] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e06] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00704] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e08] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00705] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e0a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00706] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e0c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00707] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e0e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00708] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e10] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00709] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e12] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0070a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e14] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0070b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e16] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0070c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e18] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0070d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e1a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0070e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e1c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0070f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e1e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00710] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e20] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00711] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e22] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00712] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e24] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00713] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e26] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00714] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e28] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00715] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e2a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00716] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e2c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00717] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e2e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00718] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e30] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00719] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e32] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0071a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e34] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0071b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e36] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0071c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e38] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0071d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e3a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0071e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e3c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0071f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e3e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00720] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e40] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00721] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e42] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00722] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e44] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00723] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e46] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00724] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e48] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00725] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e4a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00726] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e4c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00727] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e4e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00728] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e50] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00729] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e52] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0072a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e54] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0072b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e56] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0072c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e58] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0072d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e5a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0072e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e5c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0072f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e5e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00730] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e60] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00731] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e62] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00732] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e64] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00733] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e66] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00734] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e68] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00735] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e6a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00736] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e6c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00737] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e6e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00738] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e70] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00739] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e72] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0073a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e74] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0073b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e76] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0073c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e78] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0073d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e7a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0073e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e7c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0073f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e7e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00740] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e80] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00741] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e82] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00742] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e84] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00743] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e86] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00744] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e88] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00745] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e8a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00746] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e8c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00747] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e8e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00748] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e90] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00749] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e92] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0074a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e94] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0074b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e96] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0074c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e98] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0074d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e9a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0074e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e9c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0074f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00e9e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00750] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ea0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00751] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ea2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00752] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ea4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00753] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ea6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00754] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ea8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00755] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eaa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00756] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00757] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00758] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eb0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00759] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eb2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0075a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eb4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0075b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eb6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0075c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eb8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0075d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0075e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ebc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0075f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ebe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00760] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ec0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00761] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ec2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00762] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ec4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00763] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ec6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00764] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ec8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00765] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00766] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ecc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00767] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ece] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00768] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ed0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00769] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ed2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0076a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ed4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0076b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ed6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0076c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ed8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0076d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eda] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0076e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00edc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0076f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ede] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00770] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ee0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00771] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ee2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00772] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ee4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00773] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ee6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00774] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ee8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00775] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00776] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00777] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00eee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00778] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ef0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00779] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ef2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0077a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ef4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0077b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ef6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0077c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ef8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0077d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00efa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0077e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00efc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0077f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00efe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00780] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f00] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00781] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f02] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00782] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f04] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00783] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f06] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00784] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f08] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00785] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f0a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00786] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f0c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00787] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f0e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00788] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f10] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00789] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f12] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0078a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f14] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0078b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f16] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0078c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f18] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0078d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f1a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0078e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f1c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0078f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f1e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00790] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f20] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00791] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f22] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00792] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f24] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00793] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f26] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00794] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f28] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00795] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f2a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00796] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f2c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00797] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f2e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00798] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f30] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00799] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f32] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0079a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f34] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0079b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f36] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0079c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f38] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0079d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f3a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0079e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f3c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0079f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f3e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007a0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f40] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007a1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f42] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007a2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f44] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007a3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f46] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007a4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f48] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007a5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f4a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007a6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f4c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007a7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f4e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007a8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f50] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007a9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f52] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007aa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f54] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007ab] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f56] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007ac] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f58] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007ad] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f5a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007ae] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f5c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007af] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f5e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007b0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f60] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007b1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f62] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007b2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f64] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007b3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f66] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007b4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f68] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007b5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f6a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007b6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f6c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007b7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f6e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007b8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f70] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007b9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f72] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007ba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f74] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007bb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f76] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007bc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f78] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007bd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f7a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007be] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f7c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007bf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f7e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007c0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f80] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007c1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f82] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007c2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f84] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007c3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f86] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007c4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f88] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007c5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f8a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007c6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f8c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007c7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f8e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007c8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f90] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007c9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f92] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007ca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f94] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007cb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f96] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007cc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f98] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007cd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f9a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007ce] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f9c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007cf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00f9e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007d0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fa0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007d1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fa2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007d2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fa4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007d3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fa6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007d4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fa8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007d5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00faa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007d6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007d7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007d8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fb0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007d9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fb2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007da] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fb4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007db] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fb6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007dc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fb8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007dd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007de] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fbc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007df] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fbe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007e0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fc0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007e1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fc2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007e2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fc4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007e3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fc6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007e4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fc8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007e5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007e6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fcc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007e7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007e8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fd0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007e9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fd2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007ea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fd4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007eb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fd6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007ec] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fd8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007ed] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fda] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007ee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fdc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007ef] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fde] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007f0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fe0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007f1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fe2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007f2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fe4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007f3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fe6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007f4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fe8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007f5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007f6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007f7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00fee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007f8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ff0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007f9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ff2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007fa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ff4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007fb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ff6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007fc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ff8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007fd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ffa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007fe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ffc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007ff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h00ffe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00800] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01000] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00801] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01002] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00802] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01004] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00803] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01006] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00804] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01008] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00805] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0100a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00806] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0100c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00807] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0100e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00808] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01010] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00809] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01012] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0080a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01014] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0080b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01016] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0080c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01018] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0080d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0101a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0080e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0101c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0080f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0101e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00810] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01020] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00811] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01022] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00812] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01024] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00813] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01026] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00814] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01028] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00815] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0102a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00816] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0102c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00817] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0102e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00818] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01030] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00819] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01032] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0081a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01034] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0081b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01036] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0081c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01038] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0081d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0103a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0081e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0103c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0081f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0103e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00820] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01040] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00821] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01042] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00822] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01044] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00823] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01046] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00824] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01048] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00825] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0104a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00826] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0104c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00827] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0104e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00828] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01050] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00829] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01052] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0082a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01054] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0082b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01056] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0082c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01058] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0082d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0105a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0082e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0105c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0082f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0105e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00830] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01060] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00831] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01062] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00832] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01064] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00833] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01066] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00834] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01068] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00835] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0106a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00836] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0106c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00837] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0106e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00838] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01070] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00839] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01072] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0083a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01074] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0083b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01076] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0083c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01078] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0083d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0107a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0083e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0107c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0083f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0107e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00840] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01080] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00841] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01082] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00842] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01084] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00843] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01086] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00844] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01088] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00845] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0108a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00846] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0108c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00847] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0108e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00848] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01090] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00849] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01092] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0084a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01094] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0084b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01096] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0084c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01098] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0084d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0109a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0084e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0109c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0084f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0109e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00850] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00851] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00852] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00853] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00854] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00855] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00856] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00857] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00858] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00859] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0085a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0085b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0085c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0085d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0085e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0085f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00860] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00861] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00862] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00863] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00864] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00865] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00866] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00867] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00868] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00869] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0086a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0086b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0086c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0086d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0086e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0086f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00870] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00871] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00872] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00873] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00874] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00875] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00876] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00877] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00878] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00879] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0087a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0087b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0087c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0087d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0087e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0087f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h010fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00880] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01100] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00881] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01102] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00882] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01104] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00883] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01106] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00884] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01108] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00885] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0110a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00886] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0110c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00887] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0110e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00888] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01110] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00889] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01112] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0088a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01114] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0088b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01116] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0088c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01118] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0088d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0111a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0088e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0111c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0088f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0111e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00890] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01120] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00891] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01122] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00892] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01124] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00893] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01126] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00894] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01128] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00895] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0112a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00896] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0112c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00897] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0112e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00898] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01130] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00899] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01132] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0089a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01134] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0089b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01136] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0089c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01138] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0089d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0113a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0089e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0113c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0089f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0113e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008a0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01140] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008a1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01142] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008a2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01144] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008a3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01146] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008a4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01148] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008a5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0114a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008a6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0114c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008a7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0114e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008a8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01150] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008a9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01152] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008aa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01154] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008ab] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01156] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008ac] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01158] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008ad] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0115a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008ae] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0115c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008af] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0115e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008b0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01160] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008b1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01162] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008b2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01164] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008b3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01166] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008b4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01168] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008b5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0116a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008b6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0116c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008b7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0116e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008b8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01170] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008b9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01172] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008ba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01174] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008bb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01176] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008bc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01178] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008bd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0117a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008be] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0117c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008bf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0117e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008c0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01180] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008c1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01182] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008c2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01184] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008c3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01186] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008c4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01188] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008c5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0118a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008c6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0118c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008c7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0118e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008c8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01190] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008c9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01192] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008ca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01194] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008cb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01196] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008cc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01198] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008cd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0119a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008ce] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0119c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008cf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0119e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008d0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008d1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008d2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008d3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008d4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008d5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008d6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008d7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008d8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008d9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008da] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008db] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008dc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008dd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008de] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008df] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008e0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008e1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008e2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008e3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008e4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008e5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008e6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008e7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008e8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008e9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008ea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008eb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008ec] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008ed] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008ee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008ef] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008f0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008f1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008f2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008f3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008f4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008f5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008f6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008f7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008f8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008f9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008fa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008fb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008fc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008fd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008fe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008ff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h011fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00900] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01200] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00901] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01202] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00902] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01204] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00903] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01206] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00904] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01208] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00905] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0120a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00906] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0120c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00907] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0120e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00908] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01210] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00909] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01212] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0090a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01214] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0090b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01216] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0090c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01218] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0090d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0121a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0090e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0121c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0090f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0121e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00910] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01220] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00911] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01222] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00912] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01224] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00913] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01226] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00914] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01228] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00915] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0122a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00916] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0122c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00917] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0122e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00918] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01230] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00919] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01232] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0091a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01234] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0091b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01236] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0091c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01238] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0091d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0123a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0091e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0123c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0091f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0123e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00920] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01240] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00921] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01242] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00922] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01244] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00923] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01246] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00924] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01248] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00925] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0124a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00926] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0124c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00927] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0124e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00928] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01250] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00929] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01252] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0092a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01254] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0092b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01256] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0092c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01258] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0092d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0125a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0092e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0125c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0092f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0125e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00930] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01260] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00931] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01262] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00932] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01264] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00933] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01266] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00934] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01268] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00935] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0126a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00936] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0126c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00937] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0126e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00938] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01270] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00939] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01272] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0093a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01274] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0093b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01276] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0093c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01278] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0093d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0127a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0093e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0127c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0093f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0127e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00940] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01280] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00941] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01282] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00942] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01284] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00943] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01286] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00944] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01288] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00945] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0128a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00946] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0128c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00947] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0128e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00948] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01290] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00949] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01292] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0094a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01294] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0094b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01296] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0094c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01298] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0094d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0129a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0094e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0129c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0094f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0129e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00950] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00951] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00952] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00953] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00954] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00955] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00956] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00957] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00958] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00959] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0095a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0095b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0095c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0095d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0095e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0095f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00960] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00961] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00962] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00963] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00964] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00965] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00966] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00967] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00968] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00969] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0096a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0096b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0096c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0096d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0096e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0096f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00970] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00971] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00972] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00973] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00974] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00975] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00976] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00977] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00978] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00979] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0097a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0097b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0097c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0097d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0097e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0097f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h012fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00980] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01300] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00981] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01302] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00982] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01304] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00983] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01306] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00984] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01308] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00985] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0130a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00986] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0130c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00987] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0130e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00988] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01310] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00989] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01312] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0098a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01314] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0098b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01316] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0098c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01318] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0098d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0131a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0098e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0131c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0098f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0131e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00990] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01320] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00991] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01322] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00992] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01324] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00993] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01326] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00994] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01328] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00995] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0132a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00996] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0132c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00997] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0132e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00998] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01330] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00999] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01332] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0099a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01334] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0099b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01336] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0099c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01338] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0099d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0133a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0099e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0133c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0099f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0133e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009a0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01340] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009a1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01342] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009a2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01344] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009a3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01346] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009a4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01348] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009a5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0134a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009a6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0134c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009a7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0134e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009a8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01350] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009a9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01352] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009aa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01354] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009ab] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01356] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009ac] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01358] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009ad] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0135a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009ae] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0135c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009af] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0135e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009b0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01360] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009b1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01362] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009b2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01364] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009b3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01366] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009b4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01368] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009b5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0136a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009b6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0136c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009b7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0136e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009b8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01370] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009b9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01372] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009ba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01374] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009bb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01376] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009bc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01378] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009bd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0137a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009be] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0137c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009bf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0137e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009c0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01380] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009c1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01382] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009c2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01384] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009c3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01386] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009c4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01388] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009c5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0138a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009c6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0138c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009c7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0138e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009c8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01390] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009c9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01392] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009ca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01394] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009cb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01396] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009cc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01398] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009cd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0139a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009ce] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0139c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009cf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0139e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009d0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009d1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009d2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009d3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009d4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009d5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009d6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009d7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009d8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009d9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009da] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009db] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009dc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009dd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009de] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009df] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009e0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009e1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009e2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009e3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009e4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009e5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009e6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009e7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009e8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009e9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009ea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009eb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009ec] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009ed] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009ee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009ef] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009f0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009f1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009f2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009f3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009f4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009f5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009f6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009f7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009f8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009f9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009fa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009fb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009fc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009fd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009fe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009ff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h013fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a00] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01400] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a01] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01402] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a02] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01404] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a03] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01406] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a04] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01408] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a05] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0140a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a06] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0140c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a07] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0140e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a08] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01410] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a09] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01412] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a0a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01414] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a0b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01416] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a0c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01418] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a0d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0141a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a0e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0141c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a0f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0141e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a10] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01420] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a11] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01422] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a12] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01424] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a13] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01426] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a14] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01428] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a15] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0142a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a16] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0142c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a17] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0142e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a18] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01430] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a19] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01432] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a1a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01434] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a1b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01436] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a1c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01438] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a1d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0143a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a1e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0143c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a1f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0143e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a20] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01440] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a21] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01442] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a22] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01444] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a23] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01446] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a24] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01448] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a25] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0144a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a26] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0144c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a27] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0144e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a28] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01450] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a29] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01452] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a2a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01454] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a2b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01456] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a2c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01458] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a2d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0145a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a2e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0145c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a2f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0145e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a30] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01460] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a31] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01462] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a32] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01464] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a33] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01466] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a34] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01468] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a35] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0146a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a36] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0146c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a37] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0146e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a38] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01470] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a39] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01472] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a3a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01474] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a3b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01476] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a3c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01478] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a3d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0147a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a3e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0147c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a3f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0147e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a40] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01480] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a41] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01482] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a42] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01484] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a43] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01486] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a44] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01488] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a45] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0148a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a46] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0148c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a47] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0148e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a48] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01490] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a49] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01492] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a4a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01494] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a4b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01496] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a4c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01498] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a4d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0149a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a4e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0149c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a4f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0149e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a50] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a51] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a52] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a53] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a54] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a55] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a56] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a57] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a58] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a59] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a5a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a5b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a5c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a5d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a5e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a5f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a60] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a61] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a62] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a63] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a64] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a65] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a66] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a67] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a68] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a69] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a6a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a6b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a6c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a6d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a6e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a6f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a70] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a71] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a72] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a73] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a74] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a75] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a76] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a77] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a78] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a79] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a7a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a7b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a7c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a7d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a7e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a7f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h014fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a80] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01500] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a81] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01502] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a82] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01504] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a83] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01506] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a84] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01508] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a85] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0150a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a86] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0150c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a87] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0150e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a88] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01510] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a89] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01512] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a8a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01514] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a8b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01516] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a8c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01518] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a8d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0151a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a8e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0151c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a8f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0151e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a90] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01520] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a91] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01522] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a92] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01524] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a93] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01526] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a94] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01528] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a95] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0152a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a96] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0152c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a97] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0152e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a98] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01530] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a99] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01532] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a9a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01534] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a9b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01536] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a9c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01538] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a9d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0153a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a9e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0153c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a9f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0153e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aa0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01540] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aa1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01542] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aa2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01544] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aa3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01546] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aa4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01548] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aa5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0154a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aa6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0154c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aa7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0154e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aa8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01550] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aa9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01552] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aaa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01554] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aab] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01556] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aac] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01558] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aad] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0155a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aae] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0155c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aaf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0155e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ab0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01560] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ab1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01562] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ab2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01564] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ab3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01566] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ab4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01568] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ab5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0156a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ab6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0156c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ab7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0156e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ab8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01570] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ab9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01572] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01574] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00abb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01576] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00abc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01578] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00abd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0157a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00abe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0157c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00abf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0157e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ac0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01580] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ac1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01582] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ac2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01584] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ac3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01586] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ac4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01588] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ac5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0158a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ac6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0158c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ac7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0158e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ac8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01590] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ac9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01592] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01594] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00acb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01596] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00acc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01598] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00acd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0159a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ace] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0159c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00acf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0159e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ad0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ad1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ad2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ad3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ad4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ad5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ad6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ad7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ad8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ad9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ada] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00adb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00adc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00add] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ade] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00adf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ae0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ae1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ae2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ae3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ae4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ae5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ae6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ae7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ae8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ae9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aeb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aec] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aed] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aef] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00af0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00af1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00af2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00af3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00af4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00af5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00af6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00af7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00af8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00af9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00afa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00afb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00afc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00afd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00afe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h015fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b00] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01600] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b01] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01602] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b02] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01604] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b03] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01606] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b04] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01608] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b05] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0160a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b06] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0160c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b07] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0160e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b08] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01610] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b09] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01612] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b0a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01614] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b0b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01616] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b0c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01618] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b0d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0161a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b0e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0161c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b0f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0161e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b10] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01620] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b11] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01622] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b12] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01624] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b13] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01626] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b14] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01628] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b15] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0162a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b16] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0162c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b17] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0162e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b18] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01630] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b19] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01632] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b1a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01634] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b1b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01636] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b1c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01638] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b1d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0163a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b1e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0163c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b1f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0163e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b20] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01640] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b21] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01642] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b22] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01644] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b23] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01646] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b24] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01648] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b25] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0164a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b26] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0164c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b27] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0164e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b28] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01650] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b29] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01652] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b2a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01654] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b2b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01656] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b2c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01658] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b2d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0165a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b2e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0165c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b2f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0165e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b30] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01660] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b31] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01662] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b32] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01664] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b33] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01666] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b34] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01668] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b35] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0166a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b36] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0166c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b37] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0166e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b38] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01670] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b39] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01672] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b3a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01674] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b3b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01676] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b3c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01678] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b3d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0167a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b3e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0167c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b3f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0167e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b40] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01680] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b41] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01682] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b42] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01684] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b43] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01686] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b44] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01688] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b45] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0168a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b46] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0168c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b47] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0168e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b48] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01690] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b49] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01692] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b4a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01694] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b4b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01696] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b4c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01698] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b4d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0169a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b4e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0169c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b4f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0169e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b50] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b51] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b52] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b53] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b54] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b55] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b56] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b57] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b58] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b59] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b5a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b5b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b5c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b5d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b5e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b5f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b60] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b61] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b62] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b63] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b64] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b65] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b66] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b67] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b68] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b69] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b6a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b6b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b6c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b6d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b6e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b6f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b70] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b71] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b72] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b73] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b74] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b75] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b76] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b77] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b78] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b79] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b7a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b7b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b7c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b7d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b7e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b7f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h016fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b80] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01700] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b81] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01702] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b82] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01704] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b83] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01706] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b84] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01708] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b85] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0170a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b86] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0170c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b87] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0170e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b88] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01710] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b89] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01712] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b8a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01714] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b8b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01716] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b8c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01718] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b8d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0171a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b8e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0171c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b8f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0171e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b90] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01720] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b91] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01722] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b92] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01724] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b93] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01726] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b94] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01728] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b95] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0172a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b96] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0172c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b97] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0172e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b98] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01730] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b99] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01732] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b9a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01734] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b9b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01736] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b9c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01738] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b9d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0173a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b9e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0173c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b9f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0173e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ba0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01740] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ba1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01742] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ba2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01744] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ba3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01746] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ba4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01748] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ba5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0174a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ba6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0174c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ba7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0174e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ba8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01750] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ba9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01752] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00baa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01754] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bab] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01756] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bac] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01758] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bad] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0175a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bae] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0175c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00baf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0175e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bb0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01760] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bb1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01762] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bb2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01764] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bb3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01766] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bb4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01768] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bb5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0176a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bb6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0176c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bb7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0176e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bb8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01770] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bb9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01772] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01774] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bbb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01776] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bbc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01778] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bbd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0177a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bbe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0177c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bbf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0177e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bc0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01780] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bc1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01782] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bc2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01784] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bc3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01786] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bc4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01788] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bc5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0178a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bc6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0178c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bc7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0178e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bc8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01790] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bc9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01792] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01794] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bcb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01796] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bcc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01798] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bcd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0179a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bce] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0179c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bcf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0179e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bd0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bd1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bd2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bd3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bd4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bd5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bd6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bd7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bd8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bd9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bda] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bdb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bdc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bdd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bde] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bdf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00be0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00be1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00be2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00be3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00be4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00be5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00be6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00be7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00be8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00be9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00beb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bec] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bed] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bef] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bf0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bf1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bf2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bf3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bf4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bf5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bf6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bf7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bf8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bf9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bfa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bfb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bfc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bfd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bfe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h017fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c00] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01800] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c01] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01802] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c02] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01804] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c03] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01806] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c04] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01808] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c05] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0180a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c06] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0180c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c07] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0180e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c08] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01810] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c09] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01812] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c0a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01814] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c0b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01816] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c0c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01818] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c0d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0181a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c0e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0181c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c0f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0181e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c10] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01820] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c11] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01822] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c12] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01824] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c13] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01826] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c14] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01828] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c15] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0182a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c16] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0182c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c17] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0182e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c18] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01830] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c19] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01832] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c1a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01834] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c1b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01836] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c1c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01838] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c1d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0183a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c1e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0183c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c1f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0183e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c20] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01840] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c21] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01842] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c22] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01844] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c23] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01846] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c24] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01848] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c25] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0184a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c26] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0184c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c27] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0184e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c28] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01850] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c29] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01852] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c2a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01854] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c2b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01856] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c2c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01858] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c2d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0185a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c2e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0185c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c2f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0185e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c30] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01860] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c31] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01862] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c32] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01864] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c33] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01866] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c34] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01868] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c35] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0186a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c36] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0186c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c37] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0186e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c38] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01870] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c39] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01872] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c3a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01874] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c3b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01876] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c3c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01878] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c3d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0187a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c3e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0187c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c3f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0187e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c40] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01880] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c41] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01882] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c42] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01884] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c43] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01886] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c44] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01888] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c45] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0188a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c46] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0188c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c47] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0188e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c48] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01890] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c49] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01892] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c4a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01894] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c4b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01896] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c4c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01898] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c4d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0189a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c4e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0189c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c4f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0189e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c50] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c51] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c52] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c53] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c54] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c55] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c56] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c57] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c58] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c59] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c5a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c5b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c5c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c5d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c5e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c5f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c60] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c61] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c62] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c63] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c64] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c65] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c66] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c67] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c68] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c69] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c6a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c6b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c6c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c6d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c6e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c6f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c70] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c71] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c72] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c73] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c74] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c75] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c76] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c77] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c78] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c79] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c7a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c7b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c7c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c7d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c7e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c7f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h018fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c80] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01900] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c81] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01902] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c82] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01904] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c83] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01906] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c84] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01908] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c85] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0190a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c86] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0190c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c87] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0190e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c88] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01910] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c89] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01912] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c8a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01914] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c8b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01916] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c8c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01918] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c8d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0191a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c8e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0191c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c8f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0191e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c90] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01920] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c91] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01922] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c92] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01924] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c93] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01926] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c94] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01928] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c95] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0192a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c96] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0192c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c97] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0192e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c98] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01930] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c99] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01932] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c9a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01934] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c9b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01936] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c9c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01938] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c9d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0193a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c9e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0193c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c9f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0193e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ca0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01940] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ca1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01942] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ca2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01944] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ca3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01946] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ca4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01948] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ca5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0194a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ca6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0194c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ca7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0194e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ca8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01950] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ca9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01952] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00caa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01954] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cab] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01956] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cac] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01958] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cad] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0195a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cae] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0195c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00caf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0195e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cb0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01960] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cb1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01962] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cb2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01964] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cb3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01966] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cb4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01968] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cb5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0196a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cb6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0196c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cb7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0196e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cb8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01970] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cb9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01972] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01974] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cbb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01976] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cbc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01978] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cbd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0197a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cbe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0197c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cbf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0197e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cc0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01980] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cc1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01982] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cc2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01984] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cc3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01986] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cc4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01988] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cc5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0198a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cc6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0198c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cc7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0198e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cc8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01990] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cc9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01992] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01994] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ccb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01996] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ccc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01998] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ccd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0199a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cce] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0199c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ccf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0199e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cd0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cd1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cd2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cd3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cd4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cd5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cd6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cd7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cd8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cd9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cda] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cdb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cdc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cdd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cde] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cdf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ce0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ce1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ce2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ce3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ce4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ce5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ce6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ce7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ce8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ce9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ceb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cec] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ced] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cef] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cf0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cf1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cf2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cf3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cf4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cf5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cf6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cf7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cf8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cf9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cfa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cfb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cfc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cfd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cfe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h019fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d00] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a00] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d01] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a02] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d02] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a04] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d03] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a06] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d04] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a08] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d05] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a0a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d06] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a0c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d07] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a0e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d08] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a10] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d09] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a12] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d0a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a14] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d0b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a16] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d0c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a18] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d0d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a1a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d0e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a1c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d0f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a1e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d10] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a20] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d11] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a22] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d12] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a24] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d13] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a26] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d14] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a28] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d15] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a2a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d16] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a2c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d17] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a2e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d18] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a30] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d19] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a32] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d1a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a34] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d1b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a36] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d1c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a38] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d1d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a3a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d1e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a3c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d1f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a3e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d20] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a40] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d21] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a42] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d22] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a44] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d23] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a46] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d24] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a48] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d25] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a4a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d26] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a4c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d27] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a4e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d28] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a50] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d29] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a52] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d2a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a54] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d2b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a56] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d2c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a58] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d2d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a5a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d2e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a5c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d2f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a5e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d30] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a60] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d31] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a62] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d32] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a64] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d33] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a66] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d34] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a68] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d35] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a6a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d36] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a6c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d37] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a6e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d38] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a70] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d39] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a72] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d3a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a74] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d3b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a76] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d3c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a78] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d3d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a7a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d3e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a7c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d3f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a7e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d40] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a80] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d41] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a82] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d42] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a84] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d43] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a86] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d44] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a88] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d45] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a8a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d46] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a8c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d47] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a8e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d48] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a90] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d49] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a92] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d4a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a94] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d4b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a96] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d4c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a98] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d4d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a9a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d4e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a9c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d4f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01a9e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d50] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aa0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d51] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aa2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d52] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aa4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d53] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aa6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d54] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aa8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d55] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aaa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d56] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d57] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d58] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ab0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d59] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ab2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d5a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ab4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d5b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ab6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d5c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ab8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d5d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d5e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01abc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d5f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01abe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d60] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ac0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d61] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ac2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d62] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ac4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d63] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ac6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d64] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ac8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d65] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d66] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01acc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d67] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ace] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d68] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ad0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d69] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ad2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d6a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ad4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d6b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ad6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d6c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ad8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d6d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ada] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d6e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01adc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d6f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ade] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d70] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ae0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d71] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ae2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d72] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ae4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d73] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ae6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d74] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ae8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d75] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d76] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d77] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01aee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d78] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01af0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d79] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01af2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d7a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01af4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d7b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01af6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d7c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01af8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d7d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01afa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d7e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01afc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d7f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01afe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d80] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b00] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d81] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b02] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d82] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b04] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d83] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b06] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d84] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b08] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d85] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b0a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d86] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b0c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d87] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b0e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d88] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b10] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d89] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b12] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d8a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b14] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d8b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b16] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d8c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b18] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d8d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b1a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d8e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b1c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d8f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b1e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d90] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b20] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d91] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b22] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d92] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b24] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d93] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b26] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d94] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b28] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d95] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b2a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d96] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b2c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d97] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b2e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d98] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b30] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d99] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b32] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d9a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b34] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d9b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b36] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d9c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b38] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d9d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b3a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d9e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b3c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d9f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b3e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00da0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b40] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00da1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b42] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00da2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b44] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00da3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b46] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00da4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b48] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00da5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b4a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00da6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b4c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00da7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b4e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00da8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b50] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00da9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b52] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00daa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b54] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dab] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b56] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dac] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b58] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dad] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b5a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dae] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b5c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00daf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b5e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00db0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b60] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00db1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b62] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00db2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b64] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00db3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b66] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00db4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b68] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00db5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b6a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00db6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b6c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00db7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b6e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00db8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b70] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00db9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b72] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b74] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dbb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b76] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dbc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b78] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dbd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b7a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dbe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b7c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dbf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b7e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dc0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b80] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dc1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b82] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dc2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b84] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dc3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b86] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dc4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b88] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dc5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b8a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dc6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b8c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dc7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b8e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dc8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b90] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dc9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b92] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b94] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dcb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b96] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dcc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b98] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dcd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b9a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dce] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b9c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dcf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01b9e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dd0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ba0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dd1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ba2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dd2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ba4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dd3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ba6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dd4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ba8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dd5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01baa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dd6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dd7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dd8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bb0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dd9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bb2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dda] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bb4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ddb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bb6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ddc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bb8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ddd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dde] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bbc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ddf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bbe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00de0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bc0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00de1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bc2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00de2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bc4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00de3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bc6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00de4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bc8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00de5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00de6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bcc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00de7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00de8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bd0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00de9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bd2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bd4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00deb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bd6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dec] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bd8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ded] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bda] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bdc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00def] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bde] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00df0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01be0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00df1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01be2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00df2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01be4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00df3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01be6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00df4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01be8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00df5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00df6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00df7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00df8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bf0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00df9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bf2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dfa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bf4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dfb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bf6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dfc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bf8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dfd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bfa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dfe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bfc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01bfe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e00] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c00] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e01] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c02] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e02] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c04] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e03] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c06] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e04] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c08] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e05] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c0a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e06] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c0c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e07] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c0e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e08] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c10] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e09] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c12] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e0a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c14] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e0b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c16] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e0c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c18] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e0d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c1a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e0e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c1c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e0f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c1e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e10] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c20] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e11] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c22] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e12] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c24] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e13] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c26] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e14] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c28] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e15] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c2a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e16] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c2c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e17] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c2e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e18] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c30] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e19] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c32] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e1a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c34] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e1b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c36] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e1c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c38] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e1d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c3a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e1e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c3c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e1f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c3e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e20] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c40] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e21] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c42] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e22] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c44] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e23] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c46] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e24] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c48] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e25] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c4a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e26] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c4c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e27] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c4e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e28] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c50] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e29] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c52] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e2a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c54] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e2b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c56] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e2c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c58] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e2d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c5a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e2e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c5c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e2f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c5e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e30] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c60] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e31] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c62] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e32] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c64] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e33] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c66] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e34] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c68] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e35] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c6a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e36] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c6c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e37] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c6e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e38] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c70] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e39] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c72] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e3a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c74] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e3b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c76] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e3c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c78] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e3d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c7a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e3e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c7c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e3f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c7e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e40] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c80] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e41] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c82] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e42] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c84] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e43] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c86] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e44] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c88] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e45] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c8a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e46] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c8c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e47] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c8e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e48] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c90] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e49] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c92] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e4a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c94] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e4b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c96] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e4c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c98] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e4d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c9a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e4e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c9c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e4f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01c9e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e50] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ca0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e51] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ca2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e52] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ca4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e53] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ca6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e54] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ca8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e55] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01caa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e56] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e57] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e58] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cb0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e59] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cb2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e5a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cb4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e5b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cb6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e5c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cb8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e5d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e5e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cbc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e5f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cbe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e60] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cc0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e61] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cc2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e62] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cc4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e63] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cc6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e64] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cc8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e65] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e66] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ccc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e67] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e68] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cd0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e69] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cd2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e6a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cd4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e6b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cd6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e6c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cd8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e6d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cda] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e6e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cdc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e6f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cde] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e70] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ce0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e71] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ce2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e72] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ce4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e73] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ce6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e74] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ce8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e75] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e76] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e77] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e78] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cf0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e79] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cf2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e7a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cf4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e7b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cf6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e7c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cf8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e7d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cfa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e7e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cfc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e7f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01cfe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e80] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d00] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e81] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d02] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e82] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d04] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e83] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d06] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e84] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d08] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e85] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d0a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e86] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d0c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e87] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d0e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e88] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d10] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e89] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d12] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e8a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d14] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e8b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d16] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e8c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d18] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e8d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d1a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e8e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d1c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e8f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d1e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e90] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d20] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e91] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d22] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e92] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d24] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e93] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d26] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e94] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d28] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e95] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d2a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e96] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d2c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e97] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d2e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e98] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d30] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e99] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d32] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e9a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d34] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e9b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d36] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e9c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d38] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e9d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d3a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e9e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d3c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e9f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d3e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ea0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d40] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ea1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d42] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ea2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d44] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ea3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d46] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ea4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d48] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ea5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d4a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ea6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d4c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ea7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d4e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ea8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d50] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ea9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d52] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eaa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d54] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eab] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d56] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eac] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d58] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ead] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d5a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eae] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d5c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eaf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d5e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eb0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d60] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eb1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d62] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eb2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d64] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eb3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d66] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eb4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d68] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eb5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d6a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eb6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d6c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eb7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d6e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eb8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d70] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eb9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d72] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d74] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ebb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d76] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ebc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d78] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ebd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d7a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ebe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d7c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ebf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d7e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ec0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d80] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ec1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d82] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ec2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d84] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ec3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d86] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ec4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d88] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ec5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d8a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ec6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d8c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ec7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d8e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ec8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d90] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ec9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d92] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d94] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ecb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d96] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ecc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d98] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ecd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d9a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ece] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d9c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ecf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01d9e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ed0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01da0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ed1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01da2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ed2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01da4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ed3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01da6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ed4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01da8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ed5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01daa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ed6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ed7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ed8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01db0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ed9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01db2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eda] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01db4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00edb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01db6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00edc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01db8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00edd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ede] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dbc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00edf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dbe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ee0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dc0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ee1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dc2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ee2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dc4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ee3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dc6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ee4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dc8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ee5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ee6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dcc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ee7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ee8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dd0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ee9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dd2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dd4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eeb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dd6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eec] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dd8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eed] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dda] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ddc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eef] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dde] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ef0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01de0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ef1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01de2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ef2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01de4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ef3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01de6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ef4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01de8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ef5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ef6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ef7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ef8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01df0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ef9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01df2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00efa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01df4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00efb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01df6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00efc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01df8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00efd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dfa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00efe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dfc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01dfe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f00] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e00] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f01] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e02] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f02] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e04] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f03] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e06] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f04] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e08] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f05] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e0a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f06] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e0c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f07] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e0e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f08] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e10] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f09] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e12] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f0a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e14] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f0b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e16] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f0c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e18] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f0d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e1a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f0e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e1c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f0f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e1e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f10] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e20] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f11] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e22] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f12] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e24] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f13] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e26] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f14] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e28] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f15] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e2a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f16] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e2c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f17] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e2e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f18] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e30] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f19] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e32] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f1a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e34] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f1b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e36] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f1c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e38] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f1d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e3a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f1e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e3c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f1f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e3e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f20] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e40] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f21] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e42] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f22] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e44] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f23] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e46] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f24] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e48] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f25] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e4a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f26] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e4c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f27] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e4e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f28] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e50] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f29] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e52] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f2a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e54] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f2b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e56] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f2c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e58] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f2d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e5a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f2e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e5c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f2f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e5e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f30] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e60] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f31] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e62] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f32] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e64] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f33] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e66] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f34] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e68] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f35] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e6a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f36] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e6c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f37] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e6e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f38] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e70] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f39] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e72] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f3a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e74] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f3b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e76] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f3c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e78] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f3d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e7a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f3e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e7c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f3f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e7e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f40] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e80] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f41] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e82] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f42] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e84] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f43] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e86] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f44] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e88] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f45] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e8a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f46] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e8c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f47] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e8e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f48] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e90] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f49] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e92] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f4a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e94] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f4b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e96] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f4c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e98] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f4d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e9a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f4e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e9c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f4f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01e9e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f50] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ea0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f51] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ea2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f52] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ea4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f53] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ea6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f54] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ea8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f55] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eaa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f56] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f57] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f58] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eb0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f59] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eb2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f5a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eb4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f5b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eb6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f5c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eb8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f5d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f5e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ebc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f5f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ebe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f60] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ec0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f61] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ec2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f62] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ec4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f63] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ec6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f64] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ec8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f65] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f66] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ecc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f67] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ece] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f68] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ed0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f69] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ed2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f6a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ed4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f6b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ed6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f6c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ed8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f6d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eda] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f6e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01edc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f6f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ede] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f70] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ee0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f71] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ee2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f72] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ee4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f73] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ee6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f74] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ee8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f75] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f76] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f77] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01eee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f78] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ef0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f79] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ef2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f7a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ef4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f7b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ef6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f7c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ef8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f7d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01efa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f7e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01efc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f7f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01efe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f80] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f00] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f81] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f02] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f82] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f04] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f83] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f06] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f84] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f08] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f85] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f0a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f86] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f0c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f87] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f0e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f88] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f10] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f89] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f12] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f8a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f14] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f8b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f16] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f8c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f18] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f8d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f1a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f8e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f1c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f8f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f1e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f90] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f20] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f91] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f22] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f92] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f24] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f93] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f26] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f94] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f28] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f95] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f2a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f96] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f2c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f97] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f2e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f98] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f30] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f99] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f32] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f9a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f34] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f9b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f36] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f9c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f38] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f9d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f3a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f9e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f3c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f9f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f3e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fa0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f40] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fa1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f42] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fa2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f44] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fa3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f46] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fa4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f48] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fa5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f4a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fa6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f4c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fa7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f4e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fa8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f50] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fa9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f52] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00faa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f54] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fab] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f56] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fac] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f58] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fad] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f5a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fae] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f5c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00faf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f5e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fb0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f60] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fb1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f62] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fb2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f64] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fb3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f66] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fb4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f68] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fb5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f6a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fb6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f6c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fb7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f6e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fb8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f70] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fb9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f72] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f74] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fbb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f76] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fbc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f78] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fbd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f7a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fbe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f7c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fbf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f7e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fc0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f80] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fc1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f82] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fc2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f84] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fc3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f86] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fc4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f88] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fc5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f8a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fc6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f8c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fc7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f8e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fc8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f90] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fc9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f92] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f94] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fcb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f96] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fcc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f98] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fcd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f9a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fce] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f9c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fcf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01f9e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fd0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fa0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fd1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fa2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fd2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fa4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fd3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fa6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fd4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fa8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fd5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01faa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fd6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fd7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fd8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fb0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fd9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fb2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fda] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fb4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fdb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fb6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fdc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fb8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fdd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fde] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fbc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fdf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fbe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fe0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fc0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fe1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fc2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fe2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fc4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fe3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fc6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fe4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fc8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fe5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fe6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fcc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fe7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fe8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fd0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fe9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fd2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fd4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00feb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fd6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fec] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fd8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fed] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fda] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fdc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fef] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fde] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ff0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fe0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ff1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fe2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ff2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fe4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ff3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fe6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ff4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fe8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ff5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ff6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ff7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01fee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ff8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ff0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ff9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ff2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ffa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ff4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ffb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ff6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ffc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ff8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ffd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ffa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ffe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ffc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h01ffe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01000] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02000] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01001] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02002] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01002] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02004] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01003] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02006] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01004] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02008] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01005] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0200a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01006] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0200c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01007] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0200e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01008] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02010] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01009] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02012] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0100a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02014] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0100b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02016] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0100c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02018] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0100d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0201a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0100e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0201c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0100f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0201e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01010] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02020] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01011] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02022] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01012] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02024] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01013] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02026] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01014] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02028] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01015] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0202a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01016] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0202c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01017] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0202e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01018] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02030] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01019] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02032] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0101a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02034] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0101b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02036] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0101c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02038] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0101d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0203a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0101e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0203c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0101f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0203e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01020] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02040] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01021] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02042] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01022] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02044] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01023] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02046] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01024] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02048] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01025] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0204a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01026] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0204c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01027] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0204e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01028] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02050] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01029] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02052] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0102a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02054] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0102b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02056] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0102c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02058] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0102d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0205a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0102e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0205c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0102f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0205e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01030] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02060] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01031] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02062] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01032] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02064] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01033] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02066] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01034] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02068] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01035] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0206a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01036] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0206c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01037] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0206e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01038] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02070] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01039] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02072] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0103a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02074] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0103b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02076] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0103c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02078] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0103d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0207a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0103e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0207c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0103f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0207e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01040] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02080] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01041] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02082] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01042] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02084] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01043] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02086] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01044] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02088] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01045] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0208a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01046] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0208c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01047] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0208e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01048] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02090] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01049] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02092] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0104a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02094] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0104b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02096] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0104c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02098] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0104d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0209a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0104e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0209c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0104f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0209e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01050] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01051] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01052] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01053] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01054] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01055] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01056] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01057] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01058] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01059] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0105a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0105b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0105c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0105d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0105e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0105f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01060] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01061] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01062] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01063] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01064] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01065] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01066] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01067] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01068] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01069] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0106a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0106b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0106c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0106d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0106e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0106f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01070] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01071] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01072] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01073] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01074] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01075] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01076] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01077] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01078] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01079] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0107a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0107b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0107c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0107d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0107e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0107f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h020fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01080] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02100] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01081] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02102] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01082] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02104] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01083] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02106] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01084] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02108] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01085] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0210a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01086] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0210c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01087] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0210e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01088] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02110] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01089] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02112] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0108a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02114] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0108b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02116] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0108c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02118] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0108d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0211a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0108e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0211c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0108f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0211e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01090] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02120] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01091] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02122] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01092] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02124] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01093] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02126] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01094] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02128] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01095] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0212a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01096] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0212c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01097] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0212e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01098] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02130] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01099] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02132] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0109a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02134] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0109b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02136] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0109c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02138] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0109d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0213a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0109e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0213c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0109f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0213e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010a0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02140] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010a1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02142] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010a2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02144] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010a3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02146] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010a4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02148] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010a5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0214a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010a6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0214c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010a7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0214e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010a8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02150] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010a9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02152] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010aa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02154] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010ab] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02156] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010ac] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02158] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010ad] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0215a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010ae] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0215c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010af] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0215e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010b0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02160] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010b1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02162] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010b2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02164] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010b3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02166] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010b4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02168] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010b5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0216a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010b6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0216c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010b7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0216e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010b8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02170] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010b9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02172] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010ba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02174] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010bb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02176] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010bc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02178] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010bd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0217a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010be] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0217c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010bf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0217e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010c0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02180] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010c1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02182] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010c2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02184] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010c3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02186] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010c4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02188] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010c5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0218a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010c6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0218c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010c7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0218e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010c8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02190] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010c9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02192] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010ca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02194] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010cb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02196] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010cc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02198] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010cd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0219a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010ce] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0219c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010cf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0219e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010d0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010d1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010d2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010d3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010d4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010d5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010d6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010d7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010d8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010d9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010da] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010db] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010dc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010dd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010de] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010df] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010e0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010e1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010e2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010e3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010e4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010e5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010e6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010e7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010e8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010e9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010ea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010eb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010ec] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010ed] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010ee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010ef] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010f0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010f1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010f2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010f3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010f4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010f5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010f6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010f7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010f8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010f9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010fa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010fb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010fc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010fd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010fe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010ff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h021fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01100] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02200] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01101] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02202] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01102] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02204] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01103] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02206] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01104] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02208] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01105] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0220a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01106] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0220c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01107] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0220e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01108] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02210] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01109] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02212] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0110a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02214] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0110b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02216] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0110c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02218] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0110d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0221a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0110e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0221c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0110f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0221e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01110] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02220] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01111] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02222] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01112] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02224] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01113] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02226] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01114] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02228] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01115] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0222a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01116] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0222c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01117] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0222e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01118] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02230] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01119] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02232] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0111a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02234] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0111b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02236] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0111c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02238] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0111d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0223a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0111e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0223c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0111f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0223e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01120] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02240] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01121] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02242] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01122] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02244] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01123] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02246] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01124] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02248] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01125] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0224a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01126] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0224c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01127] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0224e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01128] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02250] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01129] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02252] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0112a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02254] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0112b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02256] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0112c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02258] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0112d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0225a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0112e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0225c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0112f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0225e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01130] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02260] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01131] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02262] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01132] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02264] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01133] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02266] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01134] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02268] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01135] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0226a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01136] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0226c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01137] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0226e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01138] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02270] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01139] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02272] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0113a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02274] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0113b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02276] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0113c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02278] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0113d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0227a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0113e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0227c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0113f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0227e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01140] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02280] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01141] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02282] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01142] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02284] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01143] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02286] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01144] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02288] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01145] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0228a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01146] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0228c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01147] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0228e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01148] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02290] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01149] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02292] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0114a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02294] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0114b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02296] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0114c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02298] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0114d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0229a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0114e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0229c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0114f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0229e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01150] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01151] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01152] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01153] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01154] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01155] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01156] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01157] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01158] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01159] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0115a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0115b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0115c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0115d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0115e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0115f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01160] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01161] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01162] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01163] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01164] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01165] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01166] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01167] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01168] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01169] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0116a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0116b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0116c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0116d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0116e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0116f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01170] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01171] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01172] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01173] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01174] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01175] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01176] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01177] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01178] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01179] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0117a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0117b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0117c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0117d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0117e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0117f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h022fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01180] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02300] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01181] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02302] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01182] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02304] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01183] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02306] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01184] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02308] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01185] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0230a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01186] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0230c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01187] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0230e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01188] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02310] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01189] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02312] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0118a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02314] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0118b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02316] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0118c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02318] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0118d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0231a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0118e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0231c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0118f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0231e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01190] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02320] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01191] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02322] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01192] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02324] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01193] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02326] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01194] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02328] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01195] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0232a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01196] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0232c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01197] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0232e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01198] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02330] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01199] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02332] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0119a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02334] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0119b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02336] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0119c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02338] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0119d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0233a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0119e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0233c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0119f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0233e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011a0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02340] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011a1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02342] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011a2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02344] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011a3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02346] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011a4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02348] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011a5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0234a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011a6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0234c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011a7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0234e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011a8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02350] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011a9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02352] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011aa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02354] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011ab] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02356] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011ac] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02358] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011ad] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0235a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011ae] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0235c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011af] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0235e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011b0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02360] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011b1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02362] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011b2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02364] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011b3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02366] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011b4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02368] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011b5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0236a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011b6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0236c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011b7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0236e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011b8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02370] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011b9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02372] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011ba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02374] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011bb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02376] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011bc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02378] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011bd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0237a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011be] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0237c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011bf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0237e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011c0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02380] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011c1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02382] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011c2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02384] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011c3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02386] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011c4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02388] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011c5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0238a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011c6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0238c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011c7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0238e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011c8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02390] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011c9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02392] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011ca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02394] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011cb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02396] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011cc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02398] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011cd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0239a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011ce] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0239c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011cf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0239e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011d0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011d1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011d2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011d3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011d4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011d5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011d6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011d7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011d8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011d9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011da] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011db] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011dc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011dd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011de] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011df] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011e0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011e1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011e2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011e3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011e4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011e5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011e6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011e7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011e8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011e9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011ea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011eb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011ec] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011ed] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011ee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011ef] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011f0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011f1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011f2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011f3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011f4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011f5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011f6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011f7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011f8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011f9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011fa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011fb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011fc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011fd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011fe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011ff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h023fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01200] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02400] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01201] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02402] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01202] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02404] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01203] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02406] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01204] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02408] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01205] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0240a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01206] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0240c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01207] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0240e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01208] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02410] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01209] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02412] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0120a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02414] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0120b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02416] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0120c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02418] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0120d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0241a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0120e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0241c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0120f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0241e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01210] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02420] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01211] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02422] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01212] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02424] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01213] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02426] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01214] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02428] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01215] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0242a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01216] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0242c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01217] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0242e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01218] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02430] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01219] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02432] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0121a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02434] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0121b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02436] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0121c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02438] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0121d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0243a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0121e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0243c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0121f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0243e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01220] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02440] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01221] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02442] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01222] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02444] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01223] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02446] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01224] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02448] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01225] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0244a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01226] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0244c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01227] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0244e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01228] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02450] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01229] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02452] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0122a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02454] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0122b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02456] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0122c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02458] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0122d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0245a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0122e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0245c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0122f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0245e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01230] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02460] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01231] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02462] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01232] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02464] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01233] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02466] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01234] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02468] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01235] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0246a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01236] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0246c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01237] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0246e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01238] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02470] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01239] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02472] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0123a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02474] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0123b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02476] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0123c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02478] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0123d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0247a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0123e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0247c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0123f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0247e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01240] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02480] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01241] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02482] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01242] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02484] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01243] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02486] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01244] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02488] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01245] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0248a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01246] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0248c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01247] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0248e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01248] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02490] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01249] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02492] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0124a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02494] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0124b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02496] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0124c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02498] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0124d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0249a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0124e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0249c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0124f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0249e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01250] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01251] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01252] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01253] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01254] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01255] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01256] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01257] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01258] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01259] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0125a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0125b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0125c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0125d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0125e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0125f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01260] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01261] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01262] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01263] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01264] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01265] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01266] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01267] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01268] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01269] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0126a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0126b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0126c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0126d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0126e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0126f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01270] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01271] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01272] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01273] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01274] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01275] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01276] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01277] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01278] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01279] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0127a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0127b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0127c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0127d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0127e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0127f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h024fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01280] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02500] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01281] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02502] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01282] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02504] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01283] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02506] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01284] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02508] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01285] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0250a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01286] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0250c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01287] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0250e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01288] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02510] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01289] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02512] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0128a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02514] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0128b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02516] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0128c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02518] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0128d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0251a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0128e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0251c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0128f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0251e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01290] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02520] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01291] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02522] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01292] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02524] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01293] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02526] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01294] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02528] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01295] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0252a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01296] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0252c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01297] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0252e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01298] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02530] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01299] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02532] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0129a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02534] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0129b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02536] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0129c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02538] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0129d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0253a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0129e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0253c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0129f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0253e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012a0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02540] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012a1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02542] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012a2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02544] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012a3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02546] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012a4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02548] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012a5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0254a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012a6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0254c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012a7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0254e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012a8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02550] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012a9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02552] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012aa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02554] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012ab] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02556] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012ac] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02558] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012ad] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0255a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012ae] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0255c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012af] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0255e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012b0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02560] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012b1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02562] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012b2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02564] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012b3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02566] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012b4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02568] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012b5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0256a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012b6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0256c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012b7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0256e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012b8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02570] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012b9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02572] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012ba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02574] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012bb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02576] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012bc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02578] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012bd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0257a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012be] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0257c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012bf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0257e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012c0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02580] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012c1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02582] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012c2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02584] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012c3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02586] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012c4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02588] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012c5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0258a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012c6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0258c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012c7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0258e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012c8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02590] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012c9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02592] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012ca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02594] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012cb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02596] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012cc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02598] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012cd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0259a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012ce] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0259c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012cf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0259e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012d0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012d1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012d2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012d3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012d4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012d5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012d6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012d7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012d8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012d9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012da] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012db] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012dc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012dd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012de] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012df] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012e0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012e1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012e2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012e3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012e4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012e5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012e6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012e7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012e8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012e9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012ea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012eb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012ec] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012ed] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012ee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012ef] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012f0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012f1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012f2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012f3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012f4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012f5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012f6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012f7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012f8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012f9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012fa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012fb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012fc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012fd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012fe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012ff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h025fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01300] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02600] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01301] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02602] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01302] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02604] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01303] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02606] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01304] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02608] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01305] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0260a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01306] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0260c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01307] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0260e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01308] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02610] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01309] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02612] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0130a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02614] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0130b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02616] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0130c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02618] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0130d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0261a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0130e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0261c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0130f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0261e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01310] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02620] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01311] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02622] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01312] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02624] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01313] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02626] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01314] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02628] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01315] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0262a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01316] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0262c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01317] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0262e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01318] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02630] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01319] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02632] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0131a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02634] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0131b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02636] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0131c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02638] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0131d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0263a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0131e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0263c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0131f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0263e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01320] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02640] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01321] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02642] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01322] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02644] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01323] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02646] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01324] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02648] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01325] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0264a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01326] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0264c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01327] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0264e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01328] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02650] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01329] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02652] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0132a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02654] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0132b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02656] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0132c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02658] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0132d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0265a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0132e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0265c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0132f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0265e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01330] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02660] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01331] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02662] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01332] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02664] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01333] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02666] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01334] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02668] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01335] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0266a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01336] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0266c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01337] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0266e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01338] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02670] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01339] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02672] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0133a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02674] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0133b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02676] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0133c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02678] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0133d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0267a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0133e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0267c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0133f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0267e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01340] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02680] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01341] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02682] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01342] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02684] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01343] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02686] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01344] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02688] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01345] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0268a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01346] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0268c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01347] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0268e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01348] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02690] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01349] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02692] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0134a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02694] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0134b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02696] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0134c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02698] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0134d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0269a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0134e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0269c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0134f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0269e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01350] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01351] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01352] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01353] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01354] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01355] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01356] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01357] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01358] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01359] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0135a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0135b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0135c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0135d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0135e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0135f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01360] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01361] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01362] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01363] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01364] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01365] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01366] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01367] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01368] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01369] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0136a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0136b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0136c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0136d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0136e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0136f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01370] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01371] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01372] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01373] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01374] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01375] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01376] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01377] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01378] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01379] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0137a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0137b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0137c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0137d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0137e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0137f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h026fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01380] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02700] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01381] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02702] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01382] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02704] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01383] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02706] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01384] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02708] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01385] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0270a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01386] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0270c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01387] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0270e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01388] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02710] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01389] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02712] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0138a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02714] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0138b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02716] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0138c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02718] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0138d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0271a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0138e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0271c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0138f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0271e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01390] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02720] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01391] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02722] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01392] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02724] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01393] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02726] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01394] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02728] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01395] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0272a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01396] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0272c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01397] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0272e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01398] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02730] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01399] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02732] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0139a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02734] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0139b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02736] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0139c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02738] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0139d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0273a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0139e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0273c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0139f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0273e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013a0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02740] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013a1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02742] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013a2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02744] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013a3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02746] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013a4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02748] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013a5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0274a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013a6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0274c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013a7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0274e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013a8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02750] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013a9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02752] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013aa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02754] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013ab] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02756] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013ac] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02758] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013ad] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0275a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013ae] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0275c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013af] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0275e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013b0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02760] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013b1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02762] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013b2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02764] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013b3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02766] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013b4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02768] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013b5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0276a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013b6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0276c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013b7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0276e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013b8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02770] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013b9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02772] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013ba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02774] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013bb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02776] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013bc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02778] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013bd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0277a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013be] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0277c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013bf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0277e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013c0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02780] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013c1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02782] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013c2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02784] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013c3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02786] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013c4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02788] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013c5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0278a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013c6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0278c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013c7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0278e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013c8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02790] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013c9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02792] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013ca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02794] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013cb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02796] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013cc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02798] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013cd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0279a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013ce] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0279c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013cf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0279e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013d0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013d1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013d2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013d3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013d4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013d5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013d6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013d7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013d8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013d9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013da] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013db] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013dc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013dd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013de] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013df] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013e0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013e1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013e2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013e3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013e4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013e5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013e6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013e7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013e8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013e9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013ea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013eb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013ec] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013ed] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013ee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013ef] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013f0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013f1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013f2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013f3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013f4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013f5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013f6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013f7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013f8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013f9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013fa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013fb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013fc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013fd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013fe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013ff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h027fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01400] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02800] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01401] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02802] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01402] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02804] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01403] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02806] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01404] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02808] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01405] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0280a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01406] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0280c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01407] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0280e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01408] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02810] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01409] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02812] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0140a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02814] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0140b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02816] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0140c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02818] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0140d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0281a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0140e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0281c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0140f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0281e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01410] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02820] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01411] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02822] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01412] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02824] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01413] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02826] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01414] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02828] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01415] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0282a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01416] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0282c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01417] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0282e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01418] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02830] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01419] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02832] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0141a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02834] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0141b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02836] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0141c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02838] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0141d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0283a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0141e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0283c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0141f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0283e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01420] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02840] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01421] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02842] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01422] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02844] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01423] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02846] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01424] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02848] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01425] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0284a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01426] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0284c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01427] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0284e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01428] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02850] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01429] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02852] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0142a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02854] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0142b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02856] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0142c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02858] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0142d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0285a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0142e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0285c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0142f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0285e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01430] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02860] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01431] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02862] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01432] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02864] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01433] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02866] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01434] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02868] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01435] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0286a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01436] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0286c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01437] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0286e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01438] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02870] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01439] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02872] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0143a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02874] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0143b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02876] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0143c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02878] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0143d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0287a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0143e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0287c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0143f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0287e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01440] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02880] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01441] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02882] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01442] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02884] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01443] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02886] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01444] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02888] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01445] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0288a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01446] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0288c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01447] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0288e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01448] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02890] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01449] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02892] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0144a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02894] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0144b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02896] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0144c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02898] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0144d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0289a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0144e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0289c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0144f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0289e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01450] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01451] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01452] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01453] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01454] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01455] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01456] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01457] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01458] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01459] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0145a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0145b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0145c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0145d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0145e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0145f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01460] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01461] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01462] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01463] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01464] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01465] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01466] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01467] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01468] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01469] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0146a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0146b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0146c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0146d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0146e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0146f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01470] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01471] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01472] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01473] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01474] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01475] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01476] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01477] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01478] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01479] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0147a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0147b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0147c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0147d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0147e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0147f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h028fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01480] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02900] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01481] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02902] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01482] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02904] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01483] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02906] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01484] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02908] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01485] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0290a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01486] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0290c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01487] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0290e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01488] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02910] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01489] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02912] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0148a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02914] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0148b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02916] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0148c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02918] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0148d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0291a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0148e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0291c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0148f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0291e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01490] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02920] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01491] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02922] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01492] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02924] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01493] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02926] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01494] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02928] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01495] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0292a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01496] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0292c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01497] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0292e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01498] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02930] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01499] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02932] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0149a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02934] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0149b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02936] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0149c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02938] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0149d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0293a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0149e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0293c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0149f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0293e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014a0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02940] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014a1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02942] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014a2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02944] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014a3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02946] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014a4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02948] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014a5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0294a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014a6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0294c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014a7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0294e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014a8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02950] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014a9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02952] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014aa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02954] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014ab] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02956] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014ac] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02958] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014ad] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0295a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014ae] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0295c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014af] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0295e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014b0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02960] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014b1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02962] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014b2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02964] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014b3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02966] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014b4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02968] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014b5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0296a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014b6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0296c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014b7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0296e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014b8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02970] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014b9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02972] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014ba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02974] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014bb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02976] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014bc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02978] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014bd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0297a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014be] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0297c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014bf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0297e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014c0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02980] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014c1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02982] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014c2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02984] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014c3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02986] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014c4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02988] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014c5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0298a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014c6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0298c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014c7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0298e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014c8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02990] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014c9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02992] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014ca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02994] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014cb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02996] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014cc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02998] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014cd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0299a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014ce] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0299c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014cf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0299e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014d0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014d1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014d2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014d3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014d4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014d5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014d6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014d7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014d8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014d9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014da] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014db] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014dc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014dd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014de] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014df] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014e0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014e1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014e2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014e3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014e4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014e5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014e6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014e7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014e8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014e9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014ea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014eb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014ec] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014ed] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014ee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014ef] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014f0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014f1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014f2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014f3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014f4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014f5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014f6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014f7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014f8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014f9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014fa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014fb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014fc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014fd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014fe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014ff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h029fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01500] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a00] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01501] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a02] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01502] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a04] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01503] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a06] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01504] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a08] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01505] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a0a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01506] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a0c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01507] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a0e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01508] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a10] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01509] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a12] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0150a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a14] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0150b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a16] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0150c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a18] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0150d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a1a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0150e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a1c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0150f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a1e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01510] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a20] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01511] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a22] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01512] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a24] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01513] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a26] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01514] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a28] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01515] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a2a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01516] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a2c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01517] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a2e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01518] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a30] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01519] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a32] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0151a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a34] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0151b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a36] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0151c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a38] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0151d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a3a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0151e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a3c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0151f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a3e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01520] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a40] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01521] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a42] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01522] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a44] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01523] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a46] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01524] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a48] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01525] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a4a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01526] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a4c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01527] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a4e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01528] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a50] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01529] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a52] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0152a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a54] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0152b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a56] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0152c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a58] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0152d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a5a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0152e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a5c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0152f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a5e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01530] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a60] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01531] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a62] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01532] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a64] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01533] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a66] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01534] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a68] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01535] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a6a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01536] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a6c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01537] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a6e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01538] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a70] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01539] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a72] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0153a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a74] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0153b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a76] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0153c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a78] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0153d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a7a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0153e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a7c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0153f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a7e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01540] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a80] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01541] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a82] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01542] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a84] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01543] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a86] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01544] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a88] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01545] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a8a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01546] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a8c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01547] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a8e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01548] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a90] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01549] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a92] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0154a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a94] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0154b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a96] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0154c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a98] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0154d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a9a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0154e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a9c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0154f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02a9e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01550] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aa0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01551] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aa2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01552] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aa4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01553] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aa6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01554] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aa8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01555] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aaa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01556] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01557] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01558] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ab0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01559] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ab2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0155a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ab4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0155b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ab6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0155c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ab8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0155d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0155e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02abc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0155f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02abe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01560] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ac0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01561] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ac2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01562] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ac4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01563] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ac6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01564] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ac8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01565] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01566] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02acc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01567] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ace] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01568] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ad0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01569] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ad2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0156a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ad4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0156b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ad6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0156c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ad8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0156d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ada] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0156e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02adc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0156f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ade] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01570] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ae0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01571] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ae2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01572] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ae4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01573] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ae6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01574] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ae8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01575] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01576] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01577] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02aee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01578] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02af0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01579] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02af2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0157a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02af4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0157b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02af6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0157c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02af8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0157d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02afa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0157e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02afc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0157f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02afe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01580] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b00] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01581] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b02] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01582] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b04] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01583] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b06] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01584] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b08] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01585] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b0a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01586] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b0c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01587] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b0e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01588] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b10] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01589] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b12] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0158a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b14] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0158b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b16] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0158c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b18] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0158d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b1a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0158e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b1c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0158f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b1e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01590] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b20] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01591] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b22] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01592] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b24] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01593] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b26] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01594] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b28] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01595] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b2a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01596] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b2c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01597] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b2e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01598] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b30] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01599] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b32] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0159a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b34] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0159b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b36] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0159c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b38] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0159d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b3a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0159e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b3c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0159f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b3e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015a0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b40] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015a1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b42] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015a2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b44] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015a3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b46] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015a4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b48] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015a5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b4a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015a6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b4c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015a7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b4e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015a8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b50] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015a9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b52] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015aa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b54] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015ab] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b56] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015ac] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b58] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015ad] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b5a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015ae] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b5c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015af] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b5e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015b0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b60] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015b1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b62] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015b2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b64] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015b3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b66] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015b4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b68] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015b5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b6a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015b6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b6c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015b7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b6e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015b8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b70] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015b9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b72] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015ba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b74] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015bb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b76] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015bc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b78] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015bd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b7a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015be] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b7c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015bf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b7e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015c0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b80] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015c1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b82] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015c2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b84] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015c3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b86] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015c4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b88] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015c5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b8a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015c6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b8c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015c7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b8e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015c8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b90] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015c9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b92] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015ca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b94] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015cb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b96] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015cc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b98] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015cd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b9a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015ce] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b9c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015cf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02b9e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015d0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ba0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015d1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ba2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015d2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ba4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015d3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ba6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015d4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ba8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015d5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02baa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015d6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015d7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015d8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bb0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015d9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bb2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015da] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bb4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015db] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bb6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015dc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bb8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015dd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015de] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bbc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015df] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bbe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015e0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bc0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015e1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bc2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015e2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bc4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015e3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bc6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015e4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bc8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015e5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015e6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bcc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015e7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015e8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bd0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015e9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bd2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015ea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bd4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015eb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bd6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015ec] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bd8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015ed] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bda] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015ee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bdc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015ef] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bde] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015f0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02be0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015f1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02be2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015f2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02be4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015f3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02be6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015f4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02be8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015f5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015f6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015f7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015f8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bf0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015f9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bf2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015fa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bf4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015fb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bf6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015fc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bf8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015fd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bfa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015fe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bfc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015ff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02bfe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01600] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c00] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01601] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c02] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01602] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c04] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01603] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c06] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01604] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c08] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01605] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c0a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01606] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c0c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01607] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c0e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01608] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c10] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01609] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c12] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0160a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c14] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0160b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c16] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0160c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c18] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0160d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c1a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0160e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c1c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0160f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c1e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01610] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c20] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01611] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c22] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01612] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c24] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01613] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c26] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01614] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c28] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01615] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c2a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01616] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c2c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01617] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c2e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01618] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c30] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01619] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c32] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0161a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c34] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0161b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c36] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0161c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c38] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0161d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c3a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0161e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c3c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0161f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c3e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01620] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c40] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01621] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c42] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01622] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c44] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01623] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c46] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01624] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c48] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01625] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c4a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01626] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c4c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01627] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c4e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01628] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c50] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01629] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c52] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0162a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c54] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0162b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c56] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0162c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c58] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0162d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c5a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0162e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c5c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0162f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c5e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01630] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c60] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01631] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c62] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01632] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c64] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01633] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c66] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01634] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c68] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01635] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c6a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01636] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c6c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01637] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c6e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01638] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c70] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01639] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c72] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0163a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c74] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0163b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c76] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0163c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c78] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0163d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c7a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0163e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c7c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0163f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c7e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01640] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c80] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01641] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c82] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01642] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c84] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01643] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c86] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01644] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c88] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01645] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c8a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01646] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c8c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01647] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c8e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01648] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c90] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01649] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c92] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0164a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c94] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0164b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c96] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0164c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c98] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0164d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c9a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0164e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c9c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0164f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02c9e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01650] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ca0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01651] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ca2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01652] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ca4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01653] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ca6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01654] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ca8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01655] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02caa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01656] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01657] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01658] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cb0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01659] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cb2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0165a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cb4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0165b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cb6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0165c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cb8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0165d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0165e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cbc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0165f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cbe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01660] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cc0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01661] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cc2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01662] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cc4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01663] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cc6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01664] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cc8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01665] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01666] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ccc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01667] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01668] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cd0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01669] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cd2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0166a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cd4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0166b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cd6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0166c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cd8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0166d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cda] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0166e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cdc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0166f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cde] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01670] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ce0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01671] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ce2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01672] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ce4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01673] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ce6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01674] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ce8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01675] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01676] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01677] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01678] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cf0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01679] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cf2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0167a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cf4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0167b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cf6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0167c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cf8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0167d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cfa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0167e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cfc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0167f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02cfe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01680] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d00] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01681] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d02] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01682] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d04] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01683] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d06] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01684] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d08] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01685] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d0a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01686] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d0c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01687] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d0e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01688] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d10] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01689] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d12] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0168a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d14] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0168b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d16] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0168c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d18] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0168d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d1a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0168e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d1c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0168f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d1e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01690] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d20] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01691] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d22] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01692] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d24] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01693] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d26] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01694] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d28] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01695] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d2a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01696] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d2c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01697] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d2e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01698] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d30] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01699] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d32] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0169a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d34] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0169b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d36] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0169c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d38] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0169d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d3a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0169e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d3c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0169f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d3e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016a0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d40] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016a1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d42] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016a2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d44] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016a3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d46] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016a4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d48] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016a5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d4a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016a6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d4c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016a7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d4e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016a8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d50] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016a9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d52] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016aa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d54] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016ab] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d56] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016ac] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d58] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016ad] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d5a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016ae] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d5c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016af] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d5e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016b0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d60] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016b1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d62] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016b2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d64] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016b3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d66] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016b4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d68] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016b5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d6a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016b6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d6c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016b7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d6e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016b8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d70] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016b9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d72] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016ba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d74] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016bb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d76] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016bc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d78] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016bd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d7a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016be] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d7c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016bf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d7e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016c0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d80] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016c1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d82] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016c2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d84] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016c3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d86] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016c4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d88] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016c5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d8a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016c6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d8c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016c7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d8e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016c8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d90] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016c9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d92] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016ca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d94] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016cb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d96] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016cc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d98] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016cd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d9a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016ce] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d9c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016cf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02d9e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016d0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02da0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016d1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02da2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016d2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02da4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016d3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02da6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016d4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02da8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016d5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02daa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016d6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016d7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016d8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02db0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016d9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02db2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016da] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02db4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016db] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02db6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016dc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02db8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016dd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016de] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dbc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016df] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dbe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016e0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dc0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016e1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dc2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016e2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dc4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016e3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dc6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016e4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dc8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016e5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016e6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dcc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016e7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016e8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dd0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016e9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dd2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016ea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dd4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016eb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dd6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016ec] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dd8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016ed] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dda] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016ee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ddc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016ef] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dde] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016f0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02de0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016f1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02de2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016f2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02de4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016f3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02de6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016f4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02de8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016f5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016f6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016f7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016f8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02df0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016f9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02df2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016fa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02df4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016fb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02df6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016fc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02df8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016fd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dfa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016fe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dfc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016ff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02dfe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01700] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e00] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01701] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e02] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01702] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e04] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01703] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e06] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01704] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e08] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01705] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e0a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01706] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e0c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01707] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e0e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01708] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e10] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01709] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e12] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0170a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e14] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0170b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e16] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0170c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e18] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0170d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e1a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0170e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e1c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0170f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e1e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01710] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e20] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01711] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e22] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01712] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e24] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01713] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e26] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01714] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e28] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01715] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e2a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01716] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e2c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01717] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e2e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01718] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e30] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01719] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e32] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0171a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e34] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0171b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e36] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0171c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e38] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0171d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e3a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0171e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e3c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0171f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e3e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01720] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e40] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01721] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e42] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01722] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e44] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01723] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e46] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01724] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e48] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01725] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e4a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01726] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e4c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01727] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e4e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01728] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e50] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01729] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e52] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0172a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e54] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0172b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e56] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0172c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e58] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0172d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e5a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0172e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e5c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0172f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e5e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01730] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e60] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01731] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e62] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01732] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e64] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01733] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e66] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01734] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e68] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01735] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e6a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01736] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e6c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01737] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e6e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01738] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e70] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01739] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e72] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0173a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e74] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0173b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e76] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0173c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e78] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0173d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e7a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0173e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e7c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0173f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e7e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01740] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e80] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01741] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e82] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01742] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e84] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01743] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e86] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01744] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e88] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01745] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e8a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01746] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e8c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01747] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e8e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01748] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e90] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01749] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e92] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0174a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e94] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0174b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e96] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0174c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e98] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0174d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e9a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0174e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e9c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0174f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02e9e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01750] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ea0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01751] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ea2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01752] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ea4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01753] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ea6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01754] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ea8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01755] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eaa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01756] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01757] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01758] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eb0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01759] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eb2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0175a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eb4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0175b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eb6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0175c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eb8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0175d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0175e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ebc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0175f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ebe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01760] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ec0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01761] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ec2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01762] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ec4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01763] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ec6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01764] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ec8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01765] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01766] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ecc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01767] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ece] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01768] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ed0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01769] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ed2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0176a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ed4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0176b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ed6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0176c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ed8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0176d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eda] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0176e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02edc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0176f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ede] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01770] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ee0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01771] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ee2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01772] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ee4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01773] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ee6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01774] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ee8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01775] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01776] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01777] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02eee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01778] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ef0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01779] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ef2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0177a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ef4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0177b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ef6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0177c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ef8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0177d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02efa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0177e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02efc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0177f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02efe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01780] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f00] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01781] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f02] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01782] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f04] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01783] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f06] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01784] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f08] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01785] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f0a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01786] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f0c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01787] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f0e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01788] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f10] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01789] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f12] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0178a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f14] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0178b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f16] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0178c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f18] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0178d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f1a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0178e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f1c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0178f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f1e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01790] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f20] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01791] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f22] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01792] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f24] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01793] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f26] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01794] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f28] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01795] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f2a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01796] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f2c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01797] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f2e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01798] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f30] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01799] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f32] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0179a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f34] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0179b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f36] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0179c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f38] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0179d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f3a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0179e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f3c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0179f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f3e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017a0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f40] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017a1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f42] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017a2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f44] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017a3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f46] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017a4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f48] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017a5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f4a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017a6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f4c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017a7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f4e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017a8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f50] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017a9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f52] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017aa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f54] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017ab] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f56] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017ac] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f58] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017ad] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f5a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017ae] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f5c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017af] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f5e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017b0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f60] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017b1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f62] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017b2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f64] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017b3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f66] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017b4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f68] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017b5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f6a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017b6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f6c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017b7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f6e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017b8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f70] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017b9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f72] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017ba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f74] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017bb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f76] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017bc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f78] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017bd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f7a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017be] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f7c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017bf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f7e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017c0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f80] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017c1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f82] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017c2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f84] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017c3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f86] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017c4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f88] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017c5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f8a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017c6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f8c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017c7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f8e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017c8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f90] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017c9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f92] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017ca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f94] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017cb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f96] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017cc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f98] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017cd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f9a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017ce] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f9c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017cf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02f9e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017d0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fa0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017d1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fa2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017d2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fa4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017d3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fa6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017d4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fa8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017d5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02faa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017d6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017d7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017d8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fb0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017d9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fb2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017da] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fb4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017db] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fb6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017dc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fb8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017dd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017de] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fbc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017df] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fbe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017e0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fc0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017e1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fc2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017e2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fc4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017e3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fc6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017e4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fc8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017e5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017e6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fcc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017e7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017e8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fd0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017e9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fd2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017ea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fd4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017eb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fd6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017ec] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fd8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017ed] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fda] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017ee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fdc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017ef] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fde] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017f0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fe0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017f1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fe2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017f2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fe4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017f3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fe6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017f4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fe8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017f5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017f6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017f7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02fee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017f8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ff0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017f9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ff2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017fa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ff4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017fb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ff6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017fc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ff8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017fd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ffa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017fe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ffc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017ff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h02ffe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01800] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03000] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01801] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03002] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01802] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03004] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01803] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03006] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01804] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03008] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01805] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0300a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01806] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0300c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01807] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0300e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01808] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03010] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01809] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03012] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0180a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03014] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0180b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03016] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0180c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03018] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0180d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0301a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0180e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0301c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0180f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0301e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01810] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03020] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01811] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03022] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01812] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03024] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01813] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03026] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01814] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03028] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01815] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0302a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01816] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0302c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01817] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0302e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01818] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03030] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01819] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03032] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0181a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03034] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0181b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03036] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0181c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03038] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0181d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0303a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0181e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0303c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0181f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0303e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01820] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03040] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01821] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03042] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01822] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03044] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01823] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03046] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01824] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03048] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01825] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0304a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01826] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0304c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01827] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0304e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01828] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03050] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01829] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03052] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0182a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03054] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0182b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03056] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0182c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03058] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0182d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0305a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0182e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0305c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0182f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0305e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01830] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03060] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01831] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03062] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01832] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03064] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01833] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03066] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01834] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03068] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01835] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0306a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01836] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0306c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01837] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0306e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01838] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03070] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01839] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03072] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0183a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03074] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0183b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03076] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0183c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03078] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0183d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0307a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0183e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0307c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0183f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0307e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01840] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03080] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01841] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03082] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01842] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03084] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01843] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03086] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01844] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03088] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01845] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0308a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01846] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0308c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01847] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0308e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01848] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03090] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01849] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03092] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0184a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03094] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0184b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03096] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0184c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03098] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0184d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0309a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0184e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0309c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0184f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0309e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01850] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01851] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01852] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01853] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01854] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01855] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01856] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01857] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01858] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01859] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0185a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0185b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0185c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0185d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0185e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0185f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01860] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01861] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01862] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01863] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01864] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01865] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01866] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01867] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01868] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01869] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0186a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0186b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0186c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0186d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0186e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0186f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01870] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01871] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01872] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01873] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01874] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01875] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01876] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01877] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01878] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01879] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0187a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0187b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0187c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0187d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0187e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0187f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h030fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01880] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03100] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01881] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03102] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01882] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03104] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01883] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03106] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01884] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03108] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01885] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0310a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01886] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0310c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01887] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0310e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01888] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03110] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01889] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03112] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0188a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03114] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0188b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03116] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0188c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03118] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0188d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0311a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0188e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0311c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0188f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0311e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01890] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03120] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01891] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03122] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01892] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03124] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01893] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03126] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01894] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03128] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01895] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0312a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01896] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0312c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01897] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0312e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01898] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03130] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01899] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03132] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0189a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03134] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0189b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03136] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0189c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03138] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0189d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0313a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0189e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0313c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0189f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0313e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018a0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03140] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018a1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03142] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018a2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03144] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018a3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03146] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018a4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03148] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018a5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0314a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018a6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0314c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018a7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0314e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018a8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03150] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018a9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03152] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018aa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03154] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018ab] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03156] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018ac] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03158] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018ad] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0315a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018ae] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0315c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018af] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0315e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018b0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03160] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018b1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03162] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018b2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03164] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018b3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03166] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018b4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03168] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018b5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0316a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018b6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0316c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018b7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0316e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018b8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03170] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018b9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03172] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018ba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03174] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018bb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03176] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018bc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03178] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018bd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0317a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018be] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0317c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018bf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0317e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018c0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03180] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018c1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03182] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018c2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03184] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018c3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03186] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018c4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03188] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018c5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0318a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018c6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0318c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018c7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0318e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018c8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03190] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018c9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03192] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018ca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03194] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018cb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03196] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018cc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03198] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018cd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0319a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018ce] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0319c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018cf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0319e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018d0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018d1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018d2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018d3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018d4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018d5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018d6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018d7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018d8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018d9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018da] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018db] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018dc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018dd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018de] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018df] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018e0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018e1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018e2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018e3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018e4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018e5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018e6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018e7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018e8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018e9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018ea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018eb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018ec] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018ed] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018ee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018ef] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018f0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018f1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018f2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018f3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018f4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018f5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018f6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018f7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018f8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018f9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018fa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018fb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018fc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018fd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018fe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018ff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h031fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01900] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03200] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01901] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03202] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01902] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03204] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01903] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03206] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01904] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03208] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01905] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0320a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01906] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0320c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01907] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0320e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01908] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03210] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01909] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03212] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0190a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03214] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0190b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03216] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0190c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03218] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0190d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0321a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0190e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0321c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0190f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0321e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01910] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03220] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01911] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03222] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01912] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03224] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01913] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03226] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01914] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03228] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01915] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0322a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01916] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0322c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01917] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0322e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01918] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03230] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01919] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03232] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0191a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03234] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0191b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03236] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0191c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03238] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0191d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0323a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0191e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0323c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0191f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0323e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01920] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03240] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01921] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03242] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01922] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03244] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01923] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03246] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01924] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03248] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01925] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0324a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01926] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0324c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01927] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0324e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01928] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03250] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01929] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03252] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0192a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03254] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0192b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03256] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0192c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03258] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0192d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0325a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0192e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0325c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0192f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0325e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01930] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03260] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01931] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03262] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01932] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03264] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01933] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03266] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01934] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03268] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01935] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0326a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01936] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0326c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01937] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0326e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01938] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03270] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01939] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03272] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0193a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03274] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0193b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03276] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0193c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03278] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0193d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0327a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0193e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0327c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0193f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0327e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01940] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03280] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01941] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03282] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01942] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03284] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01943] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03286] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01944] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03288] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01945] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0328a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01946] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0328c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01947] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0328e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01948] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03290] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01949] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03292] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0194a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03294] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0194b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03296] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0194c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03298] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0194d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0329a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0194e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0329c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0194f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0329e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01950] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01951] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01952] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01953] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01954] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01955] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01956] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01957] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01958] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01959] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0195a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0195b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0195c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0195d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0195e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0195f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01960] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01961] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01962] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01963] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01964] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01965] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01966] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01967] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01968] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01969] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0196a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0196b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0196c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0196d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0196e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0196f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01970] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01971] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01972] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01973] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01974] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01975] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01976] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01977] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01978] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01979] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0197a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0197b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0197c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0197d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0197e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0197f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h032fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01980] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03300] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01981] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03302] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01982] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03304] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01983] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03306] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01984] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03308] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01985] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0330a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01986] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0330c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01987] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0330e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01988] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03310] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01989] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03312] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0198a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03314] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0198b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03316] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0198c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03318] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0198d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0331a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0198e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0331c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0198f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0331e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01990] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03320] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01991] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03322] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01992] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03324] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01993] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03326] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01994] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03328] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01995] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0332a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01996] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0332c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01997] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0332e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01998] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03330] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01999] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03332] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0199a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03334] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0199b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03336] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0199c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03338] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0199d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0333a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0199e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0333c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0199f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0333e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019a0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03340] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019a1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03342] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019a2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03344] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019a3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03346] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019a4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03348] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019a5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0334a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019a6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0334c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019a7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0334e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019a8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03350] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019a9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03352] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019aa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03354] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019ab] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03356] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019ac] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03358] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019ad] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0335a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019ae] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0335c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019af] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0335e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019b0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03360] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019b1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03362] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019b2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03364] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019b3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03366] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019b4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03368] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019b5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0336a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019b6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0336c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019b7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0336e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019b8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03370] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019b9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03372] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019ba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03374] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019bb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03376] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019bc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03378] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019bd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0337a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019be] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0337c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019bf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0337e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019c0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03380] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019c1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03382] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019c2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03384] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019c3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03386] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019c4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03388] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019c5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0338a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019c6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0338c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019c7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0338e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019c8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03390] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019c9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03392] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019ca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03394] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019cb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03396] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019cc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03398] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019cd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0339a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019ce] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0339c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019cf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0339e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019d0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019d1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019d2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019d3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019d4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019d5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019d6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019d7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019d8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019d9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019da] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019db] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019dc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019dd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019de] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019df] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019e0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019e1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019e2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019e3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019e4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019e5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019e6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019e7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019e8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019e9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019ea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019eb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019ec] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019ed] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019ee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019ef] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019f0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019f1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019f2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019f3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019f4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019f5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019f6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019f7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019f8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019f9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019fa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019fb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019fc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019fd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019fe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019ff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h033fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a00] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03400] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a01] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03402] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a02] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03404] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a03] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03406] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a04] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03408] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a05] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0340a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a06] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0340c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a07] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0340e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a08] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03410] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a09] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03412] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a0a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03414] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a0b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03416] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a0c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03418] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a0d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0341a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a0e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0341c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a0f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0341e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a10] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03420] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a11] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03422] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a12] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03424] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a13] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03426] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a14] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03428] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a15] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0342a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a16] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0342c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a17] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0342e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a18] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03430] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a19] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03432] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a1a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03434] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a1b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03436] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a1c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03438] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a1d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0343a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a1e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0343c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a1f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0343e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a20] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03440] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a21] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03442] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a22] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03444] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a23] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03446] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a24] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03448] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a25] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0344a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a26] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0344c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a27] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0344e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a28] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03450] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a29] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03452] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a2a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03454] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a2b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03456] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a2c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03458] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a2d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0345a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a2e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0345c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a2f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0345e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a30] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03460] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a31] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03462] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a32] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03464] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a33] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03466] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a34] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03468] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a35] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0346a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a36] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0346c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a37] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0346e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a38] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03470] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a39] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03472] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a3a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03474] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a3b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03476] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a3c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03478] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a3d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0347a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a3e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0347c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a3f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0347e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a40] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03480] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a41] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03482] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a42] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03484] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a43] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03486] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a44] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03488] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a45] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0348a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a46] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0348c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a47] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0348e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a48] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03490] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a49] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03492] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a4a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03494] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a4b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03496] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a4c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03498] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a4d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0349a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a4e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0349c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a4f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0349e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a50] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a51] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a52] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a53] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a54] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a55] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a56] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a57] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a58] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a59] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a5a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a5b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a5c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a5d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a5e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a5f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a60] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a61] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a62] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a63] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a64] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a65] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a66] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a67] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a68] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a69] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a6a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a6b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a6c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a6d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a6e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a6f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a70] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a71] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a72] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a73] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a74] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a75] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a76] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a77] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a78] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a79] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a7a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a7b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a7c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a7d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a7e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a7f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h034fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a80] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03500] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a81] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03502] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a82] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03504] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a83] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03506] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a84] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03508] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a85] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0350a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a86] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0350c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a87] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0350e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a88] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03510] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a89] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03512] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a8a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03514] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a8b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03516] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a8c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03518] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a8d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0351a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a8e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0351c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a8f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0351e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a90] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03520] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a91] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03522] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a92] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03524] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a93] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03526] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a94] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03528] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a95] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0352a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a96] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0352c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a97] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0352e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a98] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03530] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a99] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03532] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a9a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03534] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a9b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03536] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a9c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03538] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a9d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0353a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a9e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0353c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a9f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0353e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aa0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03540] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aa1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03542] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aa2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03544] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aa3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03546] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aa4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03548] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aa5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0354a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aa6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0354c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aa7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0354e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aa8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03550] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aa9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03552] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aaa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03554] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aab] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03556] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aac] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03558] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aad] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0355a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aae] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0355c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aaf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0355e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ab0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03560] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ab1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03562] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ab2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03564] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ab3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03566] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ab4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03568] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ab5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0356a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ab6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0356c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ab7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0356e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ab8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03570] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ab9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03572] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03574] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01abb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03576] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01abc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03578] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01abd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0357a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01abe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0357c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01abf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0357e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ac0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03580] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ac1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03582] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ac2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03584] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ac3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03586] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ac4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03588] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ac5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0358a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ac6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0358c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ac7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0358e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ac8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03590] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ac9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03592] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03594] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01acb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03596] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01acc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03598] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01acd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0359a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ace] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0359c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01acf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0359e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ad0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ad1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ad2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ad3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ad4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ad5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ad6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ad7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ad8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ad9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ada] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01adb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01adc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01add] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ade] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01adf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ae0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ae1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ae2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ae3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ae4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ae5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ae6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ae7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ae8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ae9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aeb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aec] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aed] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aef] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01af0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01af1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01af2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01af3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01af4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01af5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01af6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01af7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01af8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01af9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01afa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01afb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01afc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01afd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01afe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h035fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b00] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03600] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b01] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03602] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b02] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03604] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b03] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03606] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b04] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03608] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b05] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0360a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b06] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0360c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b07] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0360e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b08] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03610] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b09] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03612] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b0a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03614] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b0b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03616] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b0c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03618] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b0d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0361a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b0e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0361c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b0f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0361e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b10] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03620] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b11] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03622] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b12] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03624] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b13] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03626] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b14] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03628] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b15] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0362a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b16] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0362c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b17] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0362e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b18] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03630] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b19] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03632] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b1a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03634] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b1b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03636] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b1c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03638] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b1d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0363a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b1e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0363c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b1f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0363e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b20] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03640] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b21] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03642] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b22] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03644] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b23] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03646] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b24] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03648] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b25] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0364a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b26] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0364c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b27] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0364e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b28] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03650] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b29] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03652] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b2a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03654] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b2b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03656] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b2c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03658] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b2d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0365a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b2e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0365c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b2f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0365e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b30] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03660] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b31] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03662] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b32] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03664] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b33] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03666] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b34] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03668] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b35] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0366a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b36] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0366c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b37] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0366e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b38] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03670] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b39] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03672] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b3a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03674] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b3b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03676] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b3c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03678] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b3d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0367a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b3e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0367c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b3f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0367e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b40] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03680] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b41] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03682] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b42] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03684] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b43] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03686] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b44] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03688] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b45] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0368a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b46] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0368c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b47] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0368e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b48] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03690] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b49] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03692] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b4a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03694] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b4b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03696] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b4c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03698] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b4d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0369a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b4e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0369c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b4f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0369e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b50] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b51] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b52] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b53] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b54] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b55] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b56] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b57] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b58] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b59] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b5a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b5b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b5c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b5d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b5e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b5f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b60] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b61] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b62] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b63] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b64] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b65] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b66] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b67] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b68] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b69] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b6a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b6b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b6c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b6d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b6e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b6f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b70] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b71] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b72] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b73] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b74] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b75] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b76] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b77] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b78] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b79] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b7a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b7b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b7c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b7d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b7e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b7f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h036fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b80] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03700] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b81] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03702] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b82] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03704] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b83] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03706] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b84] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03708] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b85] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0370a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b86] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0370c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b87] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0370e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b88] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03710] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b89] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03712] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b8a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03714] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b8b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03716] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b8c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03718] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b8d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0371a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b8e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0371c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b8f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0371e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b90] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03720] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b91] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03722] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b92] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03724] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b93] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03726] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b94] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03728] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b95] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0372a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b96] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0372c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b97] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0372e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b98] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03730] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b99] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03732] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b9a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03734] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b9b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03736] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b9c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03738] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b9d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0373a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b9e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0373c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b9f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0373e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ba0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03740] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ba1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03742] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ba2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03744] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ba3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03746] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ba4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03748] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ba5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0374a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ba6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0374c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ba7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0374e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ba8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03750] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ba9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03752] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01baa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03754] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bab] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03756] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bac] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03758] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bad] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0375a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bae] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0375c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01baf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0375e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bb0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03760] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bb1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03762] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bb2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03764] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bb3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03766] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bb4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03768] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bb5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0376a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bb6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0376c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bb7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0376e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bb8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03770] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bb9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03772] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03774] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bbb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03776] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bbc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03778] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bbd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0377a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bbe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0377c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bbf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0377e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bc0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03780] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bc1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03782] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bc2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03784] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bc3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03786] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bc4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03788] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bc5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0378a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bc6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0378c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bc7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0378e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bc8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03790] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bc9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03792] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03794] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bcb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03796] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bcc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03798] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bcd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0379a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bce] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0379c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bcf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0379e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bd0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bd1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bd2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bd3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bd4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bd5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bd6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bd7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bd8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bd9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bda] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bdb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bdc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bdd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bde] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bdf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01be0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01be1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01be2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01be3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01be4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01be5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01be6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01be7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01be8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01be9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01beb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bec] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bed] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bef] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bf0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bf1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bf2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bf3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bf4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bf5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bf6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bf7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bf8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bf9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bfa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bfb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bfc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bfd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bfe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h037fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c00] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03800] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c01] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03802] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c02] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03804] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c03] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03806] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c04] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03808] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c05] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0380a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c06] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0380c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c07] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0380e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c08] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03810] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c09] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03812] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c0a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03814] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c0b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03816] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c0c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03818] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c0d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0381a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c0e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0381c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c0f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0381e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c10] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03820] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c11] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03822] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c12] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03824] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c13] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03826] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c14] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03828] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c15] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0382a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c16] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0382c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c17] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0382e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c18] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03830] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c19] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03832] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c1a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03834] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c1b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03836] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c1c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03838] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c1d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0383a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c1e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0383c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c1f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0383e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c20] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03840] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c21] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03842] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c22] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03844] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c23] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03846] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c24] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03848] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c25] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0384a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c26] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0384c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c27] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0384e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c28] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03850] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c29] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03852] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c2a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03854] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c2b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03856] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c2c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03858] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c2d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0385a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c2e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0385c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c2f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0385e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c30] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03860] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c31] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03862] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c32] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03864] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c33] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03866] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c34] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03868] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c35] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0386a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c36] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0386c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c37] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0386e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c38] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03870] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c39] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03872] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c3a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03874] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c3b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03876] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c3c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03878] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c3d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0387a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c3e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0387c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c3f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0387e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c40] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03880] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c41] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03882] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c42] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03884] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c43] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03886] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c44] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03888] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c45] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0388a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c46] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0388c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c47] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0388e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c48] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03890] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c49] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03892] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c4a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03894] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c4b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03896] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c4c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03898] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c4d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0389a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c4e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0389c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c4f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0389e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c50] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c51] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c52] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c53] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c54] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c55] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c56] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c57] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c58] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c59] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c5a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c5b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c5c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c5d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c5e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c5f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c60] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c61] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c62] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c63] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c64] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c65] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c66] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c67] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c68] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c69] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c6a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c6b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c6c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c6d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c6e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c6f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c70] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c71] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c72] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c73] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c74] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c75] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c76] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c77] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c78] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c79] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c7a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c7b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c7c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c7d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c7e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c7f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h038fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c80] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03900] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c81] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03902] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c82] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03904] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c83] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03906] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c84] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03908] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c85] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0390a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c86] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0390c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c87] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0390e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c88] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03910] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c89] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03912] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c8a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03914] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c8b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03916] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c8c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03918] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c8d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0391a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c8e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0391c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c8f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0391e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c90] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03920] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c91] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03922] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c92] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03924] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c93] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03926] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c94] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03928] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c95] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0392a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c96] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0392c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c97] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0392e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c98] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03930] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c99] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03932] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c9a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03934] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c9b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03936] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c9c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03938] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c9d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0393a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c9e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0393c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c9f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0393e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ca0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03940] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ca1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03942] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ca2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03944] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ca3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03946] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ca4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03948] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ca5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0394a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ca6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0394c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ca7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0394e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ca8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03950] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ca9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03952] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01caa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03954] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cab] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03956] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cac] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03958] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cad] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0395a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cae] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0395c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01caf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0395e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cb0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03960] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cb1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03962] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cb2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03964] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cb3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03966] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cb4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03968] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cb5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0396a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cb6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0396c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cb7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0396e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cb8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03970] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cb9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03972] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03974] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cbb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03976] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cbc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03978] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cbd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0397a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cbe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0397c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cbf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0397e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cc0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03980] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cc1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03982] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cc2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03984] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cc3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03986] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cc4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03988] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cc5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0398a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cc6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0398c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cc7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0398e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cc8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03990] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cc9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03992] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03994] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ccb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03996] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ccc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03998] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ccd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0399a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cce] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0399c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ccf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h0399e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cd0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039a0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cd1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039a2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cd2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039a4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cd3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039a6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cd4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039a8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cd5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039aa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cd6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039ac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cd7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039ae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cd8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039b0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cd9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039b2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cda] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039b4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cdb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039b6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cdc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039b8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cdd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039ba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cde] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039bc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cdf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039be] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ce0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039c0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ce1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039c2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ce2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039c4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ce3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039c6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ce4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039c8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ce5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039ca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ce6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039cc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ce7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039ce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ce8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039d0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ce9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039d2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039d4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ceb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039d6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cec] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039d8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ced] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039da] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039dc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cef] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039de] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cf0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039e0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cf1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039e2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cf2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039e4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cf3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039e6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cf4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039e8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cf5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039ea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cf6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039ec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cf7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039ee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cf8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039f0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cf9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039f2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cfa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039f4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cfb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039f6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cfc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039f8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cfd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039fa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cfe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039fc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h039fe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d00] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a00] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d01] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a02] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d02] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a04] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d03] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a06] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d04] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a08] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d05] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a0a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d06] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a0c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d07] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a0e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d08] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a10] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d09] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a12] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d0a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a14] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d0b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a16] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d0c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a18] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d0d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a1a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d0e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a1c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d0f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a1e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d10] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a20] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d11] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a22] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d12] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a24] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d13] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a26] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d14] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a28] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d15] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a2a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d16] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a2c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d17] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a2e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d18] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a30] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d19] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a32] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d1a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a34] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d1b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a36] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d1c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a38] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d1d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a3a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d1e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a3c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d1f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a3e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d20] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a40] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d21] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a42] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d22] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a44] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d23] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a46] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d24] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a48] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d25] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a4a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d26] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a4c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d27] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a4e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d28] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a50] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d29] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a52] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d2a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a54] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d2b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a56] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d2c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a58] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d2d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a5a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d2e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a5c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d2f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a5e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d30] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a60] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d31] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a62] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d32] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a64] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d33] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a66] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d34] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a68] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d35] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a6a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d36] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a6c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d37] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a6e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d38] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a70] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d39] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a72] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d3a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a74] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d3b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a76] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d3c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a78] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d3d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a7a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d3e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a7c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d3f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a7e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d40] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a80] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d41] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a82] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d42] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a84] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d43] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a86] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d44] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a88] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d45] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a8a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d46] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a8c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d47] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a8e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d48] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a90] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d49] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a92] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d4a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a94] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d4b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a96] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d4c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a98] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d4d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a9a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d4e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a9c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d4f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03a9e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d50] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aa0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d51] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aa2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d52] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aa4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d53] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aa6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d54] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aa8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d55] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aaa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d56] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d57] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d58] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ab0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d59] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ab2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d5a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ab4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d5b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ab6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d5c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ab8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d5d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d5e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03abc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d5f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03abe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d60] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ac0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d61] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ac2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d62] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ac4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d63] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ac6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d64] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ac8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d65] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d66] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03acc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d67] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ace] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d68] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ad0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d69] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ad2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d6a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ad4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d6b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ad6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d6c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ad8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d6d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ada] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d6e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03adc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d6f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ade] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d70] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ae0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d71] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ae2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d72] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ae4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d73] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ae6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d74] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ae8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d75] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d76] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d77] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03aee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d78] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03af0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d79] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03af2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d7a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03af4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d7b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03af6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d7c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03af8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d7d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03afa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d7e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03afc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d7f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03afe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d80] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b00] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d81] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b02] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d82] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b04] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d83] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b06] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d84] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b08] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d85] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b0a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d86] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b0c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d87] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b0e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d88] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b10] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d89] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b12] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d8a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b14] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d8b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b16] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d8c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b18] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d8d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b1a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d8e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b1c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d8f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b1e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d90] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b20] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d91] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b22] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d92] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b24] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d93] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b26] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d94] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b28] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d95] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b2a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d96] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b2c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d97] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b2e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d98] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b30] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d99] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b32] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d9a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b34] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d9b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b36] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d9c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b38] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d9d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b3a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d9e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b3c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d9f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b3e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01da0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b40] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01da1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b42] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01da2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b44] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01da3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b46] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01da4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b48] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01da5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b4a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01da6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b4c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01da7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b4e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01da8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b50] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01da9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b52] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01daa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b54] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dab] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b56] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dac] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b58] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dad] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b5a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dae] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b5c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01daf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b5e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01db0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b60] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01db1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b62] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01db2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b64] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01db3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b66] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01db4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b68] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01db5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b6a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01db6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b6c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01db7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b6e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01db8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b70] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01db9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b72] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b74] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dbb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b76] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dbc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b78] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dbd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b7a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dbe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b7c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dbf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b7e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dc0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b80] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dc1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b82] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dc2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b84] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dc3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b86] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dc4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b88] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dc5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b8a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dc6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b8c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dc7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b8e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dc8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b90] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dc9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b92] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b94] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dcb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b96] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dcc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b98] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dcd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b9a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dce] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b9c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dcf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03b9e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dd0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ba0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dd1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ba2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dd2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ba4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dd3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ba6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dd4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ba8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dd5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03baa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dd6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dd7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dd8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bb0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dd9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bb2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dda] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bb4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ddb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bb6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ddc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bb8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ddd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dde] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bbc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ddf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bbe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01de0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bc0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01de1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bc2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01de2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bc4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01de3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bc6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01de4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bc8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01de5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01de6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bcc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01de7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01de8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bd0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01de9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bd2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bd4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01deb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bd6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dec] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bd8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ded] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bda] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bdc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01def] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bde] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01df0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03be0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01df1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03be2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01df2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03be4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01df3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03be6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01df4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03be8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01df5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01df6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01df7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01df8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bf0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01df9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bf2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dfa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bf4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dfb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bf6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dfc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bf8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dfd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bfa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dfe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bfc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03bfe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e00] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c00] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e01] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c02] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e02] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c04] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e03] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c06] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e04] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c08] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e05] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c0a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e06] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c0c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e07] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c0e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e08] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c10] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e09] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c12] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e0a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c14] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e0b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c16] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e0c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c18] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e0d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c1a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e0e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c1c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e0f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c1e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e10] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c20] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e11] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c22] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e12] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c24] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e13] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c26] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e14] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c28] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e15] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c2a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e16] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c2c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e17] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c2e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e18] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c30] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e19] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c32] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e1a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c34] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e1b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c36] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e1c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c38] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e1d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c3a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e1e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c3c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e1f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c3e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e20] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c40] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e21] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c42] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e22] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c44] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e23] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c46] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e24] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c48] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e25] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c4a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e26] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c4c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e27] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c4e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e28] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c50] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e29] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c52] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e2a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c54] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e2b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c56] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e2c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c58] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e2d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c5a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e2e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c5c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e2f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c5e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e30] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c60] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e31] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c62] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e32] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c64] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e33] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c66] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e34] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c68] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e35] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c6a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e36] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c6c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e37] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c6e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e38] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c70] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e39] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c72] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e3a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c74] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e3b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c76] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e3c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c78] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e3d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c7a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e3e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c7c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e3f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c7e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e40] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c80] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e41] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c82] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e42] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c84] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e43] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c86] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e44] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c88] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e45] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c8a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e46] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c8c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e47] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c8e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e48] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c90] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e49] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c92] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e4a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c94] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e4b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c96] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e4c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c98] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e4d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c9a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e4e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c9c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e4f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03c9e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e50] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ca0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e51] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ca2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e52] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ca4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e53] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ca6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e54] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ca8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e55] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03caa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e56] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e57] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e58] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cb0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e59] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cb2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e5a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cb4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e5b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cb6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e5c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cb8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e5d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e5e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cbc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e5f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cbe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e60] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cc0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e61] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cc2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e62] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cc4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e63] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cc6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e64] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cc8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e65] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e66] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ccc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e67] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e68] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cd0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e69] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cd2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e6a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cd4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e6b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cd6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e6c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cd8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e6d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cda] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e6e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cdc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e6f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cde] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e70] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ce0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e71] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ce2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e72] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ce4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e73] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ce6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e74] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ce8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e75] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e76] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e77] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e78] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cf0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e79] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cf2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e7a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cf4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e7b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cf6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e7c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cf8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e7d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cfa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e7e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cfc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e7f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03cfe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e80] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d00] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e81] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d02] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e82] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d04] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e83] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d06] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e84] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d08] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e85] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d0a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e86] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d0c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e87] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d0e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e88] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d10] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e89] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d12] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e8a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d14] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e8b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d16] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e8c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d18] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e8d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d1a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e8e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d1c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e8f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d1e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e90] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d20] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e91] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d22] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e92] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d24] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e93] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d26] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e94] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d28] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e95] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d2a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e96] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d2c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e97] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d2e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e98] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d30] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e99] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d32] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e9a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d34] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e9b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d36] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e9c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d38] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e9d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d3a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e9e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d3c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e9f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d3e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ea0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d40] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ea1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d42] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ea2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d44] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ea3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d46] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ea4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d48] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ea5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d4a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ea6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d4c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ea7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d4e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ea8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d50] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ea9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d52] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eaa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d54] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eab] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d56] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eac] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d58] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ead] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d5a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eae] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d5c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eaf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d5e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eb0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d60] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eb1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d62] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eb2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d64] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eb3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d66] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eb4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d68] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eb5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d6a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eb6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d6c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eb7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d6e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eb8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d70] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eb9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d72] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d74] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ebb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d76] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ebc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d78] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ebd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d7a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ebe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d7c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ebf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d7e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ec0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d80] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ec1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d82] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ec2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d84] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ec3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d86] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ec4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d88] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ec5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d8a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ec6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d8c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ec7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d8e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ec8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d90] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ec9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d92] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d94] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ecb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d96] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ecc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d98] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ecd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d9a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ece] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d9c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ecf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03d9e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ed0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03da0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ed1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03da2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ed2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03da4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ed3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03da6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ed4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03da8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ed5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03daa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ed6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ed7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ed8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03db0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ed9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03db2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eda] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03db4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01edb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03db6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01edc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03db8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01edd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ede] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dbc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01edf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dbe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ee0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dc0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ee1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dc2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ee2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dc4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ee3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dc6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ee4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dc8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ee5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ee6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dcc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ee7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ee8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dd0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ee9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dd2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dd4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eeb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dd6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eec] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dd8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eed] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dda] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ddc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eef] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dde] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ef0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03de0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ef1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03de2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ef2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03de4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ef3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03de6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ef4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03de8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ef5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ef6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ef7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ef8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03df0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ef9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03df2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01efa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03df4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01efb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03df6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01efc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03df8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01efd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dfa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01efe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dfc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03dfe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f00] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e00] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f01] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e02] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f02] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e04] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f03] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e06] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f04] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e08] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f05] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e0a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f06] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e0c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f07] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e0e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f08] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e10] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f09] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e12] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f0a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e14] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f0b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e16] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f0c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e18] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f0d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e1a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f0e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e1c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f0f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e1e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f10] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e20] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f11] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e22] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f12] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e24] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f13] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e26] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f14] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e28] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f15] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e2a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f16] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e2c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f17] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e2e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f18] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e30] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f19] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e32] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f1a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e34] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f1b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e36] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f1c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e38] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f1d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e3a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f1e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e3c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f1f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e3e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f20] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e40] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f21] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e42] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f22] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e44] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f23] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e46] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f24] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e48] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f25] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e4a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f26] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e4c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f27] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e4e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f28] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e50] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f29] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e52] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f2a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e54] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f2b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e56] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f2c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e58] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f2d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e5a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f2e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e5c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f2f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e5e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f30] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e60] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f31] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e62] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f32] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e64] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f33] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e66] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f34] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e68] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f35] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e6a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f36] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e6c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f37] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e6e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f38] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e70] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f39] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e72] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f3a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e74] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f3b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e76] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f3c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e78] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f3d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e7a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f3e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e7c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f3f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e7e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f40] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e80] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f41] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e82] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f42] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e84] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f43] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e86] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f44] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e88] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f45] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e8a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f46] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e8c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f47] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e8e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f48] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e90] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f49] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e92] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f4a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e94] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f4b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e96] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f4c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e98] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f4d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e9a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f4e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e9c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f4f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03e9e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f50] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ea0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f51] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ea2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f52] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ea4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f53] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ea6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f54] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ea8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f55] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eaa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f56] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f57] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f58] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eb0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f59] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eb2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f5a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eb4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f5b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eb6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f5c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eb8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f5d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f5e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ebc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f5f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ebe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f60] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ec0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f61] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ec2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f62] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ec4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f63] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ec6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f64] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ec8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f65] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f66] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ecc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f67] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ece] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f68] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ed0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f69] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ed2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f6a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ed4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f6b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ed6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f6c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ed8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f6d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eda] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f6e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03edc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f6f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ede] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f70] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ee0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f71] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ee2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f72] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ee4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f73] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ee6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f74] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ee8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f75] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f76] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f77] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03eee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f78] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ef0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f79] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ef2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f7a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ef4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f7b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ef6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f7c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ef8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f7d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03efa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f7e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03efc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f7f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03efe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f80] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f00] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f81] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f02] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f82] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f04] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f83] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f06] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f84] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f08] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f85] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f0a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f86] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f0c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f87] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f0e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f88] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f10] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f89] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f12] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f8a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f14] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f8b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f16] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f8c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f18] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f8d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f1a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f8e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f1c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f8f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f1e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f90] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f20] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f91] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f22] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f92] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f24] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f93] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f26] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f94] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f28] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f95] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f2a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f96] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f2c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f97] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f2e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f98] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f30] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f99] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f32] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f9a] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f34] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f9b] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f36] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f9c] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f38] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f9d] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f3a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f9e] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f3c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f9f] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f3e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fa0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f40] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fa1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f42] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fa2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f44] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fa3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f46] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fa4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f48] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fa5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f4a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fa6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f4c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fa7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f4e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fa8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f50] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fa9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f52] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01faa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f54] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fab] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f56] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fac] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f58] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fad] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f5a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fae] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f5c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01faf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f5e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fb0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f60] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fb1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f62] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fb2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f64] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fb3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f66] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fb4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f68] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fb5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f6a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fb6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f6c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fb7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f6e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fb8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f70] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fb9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f72] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fba] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f74] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fbb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f76] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fbc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f78] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fbd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f7a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fbe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f7c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fbf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f7e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fc0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f80] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fc1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f82] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fc2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f84] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fc3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f86] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fc4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f88] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fc5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f8a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fc6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f8c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fc7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f8e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fc8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f90] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fc9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f92] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fca] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f94] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fcb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f96] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fcc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f98] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fcd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f9a] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fce] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f9c] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fcf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03f9e] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fd0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fa0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fd1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fa2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fd2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fa4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fd3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fa6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fd4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fa8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fd5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03faa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fd6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fac] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fd7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fae] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fd8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fb0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fd9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fb2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fda] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fb4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fdb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fb6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fdc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fb8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fdd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fba] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fde] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fbc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fdf] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fbe] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fe0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fc0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fe1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fc2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fe2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fc4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fe3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fc6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fe4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fc8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fe5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fca] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fe6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fcc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fe7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fce] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fe8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fd0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fe9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fd2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fea] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fd4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01feb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fd6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fec] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fd8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fed] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fda] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fee] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fdc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fef] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fde] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ff0] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fe0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ff1] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fe2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ff2] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fe4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ff3] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fe6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ff4] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fe8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ff5] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fea] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ff6] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fec] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ff7] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03fee] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ff8] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ff0] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ff9] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ff2] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ffa] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ff4] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ffb] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ff6] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ffc] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ff8] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ffd] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ffa] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ffe] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ffc] ;
//end
//always_comb begin // 
               Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fff] =  Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b['h03ffe] ;
//end
