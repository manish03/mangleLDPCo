//`include "GF2_LDPC_fgallag_0x00007_assign_inc.sv"
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00000] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00000] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00001] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00001] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00002] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00003] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00002] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00004] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00005] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00003] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00006] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00007] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00004] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00008] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00009] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00005] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0000a] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0000b] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00006] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0000c] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0000d] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00007] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0000e] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0000f] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00008] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00010] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00011] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00009] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00012] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00013] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0000a] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00014] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00015] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0000b] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00016] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00017] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0000c] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00018] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00019] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0000d] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0001a] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0001b] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0000e] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0001c] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0001d] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0000f] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0001e] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0001f] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00010] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00020] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00021] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00011] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00022] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00023] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00012] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00024] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00025] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00013] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00026] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00027] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00014] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00028] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00029] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00015] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0002a] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0002b] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00016] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0002c] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0002d] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00017] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0002e] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0002f] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00018] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00030] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00031] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00019] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00032] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00033] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0001a] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00034] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00035] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0001b] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00036] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00037] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0001c] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00038] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00039] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0001d] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0003a] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0003b] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0001e] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0003c] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0003d] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0001f] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0003e] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0003f] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00020] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00040] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00041] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00021] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00042] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00043] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00022] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00044] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00045] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00023] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00046] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00047] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00024] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00048] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00049] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00025] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0004a] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0004b] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00026] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0004c] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0004d] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00027] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0004e] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0004f] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00028] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00050] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00051] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00029] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00052] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00053] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0002a] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00054] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00055] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0002b] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00056] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00057] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0002c] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00058] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00059] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0002d] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0005a] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0005b] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0002e] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0005c] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0005d] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0002f] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0005e] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0005f] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00030] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00060] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00061] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00031] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00062] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00063] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00032] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00064] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00065] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00033] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00066] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00067] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00034] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00068] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00069] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00035] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0006a] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00036] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0006c] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0006d] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00037] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0006e] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00038] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00070] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00071] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00039] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00072] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0003a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00074] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0003b] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00076] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00077] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0003c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00078] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0003d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0007a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0003e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0007c] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0003f] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0007e] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h0007f] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00040] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00080] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00041] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00082] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00042] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00084] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00043] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00086] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00044] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00088] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00045] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0008a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00046] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0008c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00047] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0008e] ;
//end
//always_comb begin
              Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00048] = 
          (!fgallag_sel['h00007]) ? 
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00090] : //%
                       Ic8a4ab93493bd6cdd4939054e46d2247['h00091] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00049] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00092] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0004a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00094] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0004b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00096] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0004c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00098] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0004d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0009a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0004e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0009c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0004f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0009e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00050] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000a0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00051] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000a2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00052] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000a4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00053] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000a6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00054] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000a8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00055] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000aa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00056] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000ac] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00057] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000ae] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00058] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000b0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00059] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000b2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0005a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000b4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0005b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000b6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0005c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000b8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0005d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000ba] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0005e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000bc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0005f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000be] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00060] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000c0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00061] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000c2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00062] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000c4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00063] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000c6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00064] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000c8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00065] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000ca] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00066] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000cc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00067] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000ce] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00068] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000d0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00069] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000d2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0006a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000d4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0006b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000d6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0006c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000d8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0006d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000da] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0006e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000dc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0006f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000de] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00070] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000e0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00071] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000e2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00072] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000e4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00073] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000e6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00074] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000e8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00075] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000ea] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00076] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000ec] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00077] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000ee] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00078] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000f0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00079] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000f2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0007a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000f4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0007b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000f6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0007c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000f8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0007d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000fa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0007e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000fc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0007f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h000fe] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00080] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00100] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00081] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00102] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00082] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00104] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00083] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00106] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00084] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00108] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00085] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0010a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00086] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0010c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00087] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0010e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00088] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00110] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00089] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00112] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0008a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00114] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0008b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00116] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0008c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00118] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0008d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0011a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0008e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0011c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0008f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0011e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00090] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00120] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00091] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00122] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00092] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00124] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00093] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00126] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00094] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00128] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00095] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0012a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00096] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0012c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00097] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0012e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00098] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00130] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00099] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00132] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0009a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00134] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0009b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00136] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0009c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00138] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0009d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0013a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0009e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0013c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0009f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0013e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000a0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00140] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000a1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00142] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000a2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00144] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000a3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00146] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000a4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00148] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000a5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0014a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000a6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0014c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000a7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0014e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000a8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00150] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000a9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00152] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000aa] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00154] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000ab] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00156] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000ac] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00158] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000ad] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0015a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000ae] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0015c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000af] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0015e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000b0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00160] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000b1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00162] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000b2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00164] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000b3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00166] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000b4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00168] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000b5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0016a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000b6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0016c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000b7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0016e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000b8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00170] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000b9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00172] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000ba] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00174] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000bb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00176] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000bc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00178] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000bd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0017a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000be] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0017c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000bf] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0017e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000c0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00180] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000c1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00182] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000c2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00184] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000c3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00186] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000c4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00188] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000c5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0018a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000c6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0018c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000c7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0018e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000c8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00190] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000c9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00192] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000ca] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00194] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000cb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00196] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000cc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00198] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000cd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0019a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000ce] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0019c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000cf] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0019e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000d0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001a0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000d1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001a2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000d2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001a4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000d3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001a6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000d4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001a8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000d5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001aa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000d6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001ac] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000d7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001ae] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000d8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001b0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000d9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001b2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000da] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001b4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000db] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001b6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000dc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001b8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000dd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001ba] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000de] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001bc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000df] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001be] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000e0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001c0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000e1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001c2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000e2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001c4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000e3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001c6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000e4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001c8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000e5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001ca] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000e6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001cc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000e7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001ce] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000e8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001d0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000e9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001d2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000ea] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001d4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000eb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001d6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000ec] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001d8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000ed] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001da] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000ee] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001dc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000ef] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001de] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000f0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001e0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000f1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001e2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000f2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001e4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000f3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001e6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000f4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001e8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000f5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001ea] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000f6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001ec] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000f7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001ee] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000f8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001f0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000f9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001f2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000fa] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001f4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000fb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001f6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000fc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001f8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000fd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001fa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000fe] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001fc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h000ff] =  Ic8a4ab93493bd6cdd4939054e46d2247['h001fe] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00100] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00200] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00101] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00202] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00102] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00204] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00103] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00206] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00104] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00208] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00105] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0020a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00106] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0020c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00107] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0020e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00108] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00210] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00109] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00212] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0010a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00214] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0010b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00216] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0010c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00218] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0010d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0021a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0010e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0021c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0010f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0021e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00110] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00220] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00111] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00222] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00112] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00224] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00113] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00226] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00114] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00228] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00115] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0022a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00116] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0022c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00117] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0022e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00118] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00230] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00119] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00232] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0011a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00234] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0011b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00236] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0011c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00238] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0011d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0023a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0011e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0023c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0011f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0023e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00120] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00240] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00121] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00242] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00122] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00244] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00123] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00246] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00124] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00248] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00125] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0024a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00126] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0024c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00127] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0024e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00128] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00250] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00129] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00252] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0012a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00254] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0012b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00256] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0012c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00258] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0012d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0025a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0012e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0025c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0012f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0025e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00130] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00260] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00131] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00262] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00132] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00264] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00133] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00266] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00134] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00268] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00135] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0026a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00136] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0026c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00137] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0026e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00138] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00270] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00139] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00272] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0013a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00274] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0013b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00276] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0013c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00278] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0013d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0027a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0013e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0027c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0013f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0027e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00140] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00280] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00141] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00282] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00142] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00284] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00143] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00286] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00144] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00288] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00145] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0028a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00146] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0028c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00147] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0028e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00148] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00290] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00149] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00292] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0014a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00294] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0014b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00296] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0014c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00298] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0014d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0029a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0014e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0029c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0014f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0029e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00150] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002a0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00151] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002a2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00152] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002a4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00153] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002a6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00154] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002a8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00155] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002aa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00156] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002ac] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00157] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002ae] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00158] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002b0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00159] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002b2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0015a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002b4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0015b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002b6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0015c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002b8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0015d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002ba] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0015e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002bc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0015f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002be] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00160] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002c0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00161] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002c2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00162] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002c4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00163] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002c6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00164] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002c8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00165] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002ca] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00166] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002cc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00167] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002ce] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00168] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002d0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00169] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002d2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0016a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002d4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0016b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002d6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0016c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002d8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0016d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002da] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0016e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002dc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0016f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002de] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00170] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002e0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00171] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002e2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00172] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002e4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00173] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002e6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00174] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002e8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00175] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002ea] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00176] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002ec] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00177] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002ee] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00178] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002f0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00179] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002f2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0017a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002f4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0017b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002f6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0017c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002f8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0017d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002fa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0017e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002fc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0017f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h002fe] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00180] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00300] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00181] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00302] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00182] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00304] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00183] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00306] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00184] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00308] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00185] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0030a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00186] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0030c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00187] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0030e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00188] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00310] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00189] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00312] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0018a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00314] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0018b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00316] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0018c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00318] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0018d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0031a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0018e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0031c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0018f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0031e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00190] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00320] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00191] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00322] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00192] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00324] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00193] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00326] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00194] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00328] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00195] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0032a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00196] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0032c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00197] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0032e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00198] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00330] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00199] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00332] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0019a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00334] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0019b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00336] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0019c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00338] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0019d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0033a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0019e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0033c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0019f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0033e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001a0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00340] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001a1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00342] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001a2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00344] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001a3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00346] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001a4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00348] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001a5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0034a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001a6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0034c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001a7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0034e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001a8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00350] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001a9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00352] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001aa] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00354] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001ab] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00356] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001ac] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00358] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001ad] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0035a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001ae] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0035c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001af] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0035e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001b0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00360] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001b1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00362] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001b2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00364] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001b3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00366] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001b4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00368] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001b5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0036a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001b6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0036c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001b7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0036e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001b8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00370] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001b9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00372] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001ba] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00374] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001bb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00376] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001bc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00378] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001bd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0037a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001be] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0037c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001bf] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0037e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001c0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00380] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001c1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00382] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001c2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00384] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001c3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00386] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001c4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00388] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001c5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0038a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001c6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0038c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001c7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0038e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001c8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00390] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001c9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00392] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001ca] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00394] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001cb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00396] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001cc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00398] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001cd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0039a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001ce] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0039c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001cf] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0039e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001d0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003a0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001d1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003a2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001d2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003a4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001d3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003a6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001d4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003a8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001d5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003aa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001d6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003ac] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001d7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003ae] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001d8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003b0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001d9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003b2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001da] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003b4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001db] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003b6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001dc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003b8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001dd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003ba] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001de] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003bc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001df] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003be] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001e0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003c0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001e1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003c2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001e2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003c4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001e3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003c6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001e4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003c8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001e5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003ca] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001e6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003cc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001e7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003ce] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001e8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003d0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001e9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003d2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001ea] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003d4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001eb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003d6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001ec] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003d8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001ed] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003da] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001ee] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003dc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001ef] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003de] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001f0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003e0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001f1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003e2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001f2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003e4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001f3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003e6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001f4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003e8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001f5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003ea] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001f6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003ec] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001f7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003ee] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001f8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003f0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001f9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003f2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001fa] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003f4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001fb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003f6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001fc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003f8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001fd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003fa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001fe] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003fc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h001ff] =  Ic8a4ab93493bd6cdd4939054e46d2247['h003fe] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00200] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00400] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00201] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00402] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00202] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00404] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00203] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00406] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00204] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00408] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00205] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0040a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00206] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0040c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00207] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0040e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00208] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00410] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00209] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00412] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0020a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00414] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0020b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00416] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0020c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00418] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0020d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0041a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0020e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0041c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0020f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0041e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00210] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00420] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00211] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00422] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00212] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00424] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00213] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00426] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00214] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00428] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00215] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0042a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00216] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0042c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00217] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0042e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00218] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00430] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00219] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00432] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0021a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00434] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0021b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00436] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0021c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00438] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0021d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0043a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0021e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0043c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0021f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0043e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00220] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00440] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00221] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00442] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00222] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00444] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00223] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00446] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00224] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00448] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00225] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0044a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00226] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0044c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00227] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0044e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00228] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00450] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00229] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00452] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0022a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00454] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0022b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00456] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0022c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00458] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0022d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0045a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0022e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0045c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0022f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0045e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00230] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00460] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00231] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00462] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00232] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00464] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00233] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00466] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00234] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00468] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00235] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0046a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00236] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0046c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00237] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0046e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00238] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00470] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00239] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00472] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0023a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00474] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0023b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00476] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0023c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00478] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0023d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0047a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0023e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0047c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0023f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0047e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00240] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00480] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00241] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00482] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00242] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00484] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00243] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00486] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00244] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00488] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00245] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0048a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00246] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0048c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00247] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0048e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00248] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00490] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00249] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00492] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0024a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00494] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0024b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00496] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0024c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00498] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0024d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0049a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0024e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0049c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0024f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0049e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00250] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004a0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00251] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004a2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00252] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004a4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00253] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004a6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00254] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004a8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00255] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004aa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00256] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004ac] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00257] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004ae] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00258] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004b0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00259] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004b2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0025a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004b4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0025b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004b6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0025c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004b8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0025d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004ba] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0025e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004bc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0025f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004be] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00260] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004c0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00261] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004c2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00262] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004c4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00263] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004c6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00264] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004c8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00265] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004ca] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00266] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004cc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00267] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004ce] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00268] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004d0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00269] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004d2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0026a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004d4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0026b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004d6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0026c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004d8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0026d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004da] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0026e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004dc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0026f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004de] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00270] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004e0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00271] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004e2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00272] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004e4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00273] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004e6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00274] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004e8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00275] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004ea] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00276] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004ec] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00277] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004ee] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00278] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004f0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00279] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004f2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0027a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004f4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0027b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004f6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0027c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004f8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0027d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004fa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0027e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004fc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0027f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h004fe] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00280] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00500] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00281] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00502] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00282] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00504] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00283] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00506] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00284] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00508] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00285] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0050a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00286] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0050c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00287] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0050e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00288] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00510] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00289] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00512] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0028a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00514] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0028b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00516] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0028c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00518] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0028d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0051a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0028e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0051c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0028f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0051e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00290] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00520] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00291] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00522] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00292] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00524] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00293] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00526] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00294] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00528] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00295] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0052a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00296] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0052c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00297] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0052e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00298] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00530] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00299] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00532] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0029a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00534] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0029b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00536] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0029c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00538] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0029d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0053a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0029e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0053c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0029f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0053e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002a0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00540] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002a1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00542] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002a2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00544] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002a3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00546] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002a4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00548] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002a5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0054a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002a6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0054c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002a7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0054e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002a8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00550] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002a9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00552] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002aa] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00554] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002ab] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00556] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002ac] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00558] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002ad] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0055a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002ae] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0055c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002af] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0055e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002b0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00560] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002b1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00562] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002b2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00564] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002b3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00566] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002b4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00568] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002b5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0056a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002b6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0056c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002b7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0056e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002b8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00570] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002b9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00572] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002ba] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00574] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002bb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00576] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002bc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00578] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002bd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0057a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002be] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0057c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002bf] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0057e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002c0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00580] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002c1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00582] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002c2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00584] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002c3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00586] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002c4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00588] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002c5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0058a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002c6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0058c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002c7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0058e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002c8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00590] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002c9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00592] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002ca] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00594] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002cb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00596] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002cc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00598] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002cd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0059a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002ce] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0059c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002cf] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0059e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002d0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005a0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002d1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005a2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002d2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005a4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002d3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005a6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002d4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005a8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002d5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005aa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002d6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005ac] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002d7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005ae] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002d8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005b0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002d9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005b2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002da] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005b4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002db] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005b6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002dc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005b8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002dd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005ba] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002de] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005bc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002df] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005be] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002e0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005c0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002e1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005c2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002e2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005c4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002e3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005c6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002e4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005c8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002e5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005ca] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002e6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005cc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002e7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005ce] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002e8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005d0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002e9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005d2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002ea] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005d4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002eb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005d6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002ec] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005d8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002ed] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005da] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002ee] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005dc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002ef] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005de] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002f0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005e0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002f1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005e2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002f2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005e4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002f3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005e6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002f4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005e8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002f5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005ea] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002f6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005ec] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002f7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005ee] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002f8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005f0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002f9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005f2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002fa] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005f4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002fb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005f6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002fc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005f8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002fd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005fa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002fe] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005fc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h002ff] =  Ic8a4ab93493bd6cdd4939054e46d2247['h005fe] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00300] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00600] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00301] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00602] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00302] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00604] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00303] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00606] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00304] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00608] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00305] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0060a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00306] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0060c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00307] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0060e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00308] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00610] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00309] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00612] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0030a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00614] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0030b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00616] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0030c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00618] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0030d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0061a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0030e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0061c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0030f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0061e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00310] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00620] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00311] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00622] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00312] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00624] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00313] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00626] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00314] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00628] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00315] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0062a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00316] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0062c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00317] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0062e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00318] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00630] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00319] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00632] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0031a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00634] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0031b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00636] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0031c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00638] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0031d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0063a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0031e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0063c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0031f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0063e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00320] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00640] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00321] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00642] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00322] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00644] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00323] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00646] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00324] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00648] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00325] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0064a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00326] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0064c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00327] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0064e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00328] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00650] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00329] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00652] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0032a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00654] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0032b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00656] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0032c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00658] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0032d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0065a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0032e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0065c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0032f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0065e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00330] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00660] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00331] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00662] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00332] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00664] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00333] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00666] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00334] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00668] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00335] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0066a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00336] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0066c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00337] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0066e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00338] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00670] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00339] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00672] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0033a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00674] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0033b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00676] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0033c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00678] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0033d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0067a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0033e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0067c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0033f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0067e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00340] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00680] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00341] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00682] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00342] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00684] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00343] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00686] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00344] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00688] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00345] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0068a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00346] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0068c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00347] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0068e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00348] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00690] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00349] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00692] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0034a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00694] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0034b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00696] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0034c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00698] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0034d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0069a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0034e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0069c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0034f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0069e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00350] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006a0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00351] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006a2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00352] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006a4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00353] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006a6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00354] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006a8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00355] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006aa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00356] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006ac] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00357] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006ae] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00358] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006b0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00359] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006b2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0035a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006b4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0035b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006b6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0035c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006b8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0035d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006ba] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0035e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006bc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0035f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006be] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00360] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006c0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00361] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006c2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00362] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006c4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00363] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006c6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00364] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006c8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00365] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006ca] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00366] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006cc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00367] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006ce] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00368] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006d0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00369] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006d2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0036a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006d4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0036b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006d6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0036c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006d8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0036d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006da] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0036e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006dc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0036f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006de] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00370] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006e0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00371] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006e2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00372] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006e4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00373] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006e6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00374] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006e8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00375] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006ea] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00376] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006ec] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00377] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006ee] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00378] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006f0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00379] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006f2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0037a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006f4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0037b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006f6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0037c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006f8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0037d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006fa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0037e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006fc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0037f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h006fe] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00380] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00700] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00381] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00702] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00382] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00704] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00383] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00706] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00384] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00708] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00385] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0070a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00386] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0070c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00387] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0070e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00388] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00710] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00389] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00712] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0038a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00714] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0038b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00716] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0038c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00718] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0038d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0071a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0038e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0071c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0038f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0071e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00390] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00720] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00391] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00722] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00392] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00724] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00393] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00726] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00394] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00728] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00395] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0072a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00396] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0072c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00397] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0072e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00398] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00730] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00399] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00732] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0039a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00734] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0039b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00736] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0039c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00738] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0039d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0073a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0039e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0073c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0039f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0073e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003a0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00740] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003a1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00742] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003a2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00744] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003a3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00746] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003a4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00748] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003a5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0074a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003a6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0074c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003a7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0074e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003a8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00750] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003a9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00752] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003aa] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00754] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003ab] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00756] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003ac] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00758] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003ad] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0075a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003ae] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0075c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003af] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0075e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003b0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00760] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003b1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00762] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003b2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00764] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003b3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00766] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003b4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00768] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003b5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0076a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003b6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0076c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003b7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0076e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003b8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00770] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003b9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00772] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003ba] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00774] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003bb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00776] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003bc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00778] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003bd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0077a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003be] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0077c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003bf] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0077e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003c0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00780] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003c1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00782] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003c2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00784] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003c3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00786] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003c4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00788] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003c5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0078a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003c6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0078c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003c7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0078e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003c8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00790] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003c9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00792] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003ca] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00794] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003cb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00796] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003cc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00798] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003cd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0079a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003ce] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0079c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003cf] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0079e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003d0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007a0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003d1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007a2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003d2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007a4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003d3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007a6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003d4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007a8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003d5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007aa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003d6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007ac] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003d7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007ae] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003d8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007b0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003d9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007b2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003da] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007b4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003db] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007b6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003dc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007b8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003dd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007ba] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003de] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007bc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003df] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007be] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003e0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007c0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003e1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007c2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003e2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007c4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003e3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007c6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003e4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007c8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003e5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007ca] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003e6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007cc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003e7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007ce] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003e8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007d0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003e9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007d2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003ea] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007d4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003eb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007d6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003ec] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007d8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003ed] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007da] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003ee] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007dc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003ef] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007de] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003f0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007e0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003f1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007e2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003f2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007e4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003f3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007e6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003f4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007e8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003f5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007ea] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003f6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007ec] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003f7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007ee] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003f8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007f0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003f9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007f2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003fa] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007f4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003fb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007f6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003fc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007f8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003fd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007fa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003fe] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007fc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h003ff] =  Ic8a4ab93493bd6cdd4939054e46d2247['h007fe] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00400] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00800] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00401] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00802] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00402] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00804] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00403] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00806] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00404] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00808] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00405] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0080a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00406] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0080c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00407] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0080e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00408] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00810] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00409] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00812] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0040a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00814] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0040b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00816] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0040c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00818] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0040d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0081a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0040e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0081c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0040f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0081e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00410] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00820] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00411] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00822] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00412] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00824] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00413] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00826] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00414] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00828] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00415] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0082a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00416] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0082c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00417] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0082e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00418] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00830] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00419] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00832] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0041a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00834] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0041b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00836] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0041c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00838] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0041d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0083a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0041e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0083c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0041f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0083e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00420] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00840] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00421] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00842] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00422] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00844] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00423] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00846] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00424] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00848] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00425] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0084a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00426] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0084c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00427] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0084e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00428] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00850] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00429] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00852] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0042a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00854] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0042b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00856] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0042c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00858] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0042d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0085a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0042e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0085c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0042f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0085e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00430] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00860] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00431] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00862] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00432] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00864] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00433] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00866] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00434] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00868] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00435] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0086a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00436] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0086c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00437] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0086e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00438] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00870] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00439] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00872] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0043a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00874] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0043b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00876] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0043c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00878] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0043d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0087a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0043e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0087c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0043f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0087e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00440] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00880] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00441] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00882] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00442] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00884] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00443] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00886] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00444] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00888] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00445] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0088a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00446] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0088c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00447] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0088e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00448] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00890] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00449] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00892] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0044a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00894] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0044b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00896] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0044c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00898] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0044d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0089a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0044e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0089c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0044f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0089e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00450] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008a0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00451] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008a2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00452] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008a4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00453] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008a6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00454] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008a8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00455] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008aa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00456] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008ac] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00457] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008ae] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00458] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008b0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00459] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008b2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0045a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008b4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0045b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008b6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0045c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008b8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0045d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008ba] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0045e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008bc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0045f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008be] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00460] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008c0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00461] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008c2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00462] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008c4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00463] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008c6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00464] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008c8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00465] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008ca] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00466] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008cc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00467] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008ce] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00468] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008d0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00469] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008d2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0046a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008d4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0046b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008d6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0046c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008d8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0046d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008da] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0046e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008dc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0046f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008de] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00470] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008e0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00471] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008e2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00472] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008e4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00473] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008e6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00474] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008e8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00475] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008ea] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00476] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008ec] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00477] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008ee] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00478] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008f0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00479] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008f2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0047a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008f4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0047b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008f6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0047c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008f8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0047d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008fa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0047e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008fc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0047f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h008fe] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00480] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00900] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00481] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00902] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00482] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00904] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00483] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00906] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00484] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00908] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00485] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0090a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00486] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0090c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00487] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0090e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00488] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00910] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00489] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00912] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0048a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00914] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0048b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00916] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0048c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00918] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0048d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0091a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0048e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0091c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0048f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0091e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00490] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00920] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00491] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00922] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00492] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00924] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00493] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00926] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00494] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00928] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00495] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0092a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00496] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0092c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00497] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0092e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00498] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00930] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00499] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00932] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0049a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00934] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0049b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00936] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0049c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00938] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0049d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0093a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0049e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0093c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0049f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0093e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004a0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00940] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004a1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00942] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004a2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00944] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004a3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00946] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004a4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00948] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004a5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0094a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004a6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0094c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004a7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0094e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004a8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00950] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004a9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00952] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004aa] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00954] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004ab] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00956] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004ac] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00958] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004ad] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0095a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004ae] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0095c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004af] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0095e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004b0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00960] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004b1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00962] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004b2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00964] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004b3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00966] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004b4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00968] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004b5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0096a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004b6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0096c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004b7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0096e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004b8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00970] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004b9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00972] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004ba] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00974] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004bb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00976] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004bc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00978] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004bd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0097a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004be] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0097c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004bf] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0097e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004c0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00980] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004c1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00982] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004c2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00984] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004c3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00986] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004c4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00988] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004c5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0098a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004c6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0098c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004c7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0098e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004c8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00990] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004c9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00992] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004ca] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00994] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004cb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00996] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004cc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00998] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004cd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0099a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004ce] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0099c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004cf] =  Ic8a4ab93493bd6cdd4939054e46d2247['h0099e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004d0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009a0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004d1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009a2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004d2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009a4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004d3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009a6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004d4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009a8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004d5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009aa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004d6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009ac] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004d7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009ae] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004d8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009b0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004d9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009b2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004da] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009b4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004db] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009b6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004dc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009b8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004dd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009ba] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004de] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009bc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004df] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009be] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004e0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009c0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004e1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009c2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004e2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009c4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004e3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009c6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004e4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009c8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004e5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009ca] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004e6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009cc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004e7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009ce] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004e8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009d0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004e9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009d2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004ea] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009d4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004eb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009d6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004ec] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009d8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004ed] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009da] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004ee] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009dc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004ef] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009de] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004f0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009e0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004f1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009e2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004f2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009e4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004f3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009e6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004f4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009e8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004f5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009ea] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004f6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009ec] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004f7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009ee] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004f8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009f0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004f9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009f2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004fa] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009f4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004fb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009f6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004fc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009f8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004fd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009fa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004fe] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009fc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h004ff] =  Ic8a4ab93493bd6cdd4939054e46d2247['h009fe] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00500] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a00] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00501] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a02] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00502] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a04] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00503] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a06] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00504] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a08] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00505] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a0a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00506] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a0c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00507] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a0e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00508] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a10] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00509] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a12] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0050a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a14] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0050b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a16] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0050c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a18] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0050d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a1a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0050e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a1c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0050f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a1e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00510] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a20] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00511] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a22] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00512] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a24] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00513] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a26] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00514] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a28] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00515] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a2a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00516] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a2c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00517] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a2e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00518] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a30] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00519] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a32] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0051a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a34] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0051b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a36] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0051c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a38] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0051d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a3a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0051e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a3c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0051f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a3e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00520] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a40] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00521] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a42] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00522] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a44] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00523] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a46] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00524] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a48] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00525] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a4a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00526] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a4c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00527] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a4e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00528] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a50] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00529] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a52] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0052a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a54] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0052b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a56] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0052c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a58] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0052d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a5a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0052e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a5c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0052f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a5e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00530] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a60] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00531] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a62] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00532] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a64] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00533] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a66] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00534] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a68] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00535] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a6a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00536] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a6c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00537] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a6e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00538] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a70] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00539] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a72] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0053a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a74] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0053b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a76] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0053c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a78] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0053d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a7a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0053e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a7c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0053f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a7e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00540] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a80] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00541] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a82] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00542] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a84] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00543] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a86] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00544] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a88] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00545] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a8a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00546] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a8c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00547] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a8e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00548] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a90] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00549] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a92] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0054a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a94] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0054b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a96] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0054c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a98] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0054d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a9a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0054e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a9c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0054f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00a9e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00550] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00aa0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00551] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00aa2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00552] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00aa4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00553] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00aa6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00554] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00aa8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00555] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00aaa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00556] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00aac] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00557] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00aae] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00558] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ab0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00559] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ab2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0055a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ab4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0055b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ab6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0055c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ab8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0055d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00aba] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0055e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00abc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0055f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00abe] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00560] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ac0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00561] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ac2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00562] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ac4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00563] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ac6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00564] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ac8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00565] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00aca] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00566] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00acc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00567] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ace] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00568] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ad0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00569] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ad2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0056a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ad4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0056b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ad6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0056c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ad8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0056d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ada] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0056e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00adc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0056f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ade] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00570] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ae0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00571] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ae2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00572] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ae4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00573] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ae6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00574] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ae8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00575] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00aea] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00576] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00aec] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00577] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00aee] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00578] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00af0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00579] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00af2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0057a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00af4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0057b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00af6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0057c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00af8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0057d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00afa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0057e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00afc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0057f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00afe] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00580] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b00] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00581] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b02] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00582] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b04] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00583] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b06] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00584] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b08] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00585] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b0a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00586] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b0c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00587] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b0e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00588] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b10] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00589] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b12] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0058a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b14] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0058b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b16] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0058c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b18] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0058d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b1a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0058e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b1c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0058f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b1e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00590] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b20] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00591] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b22] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00592] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b24] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00593] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b26] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00594] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b28] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00595] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b2a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00596] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b2c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00597] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b2e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00598] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b30] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00599] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b32] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0059a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b34] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0059b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b36] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0059c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b38] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0059d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b3a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0059e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b3c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0059f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b3e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005a0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b40] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005a1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b42] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005a2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b44] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005a3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b46] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005a4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b48] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005a5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b4a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005a6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b4c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005a7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b4e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005a8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b50] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005a9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b52] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005aa] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b54] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005ab] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b56] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005ac] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b58] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005ad] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b5a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005ae] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b5c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005af] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b5e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005b0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b60] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005b1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b62] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005b2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b64] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005b3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b66] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005b4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b68] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005b5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b6a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005b6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b6c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005b7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b6e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005b8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b70] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005b9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b72] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005ba] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b74] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005bb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b76] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005bc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b78] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005bd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b7a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005be] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b7c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005bf] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b7e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005c0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b80] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005c1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b82] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005c2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b84] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005c3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b86] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005c4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b88] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005c5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b8a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005c6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b8c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005c7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b8e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005c8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b90] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005c9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b92] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005ca] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b94] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005cb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b96] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005cc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b98] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005cd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b9a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005ce] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b9c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005cf] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00b9e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005d0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ba0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005d1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ba2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005d2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ba4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005d3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ba6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005d4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ba8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005d5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00baa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005d6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bac] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005d7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bae] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005d8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bb0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005d9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bb2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005da] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bb4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005db] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bb6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005dc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bb8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005dd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bba] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005de] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bbc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005df] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bbe] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005e0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bc0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005e1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bc2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005e2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bc4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005e3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bc6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005e4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bc8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005e5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bca] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005e6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bcc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005e7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bce] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005e8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bd0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005e9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bd2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005ea] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bd4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005eb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bd6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005ec] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bd8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005ed] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bda] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005ee] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bdc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005ef] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bde] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005f0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00be0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005f1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00be2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005f2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00be4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005f3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00be6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005f4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00be8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005f5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bea] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005f6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bec] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005f7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bee] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005f8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bf0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005f9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bf2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005fa] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bf4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005fb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bf6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005fc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bf8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005fd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bfa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005fe] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bfc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h005ff] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00bfe] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00600] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c00] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00601] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c02] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00602] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c04] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00603] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c06] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00604] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c08] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00605] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c0a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00606] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c0c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00607] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c0e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00608] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c10] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00609] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c12] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0060a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c14] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0060b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c16] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0060c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c18] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0060d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c1a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0060e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c1c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0060f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c1e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00610] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c20] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00611] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c22] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00612] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c24] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00613] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c26] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00614] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c28] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00615] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c2a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00616] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c2c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00617] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c2e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00618] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c30] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00619] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c32] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0061a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c34] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0061b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c36] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0061c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c38] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0061d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c3a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0061e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c3c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0061f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c3e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00620] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c40] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00621] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c42] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00622] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c44] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00623] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c46] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00624] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c48] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00625] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c4a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00626] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c4c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00627] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c4e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00628] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c50] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00629] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c52] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0062a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c54] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0062b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c56] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0062c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c58] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0062d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c5a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0062e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c5c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0062f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c5e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00630] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c60] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00631] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c62] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00632] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c64] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00633] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c66] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00634] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c68] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00635] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c6a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00636] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c6c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00637] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c6e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00638] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c70] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00639] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c72] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0063a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c74] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0063b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c76] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0063c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c78] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0063d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c7a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0063e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c7c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0063f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c7e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00640] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c80] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00641] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c82] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00642] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c84] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00643] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c86] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00644] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c88] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00645] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c8a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00646] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c8c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00647] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c8e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00648] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c90] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00649] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c92] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0064a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c94] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0064b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c96] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0064c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c98] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0064d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c9a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0064e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c9c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0064f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00c9e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00650] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ca0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00651] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ca2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00652] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ca4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00653] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ca6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00654] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ca8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00655] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00caa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00656] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cac] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00657] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cae] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00658] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cb0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00659] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cb2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0065a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cb4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0065b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cb6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0065c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cb8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0065d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cba] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0065e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cbc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0065f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cbe] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00660] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cc0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00661] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cc2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00662] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cc4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00663] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cc6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00664] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cc8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00665] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cca] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00666] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ccc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00667] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cce] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00668] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cd0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00669] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cd2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0066a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cd4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0066b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cd6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0066c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cd8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0066d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cda] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0066e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cdc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0066f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cde] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00670] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ce0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00671] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ce2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00672] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ce4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00673] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ce6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00674] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ce8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00675] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cea] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00676] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cec] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00677] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cee] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00678] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cf0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00679] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cf2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0067a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cf4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0067b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cf6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0067c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cf8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0067d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cfa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0067e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cfc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0067f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00cfe] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00680] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d00] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00681] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d02] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00682] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d04] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00683] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d06] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00684] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d08] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00685] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d0a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00686] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d0c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00687] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d0e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00688] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d10] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00689] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d12] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0068a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d14] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0068b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d16] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0068c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d18] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0068d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d1a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0068e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d1c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0068f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d1e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00690] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d20] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00691] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d22] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00692] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d24] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00693] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d26] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00694] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d28] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00695] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d2a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00696] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d2c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00697] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d2e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00698] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d30] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00699] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d32] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0069a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d34] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0069b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d36] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0069c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d38] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0069d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d3a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0069e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d3c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0069f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d3e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006a0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d40] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006a1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d42] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006a2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d44] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006a3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d46] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006a4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d48] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006a5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d4a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006a6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d4c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006a7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d4e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006a8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d50] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006a9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d52] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006aa] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d54] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006ab] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d56] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006ac] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d58] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006ad] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d5a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006ae] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d5c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006af] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d5e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006b0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d60] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006b1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d62] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006b2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d64] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006b3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d66] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006b4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d68] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006b5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d6a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006b6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d6c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006b7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d6e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006b8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d70] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006b9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d72] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006ba] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d74] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006bb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d76] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006bc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d78] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006bd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d7a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006be] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d7c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006bf] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d7e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006c0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d80] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006c1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d82] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006c2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d84] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006c3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d86] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006c4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d88] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006c5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d8a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006c6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d8c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006c7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d8e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006c8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d90] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006c9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d92] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006ca] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d94] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006cb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d96] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006cc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d98] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006cd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d9a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006ce] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d9c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006cf] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00d9e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006d0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00da0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006d1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00da2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006d2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00da4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006d3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00da6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006d4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00da8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006d5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00daa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006d6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00dac] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006d7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00dae] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006d8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00db0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006d9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00db2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006da] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00db4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006db] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00db6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006dc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00db8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006dd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00dba] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006de] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00dbc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006df] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00dbe] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006e0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00dc0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006e1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00dc2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006e2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00dc4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006e3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00dc6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006e4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00dc8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006e5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00dca] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006e6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00dcc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006e7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00dce] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006e8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00dd0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006e9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00dd2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006ea] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00dd4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006eb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00dd6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006ec] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00dd8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006ed] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00dda] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006ee] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ddc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006ef] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00dde] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006f0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00de0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006f1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00de2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006f2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00de4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006f3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00de6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006f4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00de8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006f5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00dea] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006f6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00dec] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006f7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00dee] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006f8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00df0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006f9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00df2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006fa] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00df4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006fb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00df6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006fc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00df8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006fd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00dfa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006fe] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00dfc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h006ff] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00dfe] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00700] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e00] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00701] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e02] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00702] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e04] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00703] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e06] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00704] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e08] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00705] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e0a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00706] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e0c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00707] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e0e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00708] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e10] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00709] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e12] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0070a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e14] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0070b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e16] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0070c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e18] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0070d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e1a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0070e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e1c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0070f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e1e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00710] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e20] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00711] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e22] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00712] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e24] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00713] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e26] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00714] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e28] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00715] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e2a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00716] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e2c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00717] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e2e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00718] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e30] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00719] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e32] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0071a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e34] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0071b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e36] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0071c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e38] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0071d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e3a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0071e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e3c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0071f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e3e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00720] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e40] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00721] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e42] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00722] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e44] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00723] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e46] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00724] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e48] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00725] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e4a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00726] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e4c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00727] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e4e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00728] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e50] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00729] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e52] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0072a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e54] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0072b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e56] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0072c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e58] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0072d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e5a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0072e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e5c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0072f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e5e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00730] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e60] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00731] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e62] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00732] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e64] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00733] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e66] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00734] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e68] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00735] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e6a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00736] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e6c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00737] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e6e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00738] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e70] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00739] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e72] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0073a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e74] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0073b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e76] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0073c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e78] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0073d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e7a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0073e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e7c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0073f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e7e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00740] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e80] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00741] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e82] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00742] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e84] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00743] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e86] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00744] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e88] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00745] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e8a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00746] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e8c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00747] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e8e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00748] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e90] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00749] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e92] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0074a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e94] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0074b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e96] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0074c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e98] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0074d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e9a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0074e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e9c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0074f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00e9e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00750] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ea0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00751] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ea2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00752] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ea4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00753] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ea6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00754] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ea8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00755] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00eaa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00756] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00eac] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00757] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00eae] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00758] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00eb0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00759] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00eb2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0075a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00eb4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0075b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00eb6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0075c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00eb8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0075d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00eba] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0075e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ebc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0075f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ebe] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00760] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ec0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00761] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ec2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00762] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ec4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00763] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ec6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00764] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ec8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00765] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00eca] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00766] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ecc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00767] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ece] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00768] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ed0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00769] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ed2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0076a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ed4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0076b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ed6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0076c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ed8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0076d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00eda] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0076e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00edc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0076f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ede] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00770] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ee0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00771] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ee2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00772] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ee4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00773] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ee6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00774] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ee8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00775] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00eea] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00776] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00eec] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00777] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00eee] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00778] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ef0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00779] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ef2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0077a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ef4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0077b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ef6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0077c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ef8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0077d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00efa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0077e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00efc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0077f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00efe] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00780] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f00] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00781] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f02] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00782] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f04] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00783] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f06] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00784] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f08] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00785] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f0a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00786] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f0c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00787] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f0e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00788] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f10] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00789] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f12] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0078a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f14] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0078b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f16] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0078c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f18] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0078d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f1a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0078e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f1c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0078f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f1e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00790] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f20] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00791] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f22] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00792] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f24] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00793] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f26] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00794] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f28] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00795] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f2a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00796] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f2c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00797] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f2e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00798] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f30] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h00799] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f32] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0079a] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f34] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0079b] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f36] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0079c] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f38] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0079d] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f3a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0079e] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f3c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h0079f] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f3e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007a0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f40] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007a1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f42] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007a2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f44] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007a3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f46] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007a4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f48] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007a5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f4a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007a6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f4c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007a7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f4e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007a8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f50] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007a9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f52] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007aa] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f54] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007ab] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f56] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007ac] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f58] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007ad] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f5a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007ae] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f5c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007af] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f5e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007b0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f60] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007b1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f62] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007b2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f64] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007b3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f66] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007b4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f68] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007b5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f6a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007b6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f6c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007b7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f6e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007b8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f70] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007b9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f72] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007ba] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f74] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007bb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f76] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007bc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f78] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007bd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f7a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007be] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f7c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007bf] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f7e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007c0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f80] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007c1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f82] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007c2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f84] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007c3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f86] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007c4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f88] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007c5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f8a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007c6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f8c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007c7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f8e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007c8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f90] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007c9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f92] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007ca] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f94] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007cb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f96] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007cc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f98] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007cd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f9a] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007ce] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f9c] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007cf] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00f9e] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007d0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fa0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007d1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fa2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007d2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fa4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007d3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fa6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007d4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fa8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007d5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00faa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007d6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fac] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007d7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fae] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007d8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fb0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007d9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fb2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007da] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fb4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007db] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fb6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007dc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fb8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007dd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fba] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007de] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fbc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007df] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fbe] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007e0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fc0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007e1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fc2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007e2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fc4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007e3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fc6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007e4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fc8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007e5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fca] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007e6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fcc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007e7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fce] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007e8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fd0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007e9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fd2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007ea] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fd4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007eb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fd6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007ec] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fd8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007ed] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fda] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007ee] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fdc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007ef] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fde] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007f0] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fe0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007f1] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fe2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007f2] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fe4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007f3] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fe6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007f4] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fe8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007f5] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fea] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007f6] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fec] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007f7] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00fee] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007f8] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ff0] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007f9] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ff2] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007fa] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ff4] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007fb] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ff6] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007fc] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ff8] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007fd] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ffa] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007fe] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ffc] ;
//end
//always_comb begin // 
               Ia940d1a12f2aecb1cf57d9d7b9e7b4aa['h007ff] =  Ic8a4ab93493bd6cdd4939054e46d2247['h00ffe] ;
//end
