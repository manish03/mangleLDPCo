 reg  ['hffff:0] [$clog2('h7000+1)-1:0] Ib26a88d1741ee737acfeaa5e34cb90db ;
