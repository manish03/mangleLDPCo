              Iad95cb311111b88124c0d2a123589b68 = 
          (!fgallag_sel[4]) ? 
                       I03b14329c0d52c7997914a8d9ab65fed: 
                       I63a4e0a46ca3426e2cb066ad3bfc245d;
              I8efbaa789c07fd87b2bd52379ef30fd6 = 
          (!fgallag_sel[4]) ? 
                       Ie21703557f53d7bf9cf79a7f6c1d5958: 
                       I3a7b809a0160dee33125934243952cdc;
              I75d6885c5406c2c71dc966efa9c6826d = 
          (!fgallag_sel[4]) ? 
                       I1cb33fdd3dac4dda0b25adbab30d2913: 
                       Ia6905a32e1257061364dd1249fa76bf2;
              I3f698aa4ba3738ea0af307eff19d7322 = 
          (!fgallag_sel[4]) ? 
                       Id2b87d69ba4c78cf41a7be349397ad5e: 
                       I7d9d74dbceb047ad0c76322038fbf229;
              I3dcfc9ea0f47bae945b7b823693115ad = 
          (!fgallag_sel[4]) ? 
                       I856e4e862c70da83553a3dba9edea1ab: 
                       Iaf42178313f7b4aa6ce6090ecbf2b3b6;
              Id1a3fd12101241027e2f457a826ed09d = 
          (!fgallag_sel[4]) ? 
                       Id7a56c8135dad1fd457d336f7a632436: 
                       I2ffc40e4b0cc841bd3c8d7519fc4512a;
              I7bfcc4e396adf33cfc50d06be12d9007 = 
          (!fgallag_sel[4]) ? 
                       I20c0389215371104437ef298cb12b3c4: 
                       Ie4e1b20f36ecda5d4d917a241ef2a1fd;
              I5ce36b9e0a8e3e118e1f1b9eae183b7b = 
          (!fgallag_sel[4]) ? 
                       Icf120a29648cb8af4bae9e4343f13a40: 
                       I1e317164e9010fb6755c65adda38ea2a;
              I98f08554298bf8e87fc54a4f8c668314 = 
          (!fgallag_sel[4]) ? 
                       I0f5a57095bb2bbf99b71f04a19e2c38f: 
                       Ib52869a26824ee42fff6262100e1ebe5;
               Ic05153bb88b7db4e173fd73841f88bf2 =  I61ff69ca863e90ffc9118f12c5aa3b14 ;
               I75df32ec8d8f7096f5f7ef1d17cfb8e7 =  I08f41ede762b72d92816c6dff8e074f9 ;
              Ia3c542d3f12470683609d561d9cd0e35 = 
          (!fgallag_sel[4]) ? 
                       I912919c7cfae1b4827ca945a92a5310c: 
                       Icd7b7d17911094c9fa48fc5906968dcd;
