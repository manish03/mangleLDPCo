//#;; Id7d2c4b2da7a6478426f10a28d9f9eba59a188d1bf2835798742825d32a11125 I8be3365cabaa6a0f90d2e64f03fa78268c135fe0b0758b576b447e9b2068d75d I18a0c098c7fb0098093fc0fd619c8032ae193215c5f695d7f5eaafa28aa64d70 I679eaac16659c013675081e715f7ef761bdd183f1d7f55d079eb46ad6e322ac5 I9ef2faffd23e7fdda264eeeb3114357fcb304142506cbb023c2894ac10f71654
/*Ic3f8d45b35548e4a4ee0b7181f1834df8a2e1aa0eea9b8c77323fcbf46bb42c8*/
////////////////////////////////////////////////////////////////////////////////
//# Copyright (c) 2018 Secantec
//# No Permission to modify and distribute this program
//# even if this copyright message remains unaltered.
//#
//# Author: Secantec 27 April, 2018
//# $Id: $//#
//# Revision History
//#       MM      17  April, 2018    Initial release
//#
////////////////////////////////////////////////////////////////////////////////

// /I51a1f05af85e342e3c849b47d387086476282d5f50dc240c19216d6edfb1eb5a/I58466ebdd352f801198118e294e38715f864985fd87977f348bfcd7db62e7c76 -I54e67ab9c29a6cfd19408098a96b2a40ede7e06aadcf77336da0dd2b57f25ba7 *I4395dc236d13a1c9b88a791fd2e1275bbb97b927d52e9b8c38248a0d57259aea* *Ic7c59e97212940ba254bbb99e5f908fec3434155e0fbb2f0a3f2ab5a6b4ba2a1* ; If0c929a9e723bc62724e30c7e396e576019dfcb8cfd0a3f264ee5d72e64e49d1 I04ad2bfad8cbdb3afbf9a26ea1454ac0a07c0eebc856992b38114cdcb5098c47.I3485639faf1591f3c16f295198e9389db5b33c949587ec48663597d4e00299d5 -If0c929a9e723bc62724e30c7e396e576019dfcb8cfd0a3f264ee5d72e64e49d1 I8803a3b234be60475d3d6498d388264bbc5edd49f43c780eee4753cddabfe052.1.sv > I8803a3b234be60475d3d6498d388264bbc5edd49f43c780eee4753cddabfe052.1.I04ad2bfad8cbdb3afbf9a26ea1454ac0a07c0eebc856992b38114cdcb5098c47.sv ; Ia8d1cfa1fc63160715eed9e8f5f39538f4520ff839d850162536352ec0a5509c -Ic572272153455b732903e10d0db7356fb56fb5d0a6a9064766547a1304406c33 -I8c2574892063f995fdf756bce07f46c1a5193e54cd52837ed91e32008ccf41ac -I4e1de0094e501762cba645b8d4663534d3eee7dc7d8bc675574f6b130d9f5302 I8803a3b234be60475d3d6498d388264bbc5edd49f43c780eee4753cddabfe052.1.I04ad2bfad8cbdb3afbf9a26ea1454ac0a07c0eebc856992b38114cdcb5098c47.sv -Iacac86c0e609ca906f632b0e2dacccb2b77d22b0621f20ebece1a4835b93f6f0 I8803a3b234be60475d3d6498d388264bbc5edd49f43c780eee4753cddabfe052.1.I04ad2bfad8cbdb3afbf9a26ea1454ac0a07c0eebc856992b38114cdcb5098c47.sv.I836ff184e7b41b1e13cb5fd89fa1de98dbbab99e9d2918913ff43b86a5c7c213

 /*Ic3f8d45b35548e4a4ee0b7181f1834df8a2e1aa0eea9b8c77323fcbf46bb42c8*/

/* I1e4d9aa7cb1ef438f80454b61c625f0c6aed19675cb2c2f865cbd2e2c3ef2ff7 Ib8a92ab2b5e2e68fc63a575fff1d62c25ec6d30209e164d82ec85f5576d9d940 I63985ce3eb57dbe35dec3a2e0dc38ffe14d2e2396edf773bd4f0298ce3ec7eff */

module  sntc_ldpc_syndrome_tb #(
// I168413ccee11e827c207105eecf061ecb7d6991383544364fda85556cdf96a57/I373a739f28b569ba97fa09dd5a21185f9bed4792859f1d9cc7fe4af7f6b9c7b7.sv
parameter MM   = 'h 000a8 ,
// parameter MM =  'h  000a8  , 
parameter NN   = 'h 000d0 ,
// parameter NN =  'h  000d0  , 
parameter cmax = 'h 00017 ,
// parameter cmax =  'h  00017  , 
parameter rmax = 'h 0000a ,
// parameter rmax =  'h  0000a  , 
// 208
// 168
parameter SUM_NN         = $clog2(NN+1), // 8 : I47c35ffcd3135a74f03fef2155c1874927bc03c22812da0a352f40ca1d7339ea
parameter SUM_MM         = $clog2(MM+1), // 8 : Ifa20411ae2befe271235475378a99513a77cfe0a9614b7cba4d2d92a1f1168c3
parameter LEN            = MM,
parameter SUM_NN_WDTH    = $clog2(SUM_NN+2),
parameter SUM_MM_WDTH    = $clog2(SUM_MM+2),
`include "sntc_LDPC_dec_param.sv"
//parameter SUM_LEN        = SUM_MM
parameter MAX_SUM_WDTH_LONG = MAX_SUM_WDTH +1,
parameter SUM_LEN        = 32

) (

input wire clk_tb,
input wire rstn_tb
);

`ifdef ENCRYPT
`endif

int Idb5f1a085a445a011e36f2e5014265ae744db959b05c5097464d6982589f26f4[int],I736b57465bc098745b079bbf59b7645dc4548bc5e23e4805c92fa6a35eb0e3a9[int], I7a475a8b0a074fa8bd3bf54dc2a172de8c70f8ad78980010b9d8e9bc5a5b978f[int];
int I86fc979a71bc09eae1f0b85d2e5f631d3e65377de57c1febb965a4085cc413eb;
int Ib95684006fa50410fdb7b71438302187c40016e386f98ca87ff6b336489bfbd5;
real Ic549779d79e5c8e9c9a6b6da5f1c5e21075eb9319852f858acb227ee855e4ef5[int];
int Ibbeebd879e1dff6918546dc0c179fdde505f2a21591c9a9c96e36b054ec5af83[int],A[int];
string Ibeac5ed31d4582212c21a5dd06959110a37c49046ed23020de290e17d4f45815[int];



// -1 : I439cd19385ab0d52df1a0893519b39c376ecee7da819b413a351d0b857b49c68
// I168413ccee11e827c207105eecf061ecb7d6991383544364fda85556cdf96a57.I53228d397d8cfe91552c5f863bd55a4d75d54e3c665004d472d6236c0c6cf139 : Ia1ea30d9838563b7809d572210298bd5939acb28235343b05c8d231255972db6 I82a3537ff0dbce7eec35d69edc3a189ee6f17d82f353a553f9aa96cb0be3ce89


// I8c64802bb57ab85b89646541ba23fdacf78b8a4697489b96c16bdb7ff1ad3d4d : Ifbcebae39bd76915a91c43d7e4f6f230b5b27bdc6ad5e6925d5eb045636df7da 2 0 4.I53228d397d8cfe91552c5f863bd55a4d75d54e3c665004d472d6236c0c6cf139
// Ibeac5ed31d4582212c21a5dd06959110a37c49046ed23020de290e17d4f45815: 2

// Ie8ca83241b10dfad19c6d317a1706e396501e7514284da760ab031d020e48459: $NR_Z





reg  [NN-1:0]                 tmp_bit;
reg  [NN-1:0] [1:0]           I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be;
wire [MM-1:0]                 syndrome;
reg  [MM-1:0]                 exp_syn;
wire [SUM_LEN-1:0]            HamDist_sum_mm;
reg  [SUM_LEN-1:0]            HamDist_loop;
reg  [SUM_LEN-1:0]            HamDist_cntr;
reg  [SUM_LEN-1:0]            HamDist_loop_max;
reg  [SUM_LEN-1:0]            HamDist_loop_percentage;
wire [1:0]                    I16bdee165138010bda1229669cf4bb78831253202a69fa31552c0ac42725776a;
wire                          I07db8da4c1a2e19e0fb67ff37bf4b2f8d5d6db2c69639497fcab892e05942ec6;
reg                           Id5607445fd3e16ebe83d7d3a46b05dfe1dc8e5eed33f51f9f795fefdac3e44cf;
wire                          Id9ac53997afa49d1b311d681cbd804894604a5574f6121604013d48a0f15afea;
reg                           clk;
reg                           rstn;
int                           Ic6c882b049984e99a95e83ce05934d4d06d0825ce52525e4e6532757001dcaf7;
reg                           clr;
reg                           Icced28c6dc3f99c2396a5eaad732bf6b28142335892b1cd0e6af6cdb53f5ccfa;
wire                          valid;
wire [31:0]                   percent_probability_int;

reg  [SUM_LEN-1:0]            HamDist_iir1;
reg  [SUM_LEN-1:0]            HamDist_iir2;
reg  [SUM_LEN-1:0]            HamDist_iir3;
reg                           I1725d63fa57c5344aa111b908a4770db8738a8217a8d458c8af741a8df7cc480 =0;

always_comb begin
          HamDist_iir1 = 85;
          HamDist_iir2 = 15;
          HamDist_iir3 = 5;

end

wire valid_cword;
wire valid_cword_dec;
wire [NN-1:0] I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6;
reg [NN-MM-1:0] y_nr_in;
reg [NN-1:0] I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd;

sntc_ldpc_syndrome_wrapper i_sntc_ldpc_syndrome_wrapper
(


                                  .y_nr_in                (tmp_bit),
                                  .I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9                 (syndrome),
/* I1e4d9aa7cb1ef438f80454b61c625f0c6aed19675cb2c2f865cbd2e2c3ef2ff7 Ib8a92ab2b5e2e68fc63a575fff1d62c25ec6d30209e164d82ec85f5576d9d940 I5fedfe54fddcdc5145ac6dd38b4c3dead65f127535af2e07a7b9790515afdb04 */
                                  .clr                    (clr),
/* I1e4d9aa7cb1ef438f80454b61c625f0c6aed19675cb2c2f865cbd2e2c3ef2ff7 I2f08a120cf6d1091827fd5d929bad0cbcaa5eff7ae0801098357ed0149cbc06e I5fedfe54fddcdc5145ac6dd38b4c3dead65f127535af2e07a7b9790515afdb04 */
                                  .valid_cword            (valid_cword),
                                  .rstn                   (rstn),
                                  .clk                    (clk)
);





`ifdef SIMULATION
 int I2ba1a21f00560d3c11f9b8906c307417a740a8dd92ccf1fe7c4c3af48da348e1 =1;
initial
begin
  clk = 0;
  Ic6c882b049984e99a95e83ce05934d4d06d0825ce52525e4e6532757001dcaf7 = 1;
  forever
  begin
    clk = ~clk;
    if (clk) Ic6c882b049984e99a95e83ce05934d4d06d0825ce52525e4e6532757001dcaf7 = Ic6c882b049984e99a95e83ce05934d4d06d0825ce52525e4e6532757001dcaf7 + 1;
    //if (clk) if ((Ic6c882b049984e99a95e83ce05934d4d06d0825ce52525e4e6532757001dcaf7 % 1000) === 0) $display("Id69a26f56dfc4cead7151d018c424aea7b4152f95aad72fe789e4ea3d643fdd7:Ic6c882b049984e99a95e83ce05934d4d06d0825ce52525e4e6532757001dcaf7:%05d %t", Ic6c882b049984e99a95e83ce05934d4d06d0825ce52525e4e6532757001dcaf7, $time);
    if (clk) $display("Id69a26f56dfc4cead7151d018c424aea7b4152f95aad72fe789e4ea3d643fdd7:Ic6c882b049984e99a95e83ce05934d4d06d0825ce52525e4e6532757001dcaf7:%05d %t", Ic6c882b049984e99a95e83ce05934d4d06d0825ce52525e4e6532757001dcaf7, $time);
    #5;
  end
end
initial
begin
  rstn = 0;
  clr = 0;
  repeat (10) @ (posedge clk);
  rstn = 1;
end


always_comb HamDist_loop_max        =  10;
always_comb HamDist_loop_percentage =  110;

initial
begin
Idb5f1a085a445a011e36f2e5014265ae744db959b05c5097464d6982589f26f4[00]=8448;I7a475a8b0a074fa8bd3bf54dc2a172de8c70f8ad78980010b9d8e9bc5a5b978f[ 0]= 9396;A[ 0]=8832;Ibeac5ed31d4582212c21a5dd06959110a37c49046ed23020de290e17d4f45815[ 0]="I65fbe7a0709a36e2f5f6295e0e45fb58ad21e0a3c0f1f5acd39a7a9f2d529f2c";
Idb5f1a085a445a011e36f2e5014265ae744db959b05c5097464d6982589f26f4[01]=8448;I7a475a8b0a074fa8bd3bf54dc2a172de8c70f8ad78980010b9d8e9bc5a5b978f[ 1]=10566;A[ 1]=8832;Ibeac5ed31d4582212c21a5dd06959110a37c49046ed23020de290e17d4f45815[ 1]="I65fbe7a0709a36e2f5f6295e0e45fb58ad21e0a3c0f1f5acd39a7a9f2d529f2c";
Idb5f1a085a445a011e36f2e5014265ae744db959b05c5097464d6982589f26f4[02]=8448;I7a475a8b0a074fa8bd3bf54dc2a172de8c70f8ad78980010b9d8e9bc5a5b978f[ 2]= 9392;A[ 2]=8832;Ibeac5ed31d4582212c21a5dd06959110a37c49046ed23020de290e17d4f45815[ 2]="I65fbe7a0709a36e2f5f6295e0e45fb58ad21e0a3c0f1f5acd39a7a9f2d529f2c";
Idb5f1a085a445a011e36f2e5014265ae744db959b05c5097464d6982589f26f4[03]=8448;I7a475a8b0a074fa8bd3bf54dc2a172de8c70f8ad78980010b9d8e9bc5a5b978f[ 3]=12368;A[ 3]=8832;Ibeac5ed31d4582212c21a5dd06959110a37c49046ed23020de290e17d4f45815[ 3]="I65fbe7a0709a36e2f5f6295e0e45fb58ad21e0a3c0f1f5acd39a7a9f2d529f2c";
Idb5f1a085a445a011e36f2e5014265ae744db959b05c5097464d6982589f26f4[04]=8448;I7a475a8b0a074fa8bd3bf54dc2a172de8c70f8ad78980010b9d8e9bc5a5b978f[ 4]=14460;A[ 4]=8832;Ibeac5ed31d4582212c21a5dd06959110a37c49046ed23020de290e17d4f45815[ 4]="I65fbe7a0709a36e2f5f6295e0e45fb58ad21e0a3c0f1f5acd39a7a9f2d529f2c";
Idb5f1a085a445a011e36f2e5014265ae744db959b05c5097464d6982589f26f4[05]=8448;I7a475a8b0a074fa8bd3bf54dc2a172de8c70f8ad78980010b9d8e9bc5a5b978f[ 5]=20768;A[ 5]=8832;Ibeac5ed31d4582212c21a5dd06959110a37c49046ed23020de290e17d4f45815[ 5]="I65fbe7a0709a36e2f5f6295e0e45fb58ad21e0a3c0f1f5acd39a7a9f2d529f2c";
Idb5f1a085a445a011e36f2e5014265ae744db959b05c5097464d6982589f26f4[06]=3840;I7a475a8b0a074fa8bd3bf54dc2a172de8c70f8ad78980010b9d8e9bc5a5b978f[ 6]=19200;A[ 6]=4032;Ibeac5ed31d4582212c21a5dd06959110a37c49046ed23020de290e17d4f45815[ 6]="Ic94885c773bb030096af27dd53a4ee4e9113981578431e30e3f1a2e794133a31" ;
Idb5f1a085a445a011e36f2e5014265ae744db959b05c5097464d6982589f26f4[07]=3840;I7a475a8b0a074fa8bd3bf54dc2a172de8c70f8ad78980010b9d8e9bc5a5b978f[ 7]=19200;A[ 7]=4032;Ibeac5ed31d4582212c21a5dd06959110a37c49046ed23020de290e17d4f45815[ 7]="Ic94885c773bb030096af27dd53a4ee4e9113981578431e30e3f1a2e794133a31" ;

Idb5f1a085a445a011e36f2e5014265ae744db959b05c5097464d6982589f26f4[ 8]=8448;I7a475a8b0a074fa8bd3bf54dc2a172de8c70f8ad78980010b9d8e9bc5a5b978f[ 8]=14556;A[ 8]=8832;Ibeac5ed31d4582212c21a5dd06959110a37c49046ed23020de290e17d4f45815[ 8]="I65fbe7a0709a36e2f5f6295e0e45fb58ad21e0a3c0f1f5acd39a7a9f2d529f2c";
Idb5f1a085a445a011e36f2e5014265ae744db959b05c5097464d6982589f26f4[ 9]=8448;I7a475a8b0a074fa8bd3bf54dc2a172de8c70f8ad78980010b9d8e9bc5a5b978f[ 9]=21048;A[ 9]=8832;Ibeac5ed31d4582212c21a5dd06959110a37c49046ed23020de290e17d4f45815[ 9]="I65fbe7a0709a36e2f5f6295e0e45fb58ad21e0a3c0f1f5acd39a7a9f2d529f2c";
Idb5f1a085a445a011e36f2e5014265ae744db959b05c5097464d6982589f26f4[10]=8448;I7a475a8b0a074fa8bd3bf54dc2a172de8c70f8ad78980010b9d8e9bc5a5b978f[10]=25344;A[10]=8832;Ibeac5ed31d4582212c21a5dd06959110a37c49046ed23020de290e17d4f45815[10]="I65fbe7a0709a36e2f5f6295e0e45fb58ad21e0a3c0f1f5acd39a7a9f2d529f2c";
Idb5f1a085a445a011e36f2e5014265ae744db959b05c5097464d6982589f26f4[11]=3840;I7a475a8b0a074fa8bd3bf54dc2a172de8c70f8ad78980010b9d8e9bc5a5b978f[11]=19200;A[11]=4032;Ibeac5ed31d4582212c21a5dd06959110a37c49046ed23020de290e17d4f45815[11]="Ic94885c773bb030096af27dd53a4ee4e9113981578431e30e3f1a2e794133a31" ;


Idb5f1a085a445a011e36f2e5014265ae744db959b05c5097464d6982589f26f4[12]= 501;I7a475a8b0a074fa8bd3bf54dc2a172de8c70f8ad78980010b9d8e9bc5a5b978f[12]= 864 ;A[12]= 546;Ibeac5ed31d4582212c21a5dd06959110a37c49046ed23020de290e17d4f45815[12]="Id6cc51d5d586252100997cbc4eb323c5241e5cf4f9e5348357a7fc8f6a5d9279" ;
Idb5f1a085a445a011e36f2e5014265ae744db959b05c5097464d6982589f26f4[13]= 231;I7a475a8b0a074fa8bd3bf54dc2a172de8c70f8ad78980010b9d8e9bc5a5b978f[13]= 576 ;A[13]= 252;Ibeac5ed31d4582212c21a5dd06959110a37c49046ed23020de290e17d4f45815[13]="Ic52ac15c21ef091ae13a668b6613a4062a8c1fb41806c3b4dfc59f97534d8532"  ;
Idb5f1a085a445a011e36f2e5014265ae744db959b05c5097464d6982589f26f4[14]=  57;I7a475a8b0a074fa8bd3bf54dc2a172de8c70f8ad78980010b9d8e9bc5a5b978f[14]= 288 ;A[14]=  84;Ibeac5ed31d4582212c21a5dd06959110a37c49046ed23020de290e17d4f45815[14]="I03831d3a895200658aa1ddfd4b58cb8ad10c77eef0430b4ee6162279c3015f15"  ;
Idb5f1a085a445a011e36f2e5014265ae744db959b05c5097464d6982589f26f4[15]=  28;I7a475a8b0a074fa8bd3bf54dc2a172de8c70f8ad78980010b9d8e9bc5a5b978f[15]= 140 ;A[15]=  84;Ibeac5ed31d4582212c21a5dd06959110a37c49046ed23020de290e17d4f45815[15]="I03831d3a895200658aa1ddfd4b58cb8ad10c77eef0430b4ee6162279c3015f15"  ;
Idb5f1a085a445a011e36f2e5014265ae744db959b05c5097464d6982589f26f4[16]=1003;I7a475a8b0a074fa8bd3bf54dc2a172de8c70f8ad78980010b9d8e9bc5a5b978f[16]=1728 ;A[16]=1096;Ibeac5ed31d4582212c21a5dd06959110a37c49046ed23020de290e17d4f45815[16]="Id9de73c234dd7a5a70738b2b45c2592cf14d4f946984fbbcfdb024de9c67c457" ;
Idb5f1a085a445a011e36f2e5014265ae744db959b05c5097464d6982589f26f4[17]= 462;I7a475a8b0a074fa8bd3bf54dc2a172de8c70f8ad78980010b9d8e9bc5a5b978f[17]=1152 ;A[17]= 504;Ibeac5ed31d4582212c21a5dd06959110a37c49046ed23020de290e17d4f45815[17]="If3e5687dc8b0205d8fd13e4bd543705974797c428838ee9a7bd83a435c1f10ec" ;
Idb5f1a085a445a011e36f2e5014265ae744db959b05c5097464d6982589f26f4[18]= 115;I7a475a8b0a074fa8bd3bf54dc2a172de8c70f8ad78980010b9d8e9bc5a5b978f[18]= 576 ;A[18]= 126;Ibeac5ed31d4582212c21a5dd06959110a37c49046ed23020de290e17d4f45815[18]="Id328fd565404dc9facd7dacd5efc5261ef9d87fe6ccbb8db46484581b7119bd8"  ;
Idb5f1a085a445a011e36f2e5014265ae744db959b05c5097464d6982589f26f4[19]=  57;I7a475a8b0a074fa8bd3bf54dc2a172de8c70f8ad78980010b9d8e9bc5a5b978f[19]= 286 ;A[19]=  84;Ibeac5ed31d4582212c21a5dd06959110a37c49046ed23020de290e17d4f45815[19]="I03831d3a895200658aa1ddfd4b58cb8ad10c77eef0430b4ee6162279c3015f15"  ;


Idb5f1a085a445a011e36f2e5014265ae744db959b05c5097464d6982589f26f4[20]=8448;I7a475a8b0a074fa8bd3bf54dc2a172de8c70f8ad78980010b9d8e9bc5a5b978f[20]=25344;A[20]=8832;Ibeac5ed31d4582212c21a5dd06959110a37c49046ed23020de290e17d4f45815[20]="I65fbe7a0709a36e2f5f6295e0e45fb58ad21e0a3c0f1f5acd39a7a9f2d529f2c";

Idb5f1a085a445a011e36f2e5014265ae744db959b05c5097464d6982589f26f4[21]=8448;I7a475a8b0a074fa8bd3bf54dc2a172de8c70f8ad78980010b9d8e9bc5a5b978f[21]=14556;A[21]=8832;Ibeac5ed31d4582212c21a5dd06959110a37c49046ed23020de290e17d4f45815[21]="I65fbe7a0709a36e2f5f6295e0e45fb58ad21e0a3c0f1f5acd39a7a9f2d529f2c";
Idb5f1a085a445a011e36f2e5014265ae744db959b05c5097464d6982589f26f4[22]=4162;I7a475a8b0a074fa8bd3bf54dc2a172de8c70f8ad78980010b9d8e9bc5a5b978f[22]=10368;A[22]=4416;Ibeac5ed31d4582212c21a5dd06959110a37c49046ed23020de290e17d4f45815[22]="I2ce9f8f34a8afa13081b150a95333c18679b12f6f8a64cf6f4ab6406accccb7d" ;
Idb5f1a085a445a011e36f2e5014265ae744db959b05c5097464d6982589f26f4[23]=1036;I7a475a8b0a074fa8bd3bf54dc2a172de8c70f8ad78980010b9d8e9bc5a5b978f[23]= 5180;A[23]=1096;Ibeac5ed31d4582212c21a5dd06959110a37c49046ed23020de290e17d4f45815[23]="Id9de73c234dd7a5a70738b2b45c2592cf14d4f946984fbbcfdb024de9c67c457" ;
Idb5f1a085a445a011e36f2e5014265ae744db959b05c5097464d6982589f26f4[24]= 518;I7a475a8b0a074fa8bd3bf54dc2a172de8c70f8ad78980010b9d8e9bc5a5b978f[24]= 2590;A[24]= 546;Ibeac5ed31d4582212c21a5dd06959110a37c49046ed23020de290e17d4f45815[24]="Id6cc51d5d586252100997cbc4eb323c5241e5cf4f9e5348357a7fc8f6a5d9279" ;

Idb5f1a085a445a011e36f2e5014265ae744db959b05c5097464d6982589f26f4[25]=4326;I7a475a8b0a074fa8bd3bf54dc2a172de8c70f8ad78980010b9d8e9bc5a5b978f[25]=4162 ;A[25]=4784;Ibeac5ed31d4582212c21a5dd06959110a37c49046ed23020de290e17d4f45815[25]="Ifcb35d944306ccef07d039274fada0f964cb1a77a01925aa585c25a2e9ecf0df";

Idb5f1a085a445a011e36f2e5014265ae744db959b05c5097464d6982589f26f4[26]=1036;I7a475a8b0a074fa8bd3bf54dc2a172de8c70f8ad78980010b9d8e9bc5a5b978f[26]=5180 ;A[26]=1092;Ibeac5ed31d4582212c21a5dd06959110a37c49046ed23020de290e17d4f45815[26]="Id9de73c234dd7a5a70738b2b45c2592cf14d4f946984fbbcfdb024de9c67c457" ;
Idb5f1a085a445a011e36f2e5014265ae744db959b05c5097464d6982589f26f4[27]=518 ;I7a475a8b0a074fa8bd3bf54dc2a172de8c70f8ad78980010b9d8e9bc5a5b978f[27]=2590 ;A[27]= 546;Ibeac5ed31d4582212c21a5dd06959110a37c49046ed23020de290e17d4f45815[27]="Id6cc51d5d586252100997cbc4eb323c5241e5cf4f9e5348357a7fc8f6a5d9279" ;

end
initial
begin

  automatic int I132ac025db10323da7e56fc77fd857c9f0d0197a23e62b72b3b47b52aae9b32d;
  automatic int I85e4aea19de2d285c91b909a8dcd3d895ad511f5c888998471db1734c996c1ee;
  automatic int Ica16285eedd36a521c6d7d12bbea6ace858611ef6e157d84a52221b529943b79;
  automatic int Ie6490d0ed1fc22607a023c6f727a12fd688ada3cd86530d53a33472e1e6ae6df;
  automatic int Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13 = 0;

  Icced28c6dc3f99c2396a5eaad732bf6b28142335892b1cd0e6af6cdb53f5ccfa                          <= 1'b0;
  Ica16285eedd36a521c6d7d12bbea6ace858611ef6e157d84a52221b529943b79 = 0;

  repeat (1) @ (posedge rstn);
  repeat (10) @ (posedge clk);

  if (I1725d63fa57c5344aa111b908a4770db8738a8217a8d458c8af741a8df7cc480) begin


              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [0] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [1] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [2] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [3] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [4] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [5] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [6] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [7] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [8] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [9] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [10] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [11] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [12] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [13] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [14] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [15] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [16] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [17] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [18] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [19] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [20] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [21] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [22] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [23] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [24] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [25] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [26] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [27] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [28] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [29] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [30] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [31] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [32] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [33] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [34] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [35] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [36] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [37] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [38] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [39] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [40] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [41] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [42] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [43] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [44] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [45] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [46] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [47] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [48] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [49] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [50] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [51] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [52] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [53] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [54] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [55] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [56] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [57] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [58] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [59] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [60] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [61] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [62] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [63] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [64] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [65] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [66] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [67] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [68] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [69] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [70] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [71] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [72] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [73] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [74] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [75] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [76] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [77] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [78] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [79] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [80] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [81] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [82] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [83] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [84] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [85] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [86] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [87] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [88] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [89] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [90] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [91] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [92] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [93] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [94] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [95] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [96] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [97] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [98] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [99] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [100] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [101] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [102] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [103] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [104] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [105] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [106] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [107] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [108] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [109] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [110] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [111] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [112] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [113] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [114] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [115] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [116] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [117] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [118] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [119] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [120] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [121] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [122] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [123] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [124] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [125] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [126] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [127] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [128] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [129] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [130] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [131] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [132] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [133] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [134] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [135] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [136] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [137] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [138] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [139] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [140] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [141] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [142] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [143] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [144] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [145] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [146] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [147] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [148] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [149] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [150] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [151] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [152] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [153] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [154] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [155] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [156] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [157] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [158] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [159] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [160] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [161] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [162] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [163] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [164] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [165] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [166] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [167] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [168] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [169] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [170] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [171] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [172] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [173] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [174] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [175] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [176] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [177] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [178] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [179] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [180] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [181] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [182] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [183] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [184] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [185] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [186] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [187] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [188] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [189] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [190] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [191] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [192] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [193] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [194] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [195] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [196] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [197] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [198] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [199] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [200] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [201] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [202] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [203] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [204] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [205] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [206] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
              I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [207] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                 // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01

         exp_syn [0] <= 1'b1;
         exp_syn [1] <= 1'b1;
         exp_syn [2] <= 1'b1;
         exp_syn [3] <= 1'b1;
         exp_syn [4] <= 1'b1;
         exp_syn [5] <= 1'b1;
         exp_syn [6] <= 1'b1;
         exp_syn [7] <= 1'b1;
         exp_syn [8] <= 1'b1;
         exp_syn [9] <= 1'b1;
         exp_syn [10] <= 1'b1;
         exp_syn [11] <= 1'b1;
         exp_syn [12] <= 1'b1;
         exp_syn [13] <= 1'b1;
         exp_syn [14] <= 1'b1;
         exp_syn [15] <= 1'b1;
         exp_syn [16] <= 1'b1;
         exp_syn [17] <= 1'b1;
         exp_syn [18] <= 1'b1;
         exp_syn [19] <= 1'b1;
         exp_syn [20] <= 1'b1;
         exp_syn [21] <= 1'b1;
         exp_syn [22] <= 1'b1;
         exp_syn [23] <= 1'b1;
         exp_syn [24] <= 1'b1;
         exp_syn [25] <= 1'b1;
         exp_syn [26] <= 1'b1;
         exp_syn [27] <= 1'b1;
         exp_syn [28] <= 1'b1;
         exp_syn [29] <= 1'b1;
         exp_syn [30] <= 1'b1;
         exp_syn [31] <= 1'b1;
         exp_syn [32] <= 1'b1;
         exp_syn [33] <= 1'b1;
         exp_syn [34] <= 1'b1;
         exp_syn [35] <= 1'b1;
         exp_syn [36] <= 1'b1;
         exp_syn [37] <= 1'b1;
         exp_syn [38] <= 1'b1;
         exp_syn [39] <= 1'b1;
         exp_syn [40] <= 1'b1;
         exp_syn [41] <= 1'b1;
         exp_syn [42] <= 1'b1;
         exp_syn [43] <= 1'b1;
         exp_syn [44] <= 1'b1;
         exp_syn [45] <= 1'b1;
         exp_syn [46] <= 1'b1;
         exp_syn [47] <= 1'b1;
         exp_syn [48] <= 1'b1;
         exp_syn [49] <= 1'b1;
         exp_syn [50] <= 1'b1;
         exp_syn [51] <= 1'b1;
         exp_syn [52] <= 1'b1;
         exp_syn [53] <= 1'b1;
         exp_syn [54] <= 1'b1;
         exp_syn [55] <= 1'b1;
         exp_syn [56] <= 1'b1;
         exp_syn [57] <= 1'b1;
         exp_syn [58] <= 1'b1;
         exp_syn [59] <= 1'b1;
         exp_syn [60] <= 1'b1;
         exp_syn [61] <= 1'b1;
         exp_syn [62] <= 1'b1;
         exp_syn [63] <= 1'b1;
         exp_syn [64] <= 1'b1;
         exp_syn [65] <= 1'b1;
         exp_syn [66] <= 1'b1;
         exp_syn [67] <= 1'b1;
         exp_syn [68] <= 1'b1;
         exp_syn [69] <= 1'b1;
         exp_syn [70] <= 1'b1;
         exp_syn [71] <= 1'b1;
         exp_syn [72] <= 1'b1;
         exp_syn [73] <= 1'b1;
         exp_syn [74] <= 1'b1;
         exp_syn [75] <= 1'b1;
         exp_syn [76] <= 1'b1;
         exp_syn [77] <= 1'b1;
         exp_syn [78] <= 1'b1;
         exp_syn [79] <= 1'b1;
         exp_syn [80] <= 1'b1;
         exp_syn [81] <= 1'b1;
         exp_syn [82] <= 1'b1;
         exp_syn [83] <= 1'b1;
         exp_syn [84] <= 1'b1;
         exp_syn [85] <= 1'b1;
         exp_syn [86] <= 1'b1;
         exp_syn [87] <= 1'b1;
         exp_syn [88] <= 1'b1;
         exp_syn [89] <= 1'b1;
         exp_syn [90] <= 1'b1;
         exp_syn [91] <= 1'b1;
         exp_syn [92] <= 1'b1;
         exp_syn [93] <= 1'b1;
         exp_syn [94] <= 1'b1;
         exp_syn [95] <= 1'b1;
         exp_syn [96] <= 1'b1;
         exp_syn [97] <= 1'b1;
         exp_syn [98] <= 1'b1;
         exp_syn [99] <= 1'b1;
         exp_syn [100] <= 1'b1;
         exp_syn [101] <= 1'b1;
         exp_syn [102] <= 1'b1;
         exp_syn [103] <= 1'b1;
         exp_syn [104] <= 1'b1;
         exp_syn [105] <= 1'b1;
         exp_syn [106] <= 1'b1;
         exp_syn [107] <= 1'b1;
         exp_syn [108] <= 1'b1;
         exp_syn [109] <= 1'b1;
         exp_syn [110] <= 1'b1;
         exp_syn [111] <= 1'b1;
         exp_syn [112] <= 1'b1;
         exp_syn [113] <= 1'b1;
         exp_syn [114] <= 1'b1;
         exp_syn [115] <= 1'b1;
         exp_syn [116] <= 1'b1;
         exp_syn [117] <= 1'b1;
         exp_syn [118] <= 1'b1;
         exp_syn [119] <= 1'b1;
         exp_syn [120] <= 1'b1;
         exp_syn [121] <= 1'b1;
         exp_syn [122] <= 1'b1;
         exp_syn [123] <= 1'b1;
         exp_syn [124] <= 1'b1;
         exp_syn [125] <= 1'b1;
         exp_syn [126] <= 1'b1;
         exp_syn [127] <= 1'b1;
         exp_syn [128] <= 1'b1;
         exp_syn [129] <= 1'b1;
         exp_syn [130] <= 1'b1;
         exp_syn [131] <= 1'b1;
         exp_syn [132] <= 1'b1;
         exp_syn [133] <= 1'b1;
         exp_syn [134] <= 1'b1;
         exp_syn [135] <= 1'b1;
         exp_syn [136] <= 1'b1;
         exp_syn [137] <= 1'b1;
         exp_syn [138] <= 1'b1;
         exp_syn [139] <= 1'b1;
         exp_syn [140] <= 1'b1;
         exp_syn [141] <= 1'b1;
         exp_syn [142] <= 1'b1;
         exp_syn [143] <= 1'b1;
         exp_syn [144] <= 1'b1;
         exp_syn [145] <= 1'b1;
         exp_syn [146] <= 1'b1;
         exp_syn [147] <= 1'b1;
         exp_syn [148] <= 1'b1;
         exp_syn [149] <= 1'b1;
         exp_syn [150] <= 1'b1;
         exp_syn [151] <= 1'b1;
         exp_syn [152] <= 1'b1;
         exp_syn [153] <= 1'b1;
         exp_syn [154] <= 1'b1;
         exp_syn [155] <= 1'b1;
         exp_syn [156] <= 1'b1;
         exp_syn [157] <= 1'b1;
         exp_syn [158] <= 1'b1;
         exp_syn [159] <= 1'b1;
         exp_syn [160] <= 1'b1;
         exp_syn [161] <= 1'b1;
         exp_syn [162] <= 1'b1;
         exp_syn [163] <= 1'b1;
         exp_syn [164] <= 1'b1;
         exp_syn [165] <= 1'b1;
         exp_syn [166] <= 1'b1;
         exp_syn [167] <= 1'b1;

  end else begin //I1725d63fa57c5344aa111b908a4770db8738a8217a8d458c8af741a8df7cc480==0
     bit Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf;
         y_nr_in[0] = 1; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[1] = 1; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[2] = 0; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[3] = 1; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[4] = 0; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[5] = 0; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[6] = 0; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[7] = 0; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[8] = 0; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[9] = 1; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[10] = 1; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[11] = 1; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[12] = 1; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[13] = 1; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[14] = 0; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[15] = 1; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[16] = 0; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[17] = 0; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[18] = 1; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[19] = 0; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[20] = 1; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[21] = 1; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[22] = 0; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[23] = 0; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[24] = 0; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[25] = 1; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[26] = 1; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[27] = 0; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[28] = 0; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[29] = 1; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[30] = 1; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[31] = 1; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[32] = 0; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[33] = 0; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[34] = 1; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[35] = 0; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[36] = 0; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[37] = 0; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[38] = 0; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
         y_nr_in[39] = 0; //I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7
     repeat (1) @ (posedge clk);
     for (int Ide7d1b721a1e0632b7cf04edf5032c8ecffa9f9a08492152b926f1a5a7e765d7=0;Ide7d1b721a1e0632b7cf04edf5032c8ecffa9f9a08492152b926f1a5a7e765d7<NN-MM;Ide7d1b721a1e0632b7cf04edf5032c8ecffa9f9a08492152b926f1a5a7e765d7++) begin
         $display("I3a6eb0790f39ac87c94f3856b2dd2c5d110e6811602261a9a923d3bb23adc8b7  y_nr_in [%0d]:%0d I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[%0d]:%0d", Ide7d1b721a1e0632b7cf04edf5032c8ecffa9f9a08492152b926f1a5a7e765d7,y_nr_in [Ide7d1b721a1e0632b7cf04edf5032c8ecffa9f9a08492152b926f1a5a7e765d7],Ide7d1b721a1e0632b7cf04edf5032c8ecffa9f9a08492152b926f1a5a7e765d7,I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[Ide7d1b721a1e0632b7cf04edf5032c8ecffa9f9a08492152b926f1a5a7e765d7]);
     end
     for (int Ide7d1b721a1e0632b7cf04edf5032c8ecffa9f9a08492152b926f1a5a7e765d7=NN-MM;Ide7d1b721a1e0632b7cf04edf5032c8ecffa9f9a08492152b926f1a5a7e765d7<NN;Ide7d1b721a1e0632b7cf04edf5032c8ecffa9f9a08492152b926f1a5a7e765d7++) begin
         $display("I65966f0faeeff2d783a9e9766d96bafb9ce7ea133ccabd263106f6d7ff1ddd14  I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6 [%0d]:%0d", Ide7d1b721a1e0632b7cf04edf5032c8ecffa9f9a08492152b926f1a5a7e765d7,I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6 [Ide7d1b721a1e0632b7cf04edf5032c8ecffa9f9a08492152b926f1a5a7e765d7]);
     end
     //if (~valid_cword)
     //     $fatal (0,"I907d4883cd4a82ba4409064cd83a1659a672e4c392eb0e34bbbc56077d3c0dc6 I20f65c28671b40937c5bf23acc7c6f37e5a5ec0622e347b57685725df5ba9e50 I9ff94c3eb0c1d350b76101c553e6e70c1178b96fc7fd738182e39e2a3f1b9ebe not a valid I5694d08a2e53ffcae0c3103e5ad6f6076abd960eb1f8a56577040bc1028f702b I98c1eb4ee93476743763878fcb96a25fbc9a175074d64004779ecb5242f645e6");
     //else
     //     $info ("Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 a valid I5694d08a2e53ffcae0c3103e5ad6f6076abd960eb1f8a56577040bc1028f702b I98c1eb4ee93476743763878fcb96a25fbc9a175074d64004779ecb5242f645e6");

       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 0, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[0] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[0] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 1, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[1] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[1] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 2, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[2] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[2] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 3, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[3] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[3] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 4, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[4] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[4] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 5, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[5] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[5] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 6, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[6] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[6] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 7, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[7] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[7] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 8, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[8] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[8] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 9, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[9] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[9] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 10, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[10] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[10] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 11, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[11] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[11] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 12, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[12] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[12] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 13, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[13] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[13] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 14, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[14] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[14] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 15, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[15] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[15] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 16, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[16] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[16] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 17, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[17] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[17] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 18, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[18] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[18] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 19, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[19] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[19] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 20, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[20] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[20] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 21, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[21] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[21] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 22, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[22] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[22] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 23, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[23] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[23] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 24, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[24] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[24] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 25, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[25] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[25] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 26, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[26] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[26] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 27, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[27] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[27] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 28, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[28] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[28] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 29, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[29] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[29] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 30, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[30] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[30] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 31, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[31] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[31] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 32, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[32] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[32] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 33, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[33] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[33] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 34, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[34] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[34] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 35, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[35] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[35] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 36, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[36] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[36] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 37, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[37] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[37] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 38, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[38] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[38] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 39, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[39] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[39] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 40, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[40] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[40] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 41, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[41] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[41] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 42, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[42] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[42] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 43, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[43] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[43] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 44, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[44] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[44] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 45, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[45] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[45] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 46, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[46] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[46] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 47, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[47] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[47] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 48, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[48] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[48] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 49, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[49] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[49] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 50, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[50] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[50] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 51, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[51] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[51] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 52, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[52] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[52] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 53, 1,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[53] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[53] ^ 1; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 54, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[54] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[54] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 55, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[55] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[55] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 56, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[56] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[56] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 57, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[57] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[57] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 58, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[58] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[58] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 59, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[59] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[59] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 60, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[60] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[60] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 61, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[61] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[61] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 62, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[62] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[62] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 63, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[63] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[63] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 64, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[64] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[64] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 65, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[65] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[65] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 66, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[66] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[66] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 67, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[67] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[67] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 68, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[68] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[68] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 69, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[69] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[69] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 70, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[70] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[70] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 71, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[71] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[71] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 72, 1,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[72] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[72] ^ 1; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 73, 1,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[73] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[73] ^ 1; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 74, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[74] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[74] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 75, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[75] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[75] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 76, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[76] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[76] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 77, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[77] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[77] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 78, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[78] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[78] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 79, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[79] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[79] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 80, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[80] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[80] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 81, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[81] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[81] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 82, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[82] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[82] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 83, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[83] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[83] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 84, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[84] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[84] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 85, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[85] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[85] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 86, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[86] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[86] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 87, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[87] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[87] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 88, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[88] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[88] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 89, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[89] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[89] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 90, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[90] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[90] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 91, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[91] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[91] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 92, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[92] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[92] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 93, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[93] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[93] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 94, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[94] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[94] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 95, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[95] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[95] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 96, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[96] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[96] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 97, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[97] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[97] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 98, 1,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[98] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[98] ^ 1; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 99, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[99] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[99] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 100, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[100] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[100] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 101, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[101] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[101] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 102, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[102] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[102] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 103, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[103] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[103] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 104, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[104] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[104] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 105, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[105] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[105] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 106, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[106] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[106] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 107, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[107] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[107] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 108, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[108] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[108] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 109, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[109] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[109] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 110, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[110] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[110] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 111, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[111] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[111] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 112, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[112] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[112] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 113, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[113] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[113] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 114, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[114] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[114] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 115, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[115] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[115] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 116, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[116] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[116] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 117, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[117] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[117] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 118, 1,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[118] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[118] ^ 1; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 119, 1,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[119] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[119] ^ 1; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 120, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[120] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[120] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 121, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[121] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[121] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 122, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[122] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[122] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 123, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[123] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[123] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 124, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[124] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[124] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 125, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[125] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[125] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 126, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[126] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[126] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 127, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[127] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[127] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 128, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[128] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[128] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 129, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[129] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[129] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 130, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[130] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[130] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 131, 1,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[131] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[131] ^ 1; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 132, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[132] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[132] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 133, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[133] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[133] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 134, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[134] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[134] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 135, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[135] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[135] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 136, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[136] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[136] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 137, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[137] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[137] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 138, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[138] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[138] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 139, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[139] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[139] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 140, 1,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[140] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[140] ^ 1; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 141, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[141] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[141] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 142, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[142] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[142] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 143, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[143] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[143] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 144, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[144] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[144] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 145, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[145] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[145] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 146, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[146] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[146] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 147, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[147] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[147] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 148, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[148] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[148] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 149, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[149] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[149] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 150, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[150] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[150] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 151, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[151] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[151] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 152, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[152] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[152] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 153, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[153] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[153] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 154, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[154] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[154] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 155, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[155] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[155] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 156, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[156] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[156] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 157, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[157] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[157] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 158, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[158] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[158] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 159, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[159] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[159] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 160, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[160] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[160] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 161, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[161] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[161] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 162, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[162] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[162] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 163, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[163] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[163] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 164, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[164] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[164] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 165, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[165] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[165] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 166, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[166] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[166] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 167, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[167] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[167] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 168, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[168] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[168] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 169, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[169] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[169] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 170, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[170] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[170] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 171, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[171] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[171] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 172, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[172] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[172] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 173, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[173] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[173] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 174, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[174] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[174] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 175, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[175] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[175] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 176, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[176] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[176] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 177, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[177] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[177] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 178, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[178] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[178] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 179, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[179] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[179] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 180, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[180] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[180] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 181, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[181] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[181] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 182, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[182] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[182] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 183, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[183] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[183] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 184, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[184] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[184] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 185, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[185] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[185] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 186, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[186] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[186] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 187, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[187] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[187] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 188, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[188] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[188] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 189, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[189] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[189] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 190, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[190] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[190] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 191, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[191] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[191] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 192, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[192] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[192] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 193, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[193] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[193] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 194, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[194] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[194] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 195, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[195] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[195] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 196, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[196] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[196] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 197, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[197] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[197] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 198, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[198] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[198] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 199, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[199] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[199] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 200, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[200] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[200] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 201, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[201] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[201] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 202, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[202] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[202] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 203, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[203] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[203] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 204, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[204] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[204] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 205, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[205] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[205] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 206, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[206] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[206] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
       $display ("Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 bit [%0d]:%0d I4aa85bde7e5621656ba1fb18520b414e58dd66e0ad07781fd8b278069054242c:%0d", 207, 0,Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13);
       I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[207] = I7135bfe2297853b87558ec0b22b5b3e070b8df3222c1e1930a310474337762e6[207] ^ 0; //Ica00fccfb408989eddc401062c4d1219a6aceb6b9b55412357f1790862e8f178 I86454204b9aa2bcb7aa26de8577832068847a0d922b2218fa2eaa964cac519ec
       Id394af78a21f8f29bdd31648d48de560f9faeed4ad0c1fa29f7e6a12efdf6f13++;
         tmp_bit[0] = 1;
         tmp_bit[1] = 1;
         tmp_bit[2] = 0;
         tmp_bit[3] = 1;
         tmp_bit[4] = 0;
         tmp_bit[5] = 0;
         tmp_bit[6] = 0;
         tmp_bit[7] = 0;
         tmp_bit[8] = 0;
         tmp_bit[9] = 1;
         tmp_bit[10] = 1;
         tmp_bit[11] = 1;
         tmp_bit[12] = 1;
         tmp_bit[13] = 1;
         tmp_bit[14] = 0;
         tmp_bit[15] = 1;
         tmp_bit[16] = 0;
         tmp_bit[17] = 0;
         tmp_bit[18] = 1;
         tmp_bit[19] = 0;
         tmp_bit[20] = 1;
         tmp_bit[21] = 1;
         tmp_bit[22] = 0;
         tmp_bit[23] = 0;
         tmp_bit[24] = 0;
         tmp_bit[25] = 1;
         tmp_bit[26] = 1;
         tmp_bit[27] = 0;
         tmp_bit[28] = 0;
         tmp_bit[29] = 1;
         tmp_bit[30] = 1;
         tmp_bit[31] = 1;
         tmp_bit[32] = 0;
         tmp_bit[33] = 0;
         tmp_bit[34] = 1;
         tmp_bit[35] = 0;
         tmp_bit[36] = 0;
         tmp_bit[37] = 0;
         tmp_bit[38] = 0;
         tmp_bit[39] = 0;
         tmp_bit[40] = 1;
         tmp_bit[41] = 0;
         tmp_bit[42] = 0;
         tmp_bit[43] = 1;
         tmp_bit[44] = 1;
         tmp_bit[45] = 1;
         tmp_bit[46] = 1;
         tmp_bit[47] = 0;
         tmp_bit[48] = 0;
         tmp_bit[49] = 1;
         tmp_bit[50] = 1;
         tmp_bit[51] = 0;
         tmp_bit[52] = 1;
         tmp_bit[53] = 1;
         tmp_bit[54] = 0;
         tmp_bit[55] = 1;
         tmp_bit[56] = 1;
         tmp_bit[57] = 0;
         tmp_bit[58] = 0;
         tmp_bit[59] = 1;
         tmp_bit[60] = 0;
         tmp_bit[61] = 0;
         tmp_bit[62] = 0;
         tmp_bit[63] = 1;
         tmp_bit[64] = 0;
         tmp_bit[65] = 1;
         tmp_bit[66] = 1;
         tmp_bit[67] = 1;
         tmp_bit[68] = 1;
         tmp_bit[69] = 1;
         tmp_bit[70] = 1;
         tmp_bit[71] = 1;
         tmp_bit[72] = 0;
         tmp_bit[73] = 0;
         tmp_bit[74] = 1;
         tmp_bit[75] = 0;
         tmp_bit[76] = 0;
         tmp_bit[77] = 0;
         tmp_bit[78] = 0;
         tmp_bit[79] = 0;
         tmp_bit[80] = 0;
         tmp_bit[81] = 1;
         tmp_bit[82] = 1;
         tmp_bit[83] = 0;
         tmp_bit[84] = 0;
         tmp_bit[85] = 0;
         tmp_bit[86] = 0;
         tmp_bit[87] = 0;
         tmp_bit[88] = 0;
         tmp_bit[89] = 1;
         tmp_bit[90] = 0;
         tmp_bit[91] = 1;
         tmp_bit[92] = 0;
         tmp_bit[93] = 0;
         tmp_bit[94] = 0;
         tmp_bit[95] = 0;
         tmp_bit[96] = 0;
         tmp_bit[97] = 0;
         tmp_bit[98] = 0;
         tmp_bit[99] = 0;
         tmp_bit[100] = 1;
         tmp_bit[101] = 1;
         tmp_bit[102] = 1;
         tmp_bit[103] = 1;
         tmp_bit[104] = 0;
         tmp_bit[105] = 1;
         tmp_bit[106] = 1;
         tmp_bit[107] = 1;
         tmp_bit[108] = 0;
         tmp_bit[109] = 0;
         tmp_bit[110] = 0;
         tmp_bit[111] = 1;
         tmp_bit[112] = 1;
         tmp_bit[113] = 0;
         tmp_bit[114] = 0;
         tmp_bit[115] = 1;
         tmp_bit[116] = 1;
         tmp_bit[117] = 1;
         tmp_bit[118] = 1;
         tmp_bit[119] = 0;
         tmp_bit[120] = 1;
         tmp_bit[121] = 0;
         tmp_bit[122] = 0;
         tmp_bit[123] = 1;
         tmp_bit[124] = 0;
         tmp_bit[125] = 0;
         tmp_bit[126] = 1;
         tmp_bit[127] = 1;
         tmp_bit[128] = 1;
         tmp_bit[129] = 0;
         tmp_bit[130] = 1;
         tmp_bit[131] = 0;
         tmp_bit[132] = 0;
         tmp_bit[133] = 0;
         tmp_bit[134] = 1;
         tmp_bit[135] = 1;
         tmp_bit[136] = 1;
         tmp_bit[137] = 0;
         tmp_bit[138] = 1;
         tmp_bit[139] = 1;
         tmp_bit[140] = 1;
         tmp_bit[141] = 0;
         tmp_bit[142] = 0;
         tmp_bit[143] = 1;
         tmp_bit[144] = 0;
         tmp_bit[145] = 1;
         tmp_bit[146] = 0;
         tmp_bit[147] = 1;
         tmp_bit[148] = 1;
         tmp_bit[149] = 1;
         tmp_bit[150] = 1;
         tmp_bit[151] = 0;
         tmp_bit[152] = 1;
         tmp_bit[153] = 0;
         tmp_bit[154] = 0;
         tmp_bit[155] = 0;
         tmp_bit[156] = 0;
         tmp_bit[157] = 1;
         tmp_bit[158] = 0;
         tmp_bit[159] = 1;
         tmp_bit[160] = 1;
         tmp_bit[161] = 0;
         tmp_bit[162] = 0;
         tmp_bit[163] = 1;
         tmp_bit[164] = 0;
         tmp_bit[165] = 0;
         tmp_bit[166] = 1;
         tmp_bit[167] = 1;
         tmp_bit[168] = 0;
         tmp_bit[169] = 0;
         tmp_bit[170] = 1;
         tmp_bit[171] = 0;
         tmp_bit[172] = 1;
         tmp_bit[173] = 1;
         tmp_bit[174] = 0;
         tmp_bit[175] = 0;
         tmp_bit[176] = 1;
         tmp_bit[177] = 0;
         tmp_bit[178] = 1;
         tmp_bit[179] = 1;
         tmp_bit[180] = 1;
         tmp_bit[181] = 0;
         tmp_bit[182] = 1;
         tmp_bit[183] = 1;
         tmp_bit[184] = 1;
         tmp_bit[185] = 1;
         tmp_bit[186] = 0;
         tmp_bit[187] = 1;
         tmp_bit[188] = 0;
         tmp_bit[189] = 0;
         tmp_bit[190] = 0;
         tmp_bit[191] = 0;
         tmp_bit[192] = 1;
         tmp_bit[193] = 0;
         tmp_bit[194] = 0;
         tmp_bit[195] = 0;
         tmp_bit[196] = 0;
         tmp_bit[197] = 0;
         tmp_bit[198] = 0;
         tmp_bit[199] = 0;
         tmp_bit[200] = 0;
         tmp_bit[201] = 0;
         tmp_bit[202] = 1;
         tmp_bit[203] = 0;
         tmp_bit[204] = 0;
         tmp_bit[205] = 0;
         tmp_bit[206] = 1;
         tmp_bit[207] = 0;
     repeat (1) @ (posedge clk);
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[0] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 0, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 0, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[1] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 1, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 1, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[2] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 2, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 2, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[3] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 3, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 3, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[4] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 4, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 4, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[5] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 5, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 5, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[6] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 6, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 6, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[7] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 7, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 7, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[8] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 8, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 8, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[9] ;
         if ( 1 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 9, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 9, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[10] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 10, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 10, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[11] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 11, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 11, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[12] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 12, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 12, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[13] ;
         if ( 1 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 13, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 13, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[14] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 14, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 14, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[15] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 15, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 15, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[16] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 16, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 16, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[17] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 17, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 17, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[18] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 18, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 18, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[19] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 19, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 19, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[20] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 20, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 20, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[21] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 21, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 21, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[22] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 22, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 22, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[23] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 23, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 23, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[24] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 24, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 24, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[25] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 25, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 25, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[26] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 26, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 26, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[27] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 27, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 27, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[28] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 28, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 28, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[29] ;
         if ( 1 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 29, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 29, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[30] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 30, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 30, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[31] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 31, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 31, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[32] ;
         if ( 1 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 32, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 32, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[33] ;
         if ( 1 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 33, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 33, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[34] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 34, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 34, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[35] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 35, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 35, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[36] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 36, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 36, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[37] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 37, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 37, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[38] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 38, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 38, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[39] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 39, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 39, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[40] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 40, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 40, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[41] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 41, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 41, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[42] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 42, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 42, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[43] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 43, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 43, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[44] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 44, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 44, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[45] ;
         if ( 1 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 45, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 45, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[46] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 46, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 46, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[47] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 47, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 47, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[48] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 48, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 48, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[49] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 49, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 49, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[50] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 50, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 50, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[51] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 51, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 51, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[52] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 52, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 52, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[53] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 53, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 53, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[54] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 54, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 54, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[55] ;
         if ( 1 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 55, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 55, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[56] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 56, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 56, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[57] ;
         if ( 1 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 57, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 57, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[58] ;
         if ( 1 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 58, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 58, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[59] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 59, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 59, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[60] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 60, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 60, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[61] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 61, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 61, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[62] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 62, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 62, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[63] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 63, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 63, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[64] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 64, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 64, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[65] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 65, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 65, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[66] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 66, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 66, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[67] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 67, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 67, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[68] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 68, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 68, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[69] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 69, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 69, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[70] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 70, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 70, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[71] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 71, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 71, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[72] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 72, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 72, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[73] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 73, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 73, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[74] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 74, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 74, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[75] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 75, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 75, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[76] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 76, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 76, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[77] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 77, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 77, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[78] ;
         if ( 1 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 78, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 78, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[79] ;
         if ( 1 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 79, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 79, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[80] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 80, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 80, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[81] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 81, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 81, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[82] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 82, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 82, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[83] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 83, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 83, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[84] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 84, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 84, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[85] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 85, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 85, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[86] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 86, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 86, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[87] ;
         if ( 1 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 87, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 87, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[88] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 88, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 88, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[89] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 89, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 89, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[90] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 90, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 90, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[91] ;
         if ( 1 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 91, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 91, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[92] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 92, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 92, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[93] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 93, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 93, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[94] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 94, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 94, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[95] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 95, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 95, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[96] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 96, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 96, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[97] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 97, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 97, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[98] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 98, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 98, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[99] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 99, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 99, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[100] ;
         if ( 1 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 100, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 100, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[101] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 101, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 101, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[102] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 102, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 102, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[103] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 103, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 103, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[104] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 104, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 104, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[105] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 105, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 105, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[106] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 106, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 106, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[107] ;
         if ( 1 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 107, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 107, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[108] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 108, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 108, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[109] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 109, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 109, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[110] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 110, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 110, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[111] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 111, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 111, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[112] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 112, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 112, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[113] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 113, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 113, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[114] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 114, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 114, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[115] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 115, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 115, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[116] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 116, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 116, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[117] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 117, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 117, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[118] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 118, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 118, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[119] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 119, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 119, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[120] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 120, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 120, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[121] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 121, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 121, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[122] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 122, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 122, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[123] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 123, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 123, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[124] ;
         if ( 1 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 124, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 124, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[125] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 125, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 125, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[126] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 126, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 126, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[127] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 127, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 127, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[128] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 128, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 128, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[129] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 129, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 129, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[130] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 130, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 130, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[131] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 131, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 131, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[132] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 132, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 132, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[133] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 133, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 133, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[134] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 134, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 134, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[135] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 135, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 135, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[136] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 136, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 136, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[137] ;
         if ( 1 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 137, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 137, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[138] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 138, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 138, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[139] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 139, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 139, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[140] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 140, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 140, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[141] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 141, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 141, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[142] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 142, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 142, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[143] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 143, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 143, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[144] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 144, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 144, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[145] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 145, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 145, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[146] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 146, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 146, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[147] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 147, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 147, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[148] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 148, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 148, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[149] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 149, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 149, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[150] ;
         if ( 1 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 150, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 150, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[151] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 151, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 151, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[152] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 152, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 152, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[153] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 153, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 153, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[154] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 154, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 154, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[155] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 155, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 155, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[156] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 156, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 156, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[157] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 157, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 157, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[158] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 158, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 158, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[159] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 159, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 159, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[160] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 160, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 160, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[161] ;
         if ( 1 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 161, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",1, 161, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[162] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 162, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 162, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[163] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 163, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 163, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[164] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 164, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 164, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[165] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 165, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 165, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[166] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 166, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 166, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
         Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf = ~  syndrome[167] ;
         if ( 0 == Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf ) begin
              $display ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 167, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end else begin
              $error   ("syndrome If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:%0d syndrome[%0d]:%0d",0, 167, Ie526c9dc13a701e0d2aa01f12baca17658d8d25bdf6a389463afc7d2b89110bf );
         end
     repeat (1) @ (posedge clk);
     $finish;

     for (int Ide7d1b721a1e0632b7cf04edf5032c8ecffa9f9a08492152b926f1a5a7e765d7=0;Ide7d1b721a1e0632b7cf04edf5032c8ecffa9f9a08492152b926f1a5a7e765d7<NN;Ide7d1b721a1e0632b7cf04edf5032c8ecffa9f9a08492152b926f1a5a7e765d7++) begin
            if (I37998cc284c9701284a5d99b4ce25aa8641fc2fe88907f05a74a38044c7d11fd[Ide7d1b721a1e0632b7cf04edf5032c8ecffa9f9a08492152b926f1a5a7e765d7]) begin
                 I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [Ide7d1b721a1e0632b7cf04edf5032c8ecffa9f9a08492152b926f1a5a7e765d7] <= 2'b11;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 1: -1 === 2'b11
                                    // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 1 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe -1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b11
            end else begin
                 I341c0a3e67c3146720fa1b9504927ece5f5daefadaad467dddfd2ff04ba039be  [Ide7d1b721a1e0632b7cf04edf5032c8ecffa9f9a08492152b926f1a5a7e765d7] <= 2'b01;  // I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a 0: 1  === 2'b01
                                    // Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 0 I70332d559269a27a08e8292a4582b0a39fc98bf0258f70d94e42a5adac26aebe 1 I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 2'b01
            end
     end
     for (int Ide7d1b721a1e0632b7cf04edf5032c8ecffa9f9a08492152b926f1a5a7e765d7=0;Ide7d1b721a1e0632b7cf04edf5032c8ecffa9f9a08492152b926f1a5a7e765d7<MM;Ide7d1b721a1e0632b7cf04edf5032c8ecffa9f9a08492152b926f1a5a7e765d7++) begin
         exp_syn [Ide7d1b721a1e0632b7cf04edf5032c8ecffa9f9a08492152b926f1a5a7e765d7] <= 1'b1;
     end

  end




  repeat (4) @ (posedge clk);
  Icced28c6dc3f99c2396a5eaad732bf6b28142335892b1cd0e6af6cdb53f5ccfa                          <= 1'b1;
  repeat (1) @ (posedge clk);
  Icced28c6dc3f99c2396a5eaad732bf6b28142335892b1cd0e6af6cdb53f5ccfa                          <= 1'b0;
  repeat (20) @(posedge clk);
  $display("Id69a26f56dfc4cead7151d018c424aea7b4152f95aad72fe789e4ea3d643fdd7:I2c9749f9e802d800d52c4b38776251298f8008aff69126f80e1035e350fbdaf6 I8c90cbf5d27d61f534ee012ea472714b0149ee526e43e0903ff7f07ce7ea4758 If77d1bb58da886e3cbeebbf35a0b3d217b003506792268052c6a730fbc5ec9bc :%0d %t", I132ac025db10323da7e56fc77fd857c9f0d0197a23e62b72b3b47b52aae9b32d, $time);
  repeat (20) @(posedge clk);
  $finish();
end


assign percent_probability_int = 32'd 6592;

initial
begin
  repeat (600) @(posedge clk);
end

initial
begin
  forever begin
      if (I16bdee165138010bda1229669cf4bb78831253202a69fa31552c0ac42725776a[1]) begin
         $display("Ie8c3f3d87ee23e76dc8a5f57f060f9a0f6a9a97fd55bb616eaad66fca7fadd1b end I52774637822c236d84ed1e221bb24d9c1840e08c9d3542efd26f16e27ac8c0a2");
         if (I16bdee165138010bda1229669cf4bb78831253202a69fa31552c0ac42725776a[0]) begin
            $display("Ie5a0eb01db902f451cdd2cbde73f951661b461ca445156da47b65b6d7e4b2106: I62c1a97974dfe6848942794be4f2f027b5f4815e1eb76db63a30f0e290b5c1c4 I54caafa49296ec47f1839e46980ed744804fb7b23264bc6801e03af643c5fbf1");
         end else begin
            $error("I02bd349299173f7fdf2dbc983d70961b26d74e6260c3755a058e25f5ee172f98: I62c1a97974dfe6848942794be4f2f027b5f4815e1eb76db63a30f0e290b5c1c4 not I54caafa49296ec47f1839e46980ed744804fb7b23264bc6801e03af643c5fbf1");
         end
         $finish();
      end
      repeat (1) @(posedge clk);
  end
end

`endif




`ifdef ENCRYPT
`endif

endmodule

//C If029c1f097c0b6dc260a6c5304ad63ce886f7b6078deb247e269b295dd8c9555: I5f75057e98eefa9da67b1a59d3d184f5c0315a905ebe0f6ddfe89aef6413c683 I148de9c5a7a44d19e56cd9ae1a554bf67847afb0c58f6e12fa29ac7ddfca9940:0.100000 I3955f8fd92cda2c17a22e4cccf13c595bc7975089af39fd576cb1be59c0b8269:2.197225 percent_probability_int:'d4500

 //I6ede6cac45f64ed08afc0391ecf38a70942e66382fdad32454a8e52bbe5673d2 I59e61154e1a87dffab5b71a93bf419a969a0a85ae8e300adf0c479acfdc2a59c valid I5694d08a2e53ffcae0c3103e5ad6f6076abd960eb1f8a56577040bc1028f702b I98c1eb4ee93476743763878fcb96a25fbc9a175074d64004779ecb5242f645e6
//y_int:
 //44010bdd34c9a17a9dc5c9798ef00a0604fe89b67904e634be0b
//If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:
 //0200400200100008100880c0000680200320002200
//C If029c1f097c0b6dc260a6c5304ad63ce886f7b6078deb247e269b295dd8c9555: I5f75057e98eefa9da67b1a59d3d184f5c0315a905ebe0f6ddfe89aef6413c683 I148de9c5a7a44d19e56cd9ae1a554bf67847afb0c58f6e12fa29ac7ddfca9940:0.038462 I3955f8fd92cda2c17a22e4cccf13c595bc7975089af39fd576cb1be59c0b8269:3.218876 percent_probability_int:'d6592
