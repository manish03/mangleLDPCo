//`include "GF2_LDPC_flogtanh_0x00007_assign_inc.sv"
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00000] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00000] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00001] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00001] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00002] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00003] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00002] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00004] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00005] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00003] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00006] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00007] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00004] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00008] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00009] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00005] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0000a] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0000b] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00006] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0000c] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0000d] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00007] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0000e] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0000f] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00008] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00010] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00011] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00009] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00012] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00013] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0000a] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00014] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00015] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0000b] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00016] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00017] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0000c] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00018] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00019] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0000d] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0001a] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0001b] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0000e] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0001c] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0001d] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0000f] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0001e] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0001f] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00010] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00020] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00021] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00011] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00022] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00023] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00012] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00024] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00025] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00013] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00026] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00027] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00014] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00028] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00029] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00015] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0002a] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0002b] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00016] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0002c] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0002d] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00017] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0002e] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0002f] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00018] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00030] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00031] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00019] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00032] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00033] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0001a] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00034] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00035] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0001b] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00036] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00037] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0001c] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00038] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00039] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0001d] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0003a] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0003b] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0001e] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0003c] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0003d] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0001f] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0003e] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0003f] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00020] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00040] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00041] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00021] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00042] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00043] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00022] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00044] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00045] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00023] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00046] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00047] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00024] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00048] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00049] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00025] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0004a] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0004b] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00026] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0004c] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0004d] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00027] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0004e] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0004f] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00028] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00050] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00051] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00029] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00052] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00053] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0002a] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00054] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00055] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0002b] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00056] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00057] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0002c] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00058] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00059] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0002d] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0005a] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0005b] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0002e] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0005c] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0005d] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0002f] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0005e] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0005f] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00030] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00060] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00061] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00031] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00062] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00063] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00032] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00064] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00065] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00033] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00066] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00067] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00034] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00068] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00069] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00035] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0006a] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00036] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0006c] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0006d] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00037] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0006e] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00038] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00070] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00071] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00039] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00072] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0003a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00074] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0003b] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00076] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00077] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0003c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00078] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0003d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0007a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0003e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0007c] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0003f] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0007e] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0007f] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00040] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00080] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00041] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00082] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00042] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00084] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00043] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00086] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00044] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00088] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00045] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0008a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00046] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0008c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00047] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0008e] ;
//end
//always_comb begin
              Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00048] = 
          (!flogtanh_sel['h00007]) ? 
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00090] : //%
                       I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00091] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00049] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00092] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0004a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00094] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0004b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00096] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0004c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00098] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0004d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0009a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0004e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0009c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0004f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0009e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00050] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000a0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00051] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000a2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00052] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000a4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00053] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000a6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00054] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000a8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00055] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000aa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00056] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000ac] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00057] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000ae] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00058] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000b0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00059] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000b2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0005a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000b4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0005b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000b6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0005c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000b8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0005d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000ba] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0005e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000bc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0005f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000be] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00060] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000c0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00061] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000c2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00062] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000c4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00063] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000c6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00064] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000c8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00065] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000ca] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00066] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000cc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00067] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000ce] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00068] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000d0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00069] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000d2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0006a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000d4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0006b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000d6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0006c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000d8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0006d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000da] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0006e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000dc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0006f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000de] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00070] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000e0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00071] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000e2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00072] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000e4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00073] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000e6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00074] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000e8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00075] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000ea] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00076] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000ec] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00077] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000ee] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00078] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000f0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00079] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000f2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0007a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000f4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0007b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000f6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0007c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000f8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0007d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000fa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0007e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000fc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0007f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000fe] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00080] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00100] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00081] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00102] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00082] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00104] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00083] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00106] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00084] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00108] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00085] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0010a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00086] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0010c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00087] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0010e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00088] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00110] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00089] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00112] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0008a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00114] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0008b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00116] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0008c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00118] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0008d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0011a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0008e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0011c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0008f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0011e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00090] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00120] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00091] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00122] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00092] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00124] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00093] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00126] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00094] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00128] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00095] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0012a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00096] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0012c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00097] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0012e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00098] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00130] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00099] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00132] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0009a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00134] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0009b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00136] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0009c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00138] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0009d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0013a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0009e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0013c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0009f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0013e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000a0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00140] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000a1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00142] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000a2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00144] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000a3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00146] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000a4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00148] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000a5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0014a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000a6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0014c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000a7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0014e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000a8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00150] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000a9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00152] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000aa] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00154] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000ab] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00156] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000ac] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00158] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000ad] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0015a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000ae] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0015c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000af] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0015e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000b0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00160] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000b1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00162] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000b2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00164] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000b3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00166] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000b4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00168] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000b5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0016a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000b6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0016c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000b7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0016e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000b8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00170] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000b9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00172] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000ba] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00174] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000bb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00176] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000bc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00178] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000bd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0017a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000be] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0017c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000bf] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0017e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000c0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00180] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000c1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00182] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000c2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00184] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000c3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00186] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000c4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00188] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000c5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0018a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000c6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0018c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000c7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0018e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000c8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00190] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000c9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00192] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000ca] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00194] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000cb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00196] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000cc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00198] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000cd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0019a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000ce] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0019c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000cf] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0019e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000d0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001a0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000d1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001a2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000d2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001a4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000d3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001a6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000d4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001a8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000d5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001aa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000d6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001ac] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000d7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001ae] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000d8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001b0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000d9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001b2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000da] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001b4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000db] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001b6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000dc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001b8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000dd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001ba] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000de] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001bc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000df] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001be] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000e0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001c0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000e1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001c2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000e2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001c4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000e3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001c6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000e4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001c8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000e5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001ca] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000e6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001cc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000e7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001ce] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000e8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001d0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000e9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001d2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000ea] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001d4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000eb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001d6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000ec] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001d8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000ed] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001da] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000ee] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001dc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000ef] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001de] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000f0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001e0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000f1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001e2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000f2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001e4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000f3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001e6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000f4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001e8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000f5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001ea] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000f6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001ec] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000f7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001ee] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000f8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001f0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000f9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001f2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000fa] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001f4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000fb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001f6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000fc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001f8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000fd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001fa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000fe] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001fc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000ff] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001fe] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00100] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00200] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00101] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00202] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00102] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00204] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00103] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00206] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00104] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00208] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00105] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0020a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00106] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0020c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00107] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0020e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00108] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00210] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00109] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00212] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0010a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00214] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0010b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00216] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0010c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00218] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0010d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0021a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0010e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0021c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0010f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0021e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00110] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00220] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00111] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00222] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00112] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00224] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00113] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00226] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00114] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00228] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00115] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0022a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00116] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0022c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00117] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0022e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00118] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00230] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00119] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00232] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0011a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00234] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0011b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00236] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0011c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00238] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0011d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0023a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0011e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0023c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0011f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0023e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00120] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00240] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00121] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00242] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00122] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00244] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00123] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00246] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00124] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00248] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00125] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0024a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00126] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0024c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00127] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0024e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00128] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00250] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00129] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00252] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0012a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00254] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0012b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00256] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0012c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00258] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0012d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0025a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0012e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0025c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0012f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0025e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00130] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00260] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00131] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00262] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00132] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00264] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00133] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00266] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00134] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00268] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00135] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0026a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00136] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0026c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00137] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0026e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00138] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00270] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00139] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00272] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0013a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00274] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0013b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00276] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0013c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00278] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0013d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0027a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0013e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0027c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0013f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0027e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00140] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00280] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00141] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00282] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00142] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00284] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00143] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00286] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00144] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00288] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00145] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0028a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00146] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0028c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00147] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0028e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00148] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00290] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00149] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00292] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0014a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00294] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0014b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00296] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0014c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00298] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0014d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0029a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0014e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0029c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0014f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0029e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00150] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002a0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00151] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002a2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00152] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002a4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00153] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002a6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00154] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002a8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00155] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002aa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00156] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002ac] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00157] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002ae] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00158] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002b0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00159] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002b2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0015a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002b4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0015b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002b6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0015c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002b8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0015d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002ba] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0015e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002bc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0015f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002be] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00160] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002c0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00161] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002c2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00162] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002c4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00163] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002c6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00164] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002c8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00165] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002ca] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00166] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002cc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00167] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002ce] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00168] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002d0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00169] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002d2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0016a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002d4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0016b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002d6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0016c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002d8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0016d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002da] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0016e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002dc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0016f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002de] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00170] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002e0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00171] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002e2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00172] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002e4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00173] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002e6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00174] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002e8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00175] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002ea] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00176] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002ec] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00177] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002ee] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00178] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002f0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00179] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002f2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0017a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002f4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0017b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002f6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0017c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002f8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0017d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002fa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0017e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002fc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0017f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002fe] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00180] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00300] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00181] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00302] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00182] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00304] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00183] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00306] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00184] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00308] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00185] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0030a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00186] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0030c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00187] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0030e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00188] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00310] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00189] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00312] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0018a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00314] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0018b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00316] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0018c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00318] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0018d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0031a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0018e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0031c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0018f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0031e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00190] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00320] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00191] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00322] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00192] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00324] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00193] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00326] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00194] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00328] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00195] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0032a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00196] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0032c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00197] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0032e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00198] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00330] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00199] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00332] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0019a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00334] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0019b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00336] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0019c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00338] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0019d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0033a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0019e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0033c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0019f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0033e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001a0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00340] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001a1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00342] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001a2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00344] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001a3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00346] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001a4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00348] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001a5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0034a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001a6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0034c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001a7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0034e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001a8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00350] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001a9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00352] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001aa] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00354] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001ab] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00356] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001ac] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00358] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001ad] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0035a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001ae] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0035c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001af] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0035e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001b0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00360] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001b1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00362] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001b2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00364] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001b3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00366] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001b4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00368] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001b5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0036a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001b6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0036c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001b7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0036e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001b8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00370] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001b9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00372] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001ba] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00374] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001bb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00376] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001bc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00378] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001bd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0037a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001be] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0037c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001bf] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0037e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001c0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00380] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001c1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00382] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001c2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00384] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001c3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00386] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001c4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00388] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001c5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0038a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001c6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0038c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001c7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0038e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001c8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00390] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001c9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00392] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001ca] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00394] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001cb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00396] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001cc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00398] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001cd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0039a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001ce] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0039c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001cf] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0039e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001d0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003a0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001d1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003a2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001d2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003a4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001d3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003a6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001d4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003a8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001d5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003aa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001d6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003ac] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001d7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003ae] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001d8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003b0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001d9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003b2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001da] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003b4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001db] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003b6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001dc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003b8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001dd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003ba] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001de] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003bc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001df] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003be] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001e0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003c0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001e1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003c2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001e2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003c4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001e3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003c6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001e4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003c8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001e5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003ca] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001e6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003cc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001e7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003ce] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001e8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003d0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001e9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003d2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001ea] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003d4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001eb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003d6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001ec] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003d8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001ed] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003da] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001ee] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003dc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001ef] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003de] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001f0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003e0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001f1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003e2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001f2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003e4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001f3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003e6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001f4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003e8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001f5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003ea] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001f6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003ec] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001f7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003ee] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001f8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003f0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001f9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003f2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001fa] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003f4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001fb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003f6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001fc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003f8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001fd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003fa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001fe] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003fc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001ff] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003fe] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00200] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00400] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00201] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00402] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00202] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00404] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00203] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00406] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00204] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00408] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00205] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0040a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00206] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0040c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00207] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0040e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00208] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00410] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00209] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00412] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0020a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00414] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0020b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00416] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0020c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00418] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0020d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0041a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0020e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0041c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0020f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0041e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00210] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00420] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00211] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00422] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00212] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00424] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00213] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00426] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00214] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00428] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00215] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0042a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00216] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0042c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00217] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0042e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00218] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00430] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00219] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00432] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0021a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00434] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0021b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00436] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0021c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00438] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0021d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0043a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0021e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0043c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0021f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0043e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00220] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00440] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00221] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00442] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00222] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00444] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00223] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00446] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00224] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00448] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00225] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0044a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00226] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0044c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00227] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0044e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00228] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00450] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00229] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00452] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0022a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00454] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0022b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00456] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0022c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00458] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0022d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0045a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0022e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0045c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0022f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0045e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00230] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00460] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00231] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00462] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00232] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00464] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00233] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00466] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00234] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00468] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00235] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0046a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00236] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0046c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00237] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0046e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00238] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00470] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00239] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00472] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0023a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00474] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0023b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00476] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0023c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00478] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0023d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0047a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0023e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0047c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0023f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0047e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00240] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00480] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00241] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00482] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00242] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00484] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00243] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00486] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00244] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00488] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00245] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0048a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00246] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0048c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00247] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0048e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00248] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00490] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00249] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00492] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0024a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00494] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0024b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00496] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0024c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00498] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0024d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0049a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0024e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0049c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0024f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0049e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00250] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004a0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00251] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004a2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00252] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004a4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00253] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004a6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00254] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004a8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00255] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004aa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00256] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004ac] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00257] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004ae] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00258] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004b0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00259] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004b2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0025a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004b4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0025b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004b6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0025c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004b8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0025d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004ba] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0025e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004bc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0025f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004be] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00260] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004c0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00261] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004c2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00262] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004c4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00263] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004c6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00264] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004c8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00265] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004ca] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00266] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004cc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00267] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004ce] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00268] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004d0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00269] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004d2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0026a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004d4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0026b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004d6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0026c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004d8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0026d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004da] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0026e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004dc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0026f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004de] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00270] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004e0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00271] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004e2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00272] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004e4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00273] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004e6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00274] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004e8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00275] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004ea] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00276] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004ec] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00277] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004ee] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00278] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004f0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00279] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004f2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0027a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004f4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0027b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004f6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0027c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004f8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0027d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004fa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0027e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004fc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0027f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004fe] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00280] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00500] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00281] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00502] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00282] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00504] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00283] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00506] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00284] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00508] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00285] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0050a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00286] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0050c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00287] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0050e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00288] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00510] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00289] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00512] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0028a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00514] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0028b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00516] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0028c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00518] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0028d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0051a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0028e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0051c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0028f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0051e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00290] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00520] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00291] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00522] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00292] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00524] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00293] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00526] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00294] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00528] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00295] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0052a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00296] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0052c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00297] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0052e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00298] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00530] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00299] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00532] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0029a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00534] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0029b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00536] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0029c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00538] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0029d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0053a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0029e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0053c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0029f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0053e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002a0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00540] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002a1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00542] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002a2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00544] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002a3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00546] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002a4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00548] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002a5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0054a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002a6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0054c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002a7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0054e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002a8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00550] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002a9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00552] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002aa] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00554] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002ab] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00556] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002ac] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00558] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002ad] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0055a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002ae] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0055c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002af] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0055e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002b0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00560] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002b1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00562] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002b2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00564] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002b3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00566] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002b4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00568] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002b5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0056a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002b6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0056c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002b7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0056e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002b8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00570] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002b9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00572] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002ba] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00574] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002bb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00576] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002bc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00578] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002bd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0057a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002be] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0057c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002bf] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0057e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002c0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00580] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002c1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00582] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002c2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00584] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002c3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00586] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002c4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00588] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002c5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0058a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002c6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0058c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002c7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0058e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002c8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00590] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002c9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00592] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002ca] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00594] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002cb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00596] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002cc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00598] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002cd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0059a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002ce] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0059c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002cf] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0059e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002d0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005a0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002d1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005a2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002d2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005a4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002d3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005a6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002d4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005a8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002d5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005aa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002d6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005ac] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002d7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005ae] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002d8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005b0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002d9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005b2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002da] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005b4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002db] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005b6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002dc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005b8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002dd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005ba] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002de] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005bc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002df] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005be] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002e0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005c0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002e1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005c2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002e2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005c4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002e3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005c6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002e4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005c8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002e5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005ca] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002e6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005cc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002e7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005ce] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002e8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005d0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002e9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005d2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002ea] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005d4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002eb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005d6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002ec] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005d8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002ed] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005da] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002ee] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005dc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002ef] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005de] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002f0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005e0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002f1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005e2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002f2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005e4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002f3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005e6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002f4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005e8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002f5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005ea] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002f6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005ec] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002f7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005ee] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002f8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005f0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002f9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005f2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002fa] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005f4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002fb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005f6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002fc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005f8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002fd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005fa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002fe] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005fc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002ff] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005fe] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00300] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00600] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00301] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00602] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00302] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00604] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00303] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00606] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00304] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00608] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00305] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0060a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00306] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0060c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00307] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0060e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00308] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00610] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00309] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00612] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0030a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00614] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0030b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00616] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0030c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00618] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0030d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0061a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0030e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0061c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0030f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0061e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00310] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00620] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00311] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00622] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00312] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00624] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00313] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00626] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00314] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00628] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00315] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0062a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00316] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0062c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00317] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0062e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00318] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00630] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00319] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00632] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0031a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00634] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0031b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00636] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0031c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00638] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0031d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0063a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0031e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0063c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0031f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0063e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00320] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00640] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00321] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00642] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00322] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00644] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00323] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00646] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00324] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00648] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00325] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0064a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00326] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0064c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00327] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0064e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00328] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00650] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00329] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00652] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0032a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00654] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0032b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00656] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0032c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00658] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0032d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0065a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0032e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0065c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0032f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0065e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00330] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00660] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00331] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00662] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00332] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00664] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00333] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00666] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00334] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00668] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00335] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0066a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00336] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0066c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00337] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0066e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00338] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00670] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00339] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00672] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0033a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00674] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0033b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00676] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0033c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00678] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0033d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0067a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0033e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0067c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0033f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0067e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00340] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00680] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00341] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00682] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00342] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00684] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00343] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00686] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00344] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00688] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00345] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0068a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00346] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0068c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00347] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0068e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00348] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00690] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00349] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00692] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0034a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00694] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0034b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00696] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0034c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00698] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0034d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0069a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0034e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0069c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0034f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0069e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00350] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006a0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00351] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006a2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00352] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006a4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00353] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006a6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00354] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006a8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00355] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006aa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00356] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006ac] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00357] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006ae] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00358] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006b0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00359] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006b2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0035a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006b4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0035b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006b6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0035c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006b8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0035d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006ba] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0035e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006bc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0035f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006be] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00360] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006c0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00361] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006c2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00362] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006c4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00363] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006c6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00364] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006c8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00365] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006ca] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00366] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006cc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00367] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006ce] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00368] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006d0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00369] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006d2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0036a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006d4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0036b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006d6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0036c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006d8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0036d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006da] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0036e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006dc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0036f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006de] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00370] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006e0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00371] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006e2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00372] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006e4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00373] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006e6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00374] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006e8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00375] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006ea] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00376] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006ec] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00377] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006ee] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00378] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006f0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00379] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006f2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0037a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006f4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0037b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006f6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0037c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006f8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0037d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006fa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0037e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006fc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0037f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006fe] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00380] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00700] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00381] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00702] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00382] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00704] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00383] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00706] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00384] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00708] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00385] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0070a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00386] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0070c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00387] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0070e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00388] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00710] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00389] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00712] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0038a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00714] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0038b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00716] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0038c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00718] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0038d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0071a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0038e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0071c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0038f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0071e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00390] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00720] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00391] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00722] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00392] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00724] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00393] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00726] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00394] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00728] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00395] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0072a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00396] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0072c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00397] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0072e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00398] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00730] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00399] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00732] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0039a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00734] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0039b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00736] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0039c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00738] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0039d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0073a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0039e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0073c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0039f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0073e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003a0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00740] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003a1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00742] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003a2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00744] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003a3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00746] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003a4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00748] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003a5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0074a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003a6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0074c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003a7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0074e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003a8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00750] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003a9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00752] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003aa] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00754] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003ab] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00756] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003ac] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00758] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003ad] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0075a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003ae] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0075c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003af] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0075e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003b0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00760] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003b1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00762] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003b2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00764] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003b3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00766] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003b4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00768] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003b5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0076a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003b6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0076c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003b7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0076e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003b8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00770] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003b9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00772] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003ba] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00774] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003bb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00776] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003bc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00778] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003bd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0077a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003be] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0077c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003bf] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0077e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003c0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00780] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003c1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00782] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003c2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00784] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003c3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00786] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003c4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00788] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003c5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0078a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003c6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0078c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003c7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0078e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003c8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00790] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003c9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00792] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003ca] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00794] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003cb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00796] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003cc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00798] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003cd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0079a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003ce] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0079c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003cf] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0079e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003d0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007a0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003d1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007a2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003d2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007a4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003d3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007a6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003d4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007a8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003d5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007aa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003d6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007ac] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003d7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007ae] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003d8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007b0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003d9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007b2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003da] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007b4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003db] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007b6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003dc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007b8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003dd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007ba] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003de] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007bc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003df] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007be] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003e0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007c0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003e1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007c2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003e2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007c4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003e3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007c6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003e4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007c8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003e5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007ca] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003e6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007cc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003e7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007ce] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003e8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007d0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003e9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007d2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003ea] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007d4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003eb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007d6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003ec] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007d8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003ed] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007da] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003ee] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007dc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003ef] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007de] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003f0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007e0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003f1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007e2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003f2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007e4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003f3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007e6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003f4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007e8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003f5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007ea] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003f6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007ec] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003f7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007ee] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003f8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007f0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003f9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007f2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003fa] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007f4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003fb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007f6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003fc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007f8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003fd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007fa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003fe] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007fc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003ff] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007fe] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00400] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00800] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00401] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00802] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00402] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00804] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00403] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00806] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00404] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00808] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00405] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0080a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00406] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0080c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00407] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0080e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00408] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00810] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00409] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00812] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0040a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00814] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0040b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00816] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0040c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00818] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0040d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0081a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0040e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0081c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0040f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0081e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00410] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00820] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00411] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00822] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00412] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00824] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00413] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00826] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00414] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00828] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00415] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0082a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00416] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0082c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00417] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0082e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00418] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00830] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00419] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00832] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0041a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00834] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0041b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00836] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0041c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00838] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0041d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0083a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0041e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0083c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0041f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0083e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00420] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00840] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00421] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00842] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00422] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00844] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00423] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00846] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00424] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00848] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00425] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0084a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00426] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0084c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00427] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0084e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00428] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00850] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00429] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00852] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0042a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00854] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0042b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00856] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0042c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00858] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0042d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0085a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0042e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0085c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0042f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0085e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00430] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00860] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00431] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00862] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00432] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00864] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00433] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00866] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00434] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00868] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00435] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0086a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00436] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0086c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00437] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0086e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00438] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00870] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00439] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00872] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0043a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00874] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0043b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00876] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0043c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00878] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0043d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0087a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0043e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0087c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0043f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0087e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00440] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00880] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00441] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00882] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00442] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00884] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00443] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00886] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00444] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00888] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00445] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0088a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00446] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0088c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00447] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0088e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00448] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00890] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00449] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00892] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0044a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00894] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0044b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00896] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0044c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00898] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0044d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0089a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0044e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0089c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0044f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0089e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00450] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008a0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00451] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008a2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00452] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008a4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00453] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008a6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00454] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008a8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00455] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008aa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00456] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008ac] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00457] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008ae] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00458] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008b0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00459] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008b2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0045a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008b4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0045b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008b6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0045c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008b8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0045d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008ba] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0045e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008bc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0045f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008be] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00460] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008c0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00461] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008c2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00462] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008c4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00463] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008c6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00464] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008c8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00465] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008ca] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00466] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008cc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00467] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008ce] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00468] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008d0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00469] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008d2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0046a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008d4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0046b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008d6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0046c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008d8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0046d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008da] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0046e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008dc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0046f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008de] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00470] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008e0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00471] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008e2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00472] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008e4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00473] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008e6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00474] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008e8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00475] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008ea] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00476] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008ec] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00477] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008ee] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00478] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008f0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00479] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008f2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0047a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008f4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0047b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008f6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0047c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008f8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0047d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008fa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0047e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008fc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0047f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008fe] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00480] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00900] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00481] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00902] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00482] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00904] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00483] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00906] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00484] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00908] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00485] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0090a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00486] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0090c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00487] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0090e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00488] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00910] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00489] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00912] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0048a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00914] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0048b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00916] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0048c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00918] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0048d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0091a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0048e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0091c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0048f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0091e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00490] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00920] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00491] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00922] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00492] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00924] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00493] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00926] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00494] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00928] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00495] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0092a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00496] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0092c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00497] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0092e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00498] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00930] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00499] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00932] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0049a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00934] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0049b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00936] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0049c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00938] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0049d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0093a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0049e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0093c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0049f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0093e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004a0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00940] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004a1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00942] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004a2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00944] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004a3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00946] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004a4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00948] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004a5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0094a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004a6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0094c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004a7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0094e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004a8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00950] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004a9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00952] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004aa] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00954] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004ab] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00956] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004ac] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00958] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004ad] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0095a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004ae] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0095c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004af] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0095e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004b0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00960] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004b1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00962] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004b2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00964] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004b3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00966] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004b4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00968] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004b5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0096a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004b6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0096c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004b7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0096e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004b8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00970] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004b9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00972] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004ba] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00974] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004bb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00976] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004bc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00978] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004bd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0097a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004be] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0097c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004bf] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0097e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004c0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00980] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004c1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00982] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004c2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00984] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004c3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00986] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004c4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00988] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004c5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0098a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004c6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0098c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004c7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0098e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004c8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00990] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004c9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00992] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004ca] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00994] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004cb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00996] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004cc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00998] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004cd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0099a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004ce] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0099c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004cf] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0099e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004d0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009a0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004d1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009a2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004d2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009a4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004d3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009a6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004d4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009a8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004d5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009aa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004d6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009ac] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004d7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009ae] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004d8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009b0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004d9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009b2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004da] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009b4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004db] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009b6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004dc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009b8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004dd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009ba] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004de] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009bc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004df] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009be] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004e0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009c0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004e1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009c2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004e2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009c4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004e3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009c6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004e4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009c8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004e5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009ca] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004e6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009cc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004e7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009ce] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004e8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009d0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004e9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009d2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004ea] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009d4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004eb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009d6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004ec] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009d8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004ed] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009da] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004ee] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009dc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004ef] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009de] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004f0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009e0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004f1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009e2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004f2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009e4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004f3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009e6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004f4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009e8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004f5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009ea] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004f6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009ec] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004f7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009ee] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004f8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009f0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004f9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009f2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004fa] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009f4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004fb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009f6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004fc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009f8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004fd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009fa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004fe] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009fc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004ff] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009fe] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00500] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a00] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00501] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a02] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00502] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a04] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00503] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a06] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00504] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a08] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00505] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a0a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00506] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a0c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00507] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a0e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00508] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a10] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00509] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a12] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0050a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a14] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0050b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a16] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0050c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a18] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0050d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a1a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0050e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a1c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0050f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a1e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00510] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a20] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00511] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a22] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00512] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a24] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00513] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a26] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00514] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a28] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00515] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a2a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00516] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a2c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00517] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a2e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00518] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a30] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00519] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a32] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0051a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a34] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0051b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a36] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0051c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a38] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0051d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a3a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0051e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a3c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0051f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a3e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00520] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a40] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00521] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a42] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00522] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a44] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00523] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a46] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00524] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a48] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00525] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a4a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00526] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a4c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00527] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a4e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00528] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a50] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00529] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a52] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0052a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a54] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0052b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a56] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0052c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a58] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0052d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a5a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0052e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a5c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0052f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a5e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00530] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a60] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00531] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a62] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00532] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a64] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00533] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a66] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00534] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a68] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00535] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a6a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00536] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a6c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00537] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a6e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00538] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a70] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00539] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a72] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0053a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a74] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0053b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a76] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0053c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a78] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0053d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a7a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0053e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a7c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0053f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a7e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00540] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a80] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00541] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a82] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00542] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a84] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00543] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a86] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00544] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a88] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00545] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a8a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00546] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a8c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00547] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a8e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00548] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a90] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00549] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a92] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0054a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a94] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0054b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a96] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0054c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a98] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0054d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a9a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0054e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a9c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0054f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a9e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00550] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aa0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00551] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aa2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00552] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aa4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00553] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aa6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00554] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aa8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00555] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aaa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00556] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aac] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00557] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aae] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00558] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ab0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00559] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ab2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0055a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ab4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0055b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ab6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0055c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ab8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0055d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aba] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0055e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00abc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0055f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00abe] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00560] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ac0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00561] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ac2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00562] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ac4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00563] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ac6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00564] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ac8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00565] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aca] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00566] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00acc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00567] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ace] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00568] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ad0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00569] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ad2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0056a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ad4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0056b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ad6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0056c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ad8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0056d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ada] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0056e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00adc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0056f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ade] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00570] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ae0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00571] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ae2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00572] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ae4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00573] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ae6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00574] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ae8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00575] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aea] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00576] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aec] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00577] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aee] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00578] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00af0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00579] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00af2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0057a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00af4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0057b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00af6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0057c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00af8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0057d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00afa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0057e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00afc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0057f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00afe] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00580] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b00] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00581] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b02] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00582] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b04] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00583] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b06] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00584] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b08] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00585] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b0a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00586] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b0c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00587] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b0e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00588] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b10] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00589] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b12] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0058a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b14] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0058b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b16] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0058c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b18] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0058d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b1a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0058e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b1c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0058f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b1e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00590] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b20] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00591] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b22] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00592] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b24] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00593] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b26] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00594] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b28] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00595] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b2a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00596] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b2c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00597] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b2e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00598] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b30] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00599] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b32] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0059a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b34] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0059b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b36] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0059c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b38] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0059d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b3a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0059e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b3c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0059f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b3e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005a0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b40] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005a1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b42] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005a2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b44] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005a3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b46] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005a4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b48] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005a5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b4a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005a6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b4c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005a7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b4e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005a8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b50] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005a9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b52] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005aa] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b54] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005ab] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b56] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005ac] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b58] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005ad] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b5a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005ae] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b5c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005af] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b5e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005b0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b60] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005b1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b62] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005b2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b64] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005b3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b66] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005b4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b68] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005b5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b6a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005b6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b6c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005b7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b6e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005b8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b70] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005b9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b72] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005ba] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b74] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005bb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b76] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005bc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b78] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005bd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b7a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005be] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b7c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005bf] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b7e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005c0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b80] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005c1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b82] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005c2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b84] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005c3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b86] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005c4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b88] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005c5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b8a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005c6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b8c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005c7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b8e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005c8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b90] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005c9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b92] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005ca] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b94] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005cb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b96] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005cc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b98] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005cd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b9a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005ce] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b9c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005cf] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b9e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005d0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ba0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005d1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ba2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005d2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ba4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005d3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ba6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005d4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ba8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005d5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00baa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005d6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bac] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005d7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bae] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005d8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bb0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005d9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bb2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005da] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bb4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005db] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bb6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005dc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bb8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005dd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bba] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005de] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bbc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005df] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bbe] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005e0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bc0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005e1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bc2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005e2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bc4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005e3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bc6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005e4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bc8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005e5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bca] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005e6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bcc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005e7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bce] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005e8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bd0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005e9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bd2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005ea] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bd4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005eb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bd6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005ec] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bd8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005ed] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bda] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005ee] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bdc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005ef] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bde] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005f0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00be0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005f1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00be2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005f2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00be4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005f3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00be6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005f4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00be8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005f5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bea] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005f6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bec] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005f7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bee] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005f8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bf0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005f9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bf2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005fa] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bf4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005fb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bf6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005fc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bf8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005fd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bfa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005fe] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bfc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005ff] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bfe] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00600] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c00] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00601] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c02] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00602] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c04] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00603] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c06] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00604] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c08] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00605] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c0a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00606] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c0c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00607] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c0e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00608] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c10] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00609] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c12] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0060a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c14] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0060b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c16] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0060c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c18] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0060d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c1a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0060e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c1c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0060f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c1e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00610] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c20] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00611] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c22] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00612] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c24] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00613] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c26] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00614] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c28] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00615] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c2a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00616] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c2c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00617] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c2e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00618] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c30] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00619] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c32] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0061a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c34] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0061b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c36] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0061c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c38] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0061d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c3a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0061e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c3c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0061f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c3e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00620] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c40] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00621] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c42] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00622] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c44] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00623] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c46] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00624] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c48] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00625] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c4a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00626] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c4c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00627] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c4e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00628] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c50] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00629] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c52] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0062a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c54] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0062b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c56] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0062c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c58] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0062d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c5a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0062e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c5c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0062f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c5e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00630] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c60] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00631] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c62] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00632] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c64] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00633] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c66] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00634] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c68] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00635] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c6a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00636] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c6c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00637] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c6e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00638] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c70] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00639] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c72] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0063a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c74] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0063b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c76] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0063c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c78] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0063d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c7a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0063e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c7c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0063f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c7e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00640] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c80] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00641] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c82] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00642] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c84] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00643] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c86] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00644] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c88] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00645] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c8a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00646] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c8c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00647] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c8e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00648] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c90] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00649] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c92] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0064a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c94] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0064b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c96] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0064c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c98] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0064d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c9a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0064e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c9c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0064f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c9e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00650] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ca0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00651] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ca2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00652] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ca4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00653] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ca6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00654] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ca8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00655] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00caa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00656] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cac] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00657] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cae] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00658] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cb0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00659] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cb2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0065a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cb4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0065b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cb6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0065c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cb8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0065d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cba] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0065e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cbc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0065f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cbe] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00660] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cc0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00661] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cc2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00662] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cc4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00663] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cc6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00664] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cc8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00665] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cca] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00666] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ccc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00667] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cce] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00668] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cd0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00669] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cd2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0066a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cd4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0066b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cd6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0066c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cd8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0066d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cda] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0066e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cdc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0066f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cde] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00670] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ce0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00671] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ce2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00672] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ce4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00673] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ce6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00674] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ce8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00675] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cea] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00676] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cec] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00677] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cee] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00678] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cf0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00679] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cf2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0067a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cf4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0067b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cf6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0067c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cf8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0067d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cfa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0067e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cfc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0067f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cfe] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00680] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d00] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00681] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d02] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00682] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d04] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00683] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d06] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00684] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d08] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00685] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d0a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00686] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d0c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00687] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d0e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00688] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d10] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00689] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d12] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0068a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d14] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0068b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d16] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0068c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d18] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0068d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d1a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0068e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d1c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0068f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d1e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00690] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d20] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00691] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d22] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00692] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d24] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00693] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d26] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00694] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d28] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00695] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d2a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00696] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d2c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00697] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d2e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00698] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d30] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00699] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d32] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0069a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d34] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0069b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d36] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0069c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d38] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0069d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d3a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0069e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d3c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0069f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d3e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006a0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d40] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006a1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d42] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006a2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d44] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006a3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d46] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006a4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d48] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006a5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d4a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006a6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d4c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006a7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d4e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006a8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d50] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006a9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d52] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006aa] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d54] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006ab] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d56] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006ac] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d58] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006ad] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d5a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006ae] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d5c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006af] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d5e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006b0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d60] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006b1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d62] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006b2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d64] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006b3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d66] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006b4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d68] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006b5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d6a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006b6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d6c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006b7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d6e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006b8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d70] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006b9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d72] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006ba] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d74] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006bb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d76] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006bc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d78] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006bd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d7a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006be] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d7c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006bf] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d7e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006c0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d80] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006c1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d82] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006c2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d84] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006c3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d86] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006c4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d88] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006c5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d8a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006c6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d8c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006c7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d8e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006c8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d90] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006c9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d92] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006ca] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d94] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006cb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d96] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006cc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d98] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006cd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d9a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006ce] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d9c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006cf] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d9e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006d0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00da0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006d1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00da2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006d2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00da4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006d3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00da6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006d4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00da8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006d5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00daa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006d6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dac] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006d7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dae] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006d8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00db0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006d9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00db2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006da] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00db4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006db] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00db6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006dc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00db8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006dd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dba] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006de] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dbc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006df] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dbe] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006e0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dc0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006e1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dc2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006e2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dc4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006e3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dc6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006e4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dc8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006e5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dca] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006e6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dcc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006e7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dce] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006e8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dd0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006e9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dd2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006ea] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dd4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006eb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dd6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006ec] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dd8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006ed] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dda] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006ee] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ddc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006ef] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dde] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006f0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00de0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006f1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00de2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006f2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00de4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006f3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00de6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006f4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00de8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006f5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dea] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006f6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dec] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006f7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dee] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006f8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00df0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006f9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00df2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006fa] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00df4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006fb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00df6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006fc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00df8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006fd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dfa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006fe] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dfc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006ff] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dfe] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00700] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e00] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00701] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e02] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00702] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e04] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00703] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e06] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00704] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e08] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00705] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e0a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00706] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e0c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00707] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e0e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00708] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e10] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00709] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e12] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0070a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e14] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0070b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e16] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0070c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e18] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0070d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e1a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0070e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e1c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0070f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e1e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00710] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e20] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00711] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e22] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00712] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e24] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00713] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e26] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00714] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e28] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00715] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e2a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00716] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e2c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00717] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e2e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00718] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e30] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00719] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e32] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0071a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e34] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0071b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e36] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0071c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e38] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0071d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e3a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0071e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e3c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0071f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e3e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00720] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e40] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00721] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e42] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00722] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e44] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00723] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e46] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00724] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e48] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00725] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e4a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00726] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e4c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00727] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e4e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00728] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e50] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00729] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e52] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0072a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e54] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0072b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e56] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0072c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e58] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0072d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e5a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0072e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e5c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0072f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e5e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00730] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e60] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00731] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e62] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00732] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e64] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00733] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e66] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00734] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e68] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00735] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e6a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00736] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e6c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00737] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e6e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00738] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e70] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00739] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e72] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0073a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e74] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0073b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e76] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0073c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e78] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0073d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e7a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0073e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e7c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0073f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e7e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00740] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e80] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00741] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e82] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00742] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e84] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00743] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e86] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00744] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e88] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00745] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e8a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00746] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e8c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00747] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e8e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00748] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e90] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00749] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e92] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0074a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e94] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0074b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e96] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0074c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e98] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0074d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e9a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0074e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e9c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0074f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e9e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00750] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ea0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00751] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ea2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00752] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ea4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00753] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ea6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00754] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ea8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00755] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eaa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00756] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eac] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00757] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eae] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00758] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eb0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00759] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eb2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0075a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eb4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0075b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eb6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0075c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eb8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0075d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eba] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0075e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ebc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0075f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ebe] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00760] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ec0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00761] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ec2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00762] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ec4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00763] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ec6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00764] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ec8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00765] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eca] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00766] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ecc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00767] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ece] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00768] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ed0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00769] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ed2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0076a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ed4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0076b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ed6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0076c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ed8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0076d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eda] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0076e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00edc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0076f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ede] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00770] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ee0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00771] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ee2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00772] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ee4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00773] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ee6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00774] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ee8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00775] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eea] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00776] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eec] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00777] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eee] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00778] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ef0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00779] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ef2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0077a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ef4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0077b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ef6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0077c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ef8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0077d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00efa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0077e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00efc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0077f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00efe] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00780] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f00] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00781] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f02] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00782] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f04] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00783] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f06] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00784] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f08] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00785] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f0a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00786] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f0c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00787] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f0e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00788] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f10] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00789] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f12] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0078a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f14] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0078b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f16] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0078c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f18] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0078d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f1a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0078e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f1c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0078f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f1e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00790] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f20] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00791] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f22] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00792] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f24] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00793] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f26] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00794] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f28] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00795] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f2a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00796] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f2c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00797] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f2e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00798] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f30] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00799] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f32] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0079a] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f34] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0079b] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f36] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0079c] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f38] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0079d] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f3a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0079e] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f3c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0079f] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f3e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007a0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f40] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007a1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f42] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007a2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f44] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007a3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f46] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007a4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f48] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007a5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f4a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007a6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f4c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007a7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f4e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007a8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f50] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007a9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f52] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007aa] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f54] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007ab] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f56] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007ac] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f58] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007ad] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f5a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007ae] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f5c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007af] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f5e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007b0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f60] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007b1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f62] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007b2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f64] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007b3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f66] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007b4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f68] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007b5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f6a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007b6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f6c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007b7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f6e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007b8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f70] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007b9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f72] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007ba] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f74] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007bb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f76] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007bc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f78] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007bd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f7a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007be] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f7c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007bf] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f7e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007c0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f80] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007c1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f82] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007c2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f84] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007c3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f86] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007c4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f88] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007c5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f8a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007c6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f8c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007c7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f8e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007c8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f90] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007c9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f92] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007ca] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f94] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007cb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f96] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007cc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f98] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007cd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f9a] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007ce] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f9c] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007cf] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f9e] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007d0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fa0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007d1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fa2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007d2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fa4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007d3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fa6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007d4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fa8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007d5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00faa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007d6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fac] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007d7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fae] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007d8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fb0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007d9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fb2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007da] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fb4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007db] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fb6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007dc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fb8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007dd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fba] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007de] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fbc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007df] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fbe] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007e0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fc0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007e1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fc2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007e2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fc4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007e3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fc6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007e4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fc8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007e5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fca] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007e6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fcc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007e7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fce] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007e8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fd0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007e9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fd2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007ea] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fd4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007eb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fd6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007ec] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fd8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007ed] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fda] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007ee] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fdc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007ef] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fde] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007f0] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fe0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007f1] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fe2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007f2] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fe4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007f3] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fe6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007f4] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fe8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007f5] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fea] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007f6] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fec] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007f7] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fee] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007f8] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ff0] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007f9] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ff2] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007fa] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ff4] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007fb] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ff6] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007fc] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ff8] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007fd] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ffa] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007fe] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ffc] ;
//end
//always_comb begin // 
               Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007ff] =  I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ffe] ;
//end
