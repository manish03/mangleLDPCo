 reg  ['h3ffff:0] [$clog2('h7000+1)-1:0] Ie48b0bc6f48b1df342b20ff8b41da9d9 ;
