//#;; Id7d2c4b2da7a6478426f10a28d9f9eba59a188d1bf2835798742825d32a11125 I8be3365cabaa6a0f90d2e64f03fa78268c135fe0b0758b576b447e9b2068d75d I18a0c098c7fb0098093fc0fd619c8032ae193215c5f695d7f5eaafa28aa64d70 I679eaac16659c013675081e715f7ef761bdd183f1d7f55d079eb46ad6e322ac5 I9ef2faffd23e7fdda264eeeb3114357fcb304142506cbb023c2894ac10f71654
/*Ic3f8d45b35548e4a4ee0b7181f1834df8a2e1aa0eea9b8c77323fcbf46bb42c8*/
////////////////////////////////////////////////////////////////////////////////
//# Copyright (c) 2018 Secantec
//# No Permission to modify and distribute this program
//# even if this copyright message remains unaltered.
//#
//# Author: Secantec 27 April, 2018
//# $Id: $//#
//# Revision History
//#       MM      17  April, 2018    Initial release
//#
////////////////////////////////////////////////////////////////////////////////

// /I51a1f05af85e342e3c849b47d387086476282d5f50dc240c19216d6edfb1eb5a/I58466ebdd352f801198118e294e38715f864985fd87977f348bfcd7db62e7c76 -I54e67ab9c29a6cfd19408098a96b2a40ede7e06aadcf77336da0dd2b57f25ba7 *I4395dc236d13a1c9b88a791fd2e1275bbb97b927d52e9b8c38248a0d57259aea* *Ic7c59e97212940ba254bbb99e5f908fec3434155e0fbb2f0a3f2ab5a6b4ba2a1* ; If0c929a9e723bc62724e30c7e396e576019dfcb8cfd0a3f264ee5d72e64e49d1 I04ad2bfad8cbdb3afbf9a26ea1454ac0a07c0eebc856992b38114cdcb5098c47.I3485639faf1591f3c16f295198e9389db5b33c949587ec48663597d4e00299d5 -If0c929a9e723bc62724e30c7e396e576019dfcb8cfd0a3f264ee5d72e64e49d1 I8803a3b234be60475d3d6498d388264bbc5edd49f43c780eee4753cddabfe052.1.sv > I8803a3b234be60475d3d6498d388264bbc5edd49f43c780eee4753cddabfe052.1.I04ad2bfad8cbdb3afbf9a26ea1454ac0a07c0eebc856992b38114cdcb5098c47.sv ; Ia8d1cfa1fc63160715eed9e8f5f39538f4520ff839d850162536352ec0a5509c -Ic572272153455b732903e10d0db7356fb56fb5d0a6a9064766547a1304406c33 -I8c2574892063f995fdf756bce07f46c1a5193e54cd52837ed91e32008ccf41ac -I4e1de0094e501762cba645b8d4663534d3eee7dc7d8bc675574f6b130d9f5302 I8803a3b234be60475d3d6498d388264bbc5edd49f43c780eee4753cddabfe052.1.I04ad2bfad8cbdb3afbf9a26ea1454ac0a07c0eebc856992b38114cdcb5098c47.sv -Iacac86c0e609ca906f632b0e2dacccb2b77d22b0621f20ebece1a4835b93f6f0 I8803a3b234be60475d3d6498d388264bbc5edd49f43c780eee4753cddabfe052.1.I04ad2bfad8cbdb3afbf9a26ea1454ac0a07c0eebc856992b38114cdcb5098c47.sv.I836ff184e7b41b1e13cb5fd89fa1de98dbbab99e9d2918913ff43b86a5c7c213

 /*Ic3f8d45b35548e4a4ee0b7181f1834df8a2e1aa0eea9b8c77323fcbf46bb42c8*/

/* I1e4d9aa7cb1ef438f80454b61c625f0c6aed19675cb2c2f865cbd2e2c3ef2ff7 Ib8a92ab2b5e2e68fc63a575fff1d62c25ec6d30209e164d82ec85f5576d9d940 I63985ce3eb57dbe35dec3a2e0dc38ffe14d2e2396edf773bd4f0298ce3ec7eff */

module  sntc_HamDist#(
// I168413ccee11e827c207105eecf061ecb7d6991383544364fda85556cdf96a57/I373a739f28b569ba97fa09dd5a21185f9bed4792859f1d9cc7fe4af7f6b9c7b7.sv
parameter MM   = 'h 000a8 ,
// parameter MM =  'h  000a8  , 
parameter NN   = 'h 000d0 ,
// parameter NN =  'h  000d0  , 
parameter cmax = 'h 00017 ,
// parameter cmax =  'h  00017  , 
parameter rmax = 'h 0000a ,
// parameter rmax =  'h  0000a  , 
// 208
// 168
parameter SUM_NN=$clog2(NN+1), // 8 : I47c35ffcd3135a74f03fef2155c1874927bc03c22812da0a352f40ca1d7339ea
parameter SUM_MM=$clog2(MM+1), // 8 : Ifa20411ae2befe271235475378a99513a77cfe0a9614b7cba4d2d92a1f1168c3
parameter LEN=MM,
//parameter SUM_LEN= SUM_MM
parameter SUM_LEN= 32
) (


input  wire [LEN-1:0]                         Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa,
input  wire [LEN-1:0]                         I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881,
output wire [SUM_LEN-1:0]                     sum_mm,

/* I1e4d9aa7cb1ef438f80454b61c625f0c6aed19675cb2c2f865cbd2e2c3ef2ff7 Ib8a92ab2b5e2e68fc63a575fff1d62c25ec6d30209e164d82ec85f5576d9d940 I5fedfe54fddcdc5145ac6dd38b4c3dead65f127535af2e07a7b9790515afdb04 */
input wire                                    clr,
/* I1e4d9aa7cb1ef438f80454b61c625f0c6aed19675cb2c2f865cbd2e2c3ef2ff7 I2f08a120cf6d1091827fd5d929bad0cbcaa5eff7ae0801098357ed0149cbc06e I5fedfe54fddcdc5145ac6dd38b4c3dead65f127535af2e07a7b9790515afdb04 */
input wire                                    rstn,
input wire                                    clk
);

`ifdef ENCRYPT
`endif

//  4 : Ifd0eae413952a156de9687eed7bb6378dedf004b3c5116c6a33c7ba5029d49a2

wire [SUM_LEN -1:0] I9015db1921f25e12204c6d0f9e52c76efabda6f8ad61870bd211efa68a974de0;
wire [SUM_LEN -1:0] Ie363a56342202df3680e91aea79f32ff8e2a62029212433aed75dce9fcc07bb4;
wire [SUM_LEN -1:0] Ic05031867d0c296a72de6ce5b1530277ba9d453fb21c2dcabad50817cac3baeb;
wire [SUM_LEN -1:0] I2f5c8c31c2c9a49215a291a3320e2951f741925115ce4f08d4e87641a9c6d286;
wire [SUM_LEN -1:0] I4e2fa42b4d9fc334936ac5b979d3d6098a764a79053bffc7051743cef60115c7;
wire [SUM_LEN -1:0] Ibcd479f48a16eb61d8e4bd6d59d735c5a1a54b123abf184b92bdb427b5f3f837;
wire [SUM_LEN -1:0] Idaca540dbf567c230af1c005a39b2fe1a058bea28b5dff26e45bc5bdb05f47e2;
wire [SUM_LEN -1:0] I88a90a0d707226b4fdd2b7c3425fa931d82cce4288bf4f9e15071c949eefcdc7;
wire [SUM_LEN -1:0] I7e1405f189f1c1a1d30ffe71069d6c718308281a467530c5d30b0730e96767d2;
wire [SUM_LEN -1:0] I9cc184be873d7a7a542eaa06c8c54877d964b05246097a857e50aec1d2d27e55;
wire [SUM_LEN -1:0] I119d576b67a1cd3cde6f756d53268817be990789873d05a8abaa97ce219170cc;
wire [SUM_LEN -1:0] I7d069d89dccfd691590505cc8ab2e7119be807e697e7a383434e79f0e561ee39;
wire [SUM_LEN -1:0] I96babb7e4864759d56a082de49b9ba922209a8b7f9c7d5c1f1ffacb69fd323cb;
wire [SUM_LEN -1:0] I472c8d1cd6c06f6b45c6a7e3eeea688c3ade09e0d2e65b47c7e0039f9ba3e2e8;
wire [SUM_LEN -1:0] I98120c2391baf4134cc30f567cdf58cebf0efb7336ea27358d040f4a9322d493;
wire [SUM_LEN -1:0] I872635255dfa96019499e3c343a1e00209328aa1a0786dee3184b4b2b4144f64;
wire [SUM_LEN -1:0] I144f6032be01c7c4715d215d24c3b26b3733a5c0561ae782105e9fe89e2e9be6;
wire [SUM_LEN -1:0] I0846a8903885db4cc60c2aaefb18ad455bcda9eca7b605ce4034b8137777fbae;
wire [SUM_LEN -1:0] I6b216f79c8be0cb8cf2ec3c5e25c118112a7d41eea659f34507a01b606d91e3a;
wire [SUM_LEN -1:0] I96ffec0fb72bb1de0b91ccab51b60c3b322c7311a3d6e80c4292539e95bf102a;
wire [SUM_LEN -1:0] I50b23de2cb7473fbb4f4097b53fc593e1a432b0d0b068703b13c1e4545d1254d;
wire [SUM_LEN -1:0] I2cdf3d868226af0127c35cb87aa18a5c79743a175363bd90b0229aeebbd904c9;
wire [SUM_LEN -1:0] I506eb86b96c16e51a96e7dffdc77922b117f2ad92e85ff1f0da0d1c35c1e9abf;
wire [SUM_LEN -1:0] I4750c0e01066ba7923ed9bba7eb616674d0160aeed7cf42042e2f7980f228682;

wire [LEN-1:0] Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e;
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00000] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00000] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00000];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00001] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00001] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00001];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00002] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00002] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00002];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00003] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00003] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00003];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00004] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00004] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00004];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00005] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00005] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00005];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00006] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00006] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00006];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00007] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00007] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00007];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00008] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00008] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00008];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00009] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00009] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00009];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00010] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00010] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00010];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00011] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00011] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00011];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00012] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00012] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00012];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00013] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00013] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00013];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00014] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00014] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00014];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00015] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00015] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00015];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00016] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00016] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00016];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00017] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00017] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00017];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00018] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00018] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00018];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00019] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00019] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00019];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00020] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00020] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00020];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00021] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00021] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00021];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00022] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00022] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00022];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00023] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00023] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00023];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00024] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00024] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00024];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00025] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00025] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00025];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00026] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00026] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00026];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00027] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00027] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00027];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00028] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00028] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00028];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00029] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00029] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00029];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00030] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00030] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00030];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00031] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00031] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00031];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00032] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00032] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00032];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00033] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00033] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00033];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00034] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00034] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00034];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00035] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00035] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00035];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00036] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00036] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00036];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00037] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00037] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00037];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00038] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00038] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00038];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00039] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00039] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00039];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00040] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00040] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00040];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00041] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00041] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00041];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00042] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00042] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00042];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00043] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00043] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00043];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00044] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00044] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00044];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00045] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00045] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00045];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00046] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00046] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00046];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00047] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00047] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00047];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00048] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00048] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00048];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00049] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00049] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00049];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00050] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00050] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00050];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00051] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00051] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00051];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00052] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00052] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00052];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00053] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00053] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00053];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00054] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00054] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00054];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00055] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00055] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00055];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00056] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00056] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00056];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00057] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00057] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00057];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00058] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00058] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00058];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00059] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00059] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00059];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00060] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00060] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00060];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00061] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00061] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00061];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00062] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00062] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00062];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00063] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00063] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00063];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00064] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00064] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00064];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00065] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00065] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00065];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00066] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00066] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00066];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00067] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00067] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00067];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00068] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00068] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00068];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00069] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00069] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00069];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00070] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00070] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00070];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00071] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00071] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00071];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00072] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00072] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00072];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00073] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00073] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00073];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00074] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00074] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00074];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00075] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00075] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00075];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00076] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00076] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00076];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00077] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00077] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00077];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00078] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00078] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00078];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00079] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00079] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00079];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00080] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00080] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00080];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00081] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00081] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00081];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00082] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00082] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00082];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00083] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00083] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00083];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00084] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00084] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00084];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00085] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00085] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00085];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00086] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00086] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00086];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00087] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00087] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00087];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00088] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00088] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00088];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00089] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00089] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00089];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00090] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00090] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00090];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00091] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00091] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00091];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00092] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00092] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00092];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00093] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00093] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00093];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00094] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00094] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00094];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00095] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00095] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00095];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00096] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00096] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00096];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00097] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00097] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00097];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00098] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00098] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00098];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00099] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00099] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00099];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00100] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00100] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00100];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00101] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00101] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00101];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00102] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00102] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00102];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00103] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00103] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00103];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00104] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00104] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00104];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00105] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00105] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00105];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00106] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00106] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00106];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00107] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00107] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00107];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00108] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00108] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00108];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00109] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00109] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00109];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00110] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00110] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00110];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00111] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00111] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00111];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00112] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00112] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00112];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00113] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00113] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00113];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00114] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00114] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00114];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00115] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00115] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00115];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00116] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00116] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00116];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00117] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00117] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00117];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00118] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00118] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00118];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00119] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00119] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00119];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00120] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00120] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00120];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00121] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00121] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00121];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00122] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00122] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00122];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00123] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00123] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00123];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00124] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00124] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00124];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00125] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00125] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00125];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00126] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00126] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00126];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00127] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00127] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00127];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00128] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00128] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00128];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00129] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00129] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00129];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00130] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00130] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00130];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00131] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00131] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00131];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00132] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00132] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00132];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00133] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00133] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00133];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00134] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00134] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00134];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00135] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00135] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00135];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00136] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00136] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00136];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00137] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00137] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00137];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00138] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00138] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00138];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00139] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00139] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00139];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00140] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00140] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00140];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00141] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00141] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00141];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00142] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00142] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00142];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00143] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00143] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00143];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00144] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00144] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00144];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00145] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00145] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00145];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00146] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00146] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00146];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00147] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00147] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00147];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00148] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00148] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00148];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00149] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00149] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00149];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00150] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00150] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00150];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00151] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00151] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00151];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00152] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00152] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00152];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00153] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00153] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00153];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00154] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00154] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00154];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00155] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00155] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00155];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00156] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00156] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00156];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00157] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00157] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00157];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00158] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00158] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00158];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00159] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00159] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00159];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00160] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00160] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00160];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00161] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00161] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00161];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00162] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00162] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00162];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00163] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00163] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00163];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00164] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00164] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00164];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00165] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00165] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00165];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00166] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00166] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00166];
assign       Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e['d 00167] = I2d711642b726b04401627ca9fbac32f5c8530fb1903cc4db02258717921a4881['d 00167] != Ia1fce4363854ff888cff4b8e7875d600c2682390412a8cf79b37d0b11148b0fa ['d 00167];


wire [3-1:0] I944779deeb85d7d8a0dba4d680192b22dbfb7a08a0577860a8d76104eaeb23a0;
            assign I944779deeb85d7d8a0dba4d680192b22dbfb7a08a0577860a8d76104eaeb23a0 =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[0] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[1] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[2] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[3] +
                                                0;
wire [3-1:0] I30ae112f8fb5e53f74e3988bc61fa8ea49accfe350f847a0ae85c922bd66aa3c;
            assign I30ae112f8fb5e53f74e3988bc61fa8ea49accfe350f847a0ae85c922bd66aa3c =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[4] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[5] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[6] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[7] +
                                                0;
wire [3-1:0] Ib0dcc7e27183fc209f5592897dda4d6e12e66396484354bf7ff51ab939d5a3dd;
            assign Ib0dcc7e27183fc209f5592897dda4d6e12e66396484354bf7ff51ab939d5a3dd =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[8] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[9] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[10] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[11] +
                                                0;
wire [3-1:0] I681e8f930bdf6be123094f5e6096415a9ee6b6d5615ba550505b413202be2e35;
            assign I681e8f930bdf6be123094f5e6096415a9ee6b6d5615ba550505b413202be2e35 =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[12] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[13] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[14] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[15] +
                                                0;
wire [3-1:0] I9b264334cf0f94f12d345114acfc1fcae739be55ce0050e4d9064477aa338002;
            assign I9b264334cf0f94f12d345114acfc1fcae739be55ce0050e4d9064477aa338002 =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[16] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[17] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[18] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[19] +
                                                0;
wire [3-1:0] If58eeaaf40ddd66bded568d044d3cbbcab3bf8f1d7bd52684093db555b679d53;
            assign If58eeaaf40ddd66bded568d044d3cbbcab3bf8f1d7bd52684093db555b679d53 =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[20] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[21] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[22] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[23] +
                                                0;
wire [3-1:0] I6f7e327d05991e592e81d9b7886844896adb5bc0d28a98830f1e3173c96b49ae;
            assign I6f7e327d05991e592e81d9b7886844896adb5bc0d28a98830f1e3173c96b49ae =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[24] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[25] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[26] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[27] +
                                                0;
wire [3-1:0] Iadc65eb532b959fb535efab73abbd460fc9ad3c6de17d9b767f41f23c97831e2;
            assign Iadc65eb532b959fb535efab73abbd460fc9ad3c6de17d9b767f41f23c97831e2 =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[28] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[29] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[30] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[31] +
                                                0;
wire [3-1:0] Idef1287e81d9b31855e0107e1f1fd5c155db49f96de751047ffde3ac6a8d303d;
            assign Idef1287e81d9b31855e0107e1f1fd5c155db49f96de751047ffde3ac6a8d303d =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[32] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[33] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[34] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[35] +
                                                0;
wire [3-1:0] I534b3818e2a9a99d41f89a2aa87b790cd94bb3deeac1eae7cbe0bffcc5886173;
            assign I534b3818e2a9a99d41f89a2aa87b790cd94bb3deeac1eae7cbe0bffcc5886173 =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[36] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[37] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[38] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[39] +
                                                0;
wire [3-1:0] I301afb5269dbacefd4c6a29e4e98eb3e8451091965013943d6892e582e25a18e;
            assign I301afb5269dbacefd4c6a29e4e98eb3e8451091965013943d6892e582e25a18e =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[40] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[41] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[42] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[43] +
                                                0;
wire [3-1:0] I8ffa56f768dd4ab0019c8b9b4b308eb832d2dfb97fe3b3f810fdc39dc509f03e;
            assign I8ffa56f768dd4ab0019c8b9b4b308eb832d2dfb97fe3b3f810fdc39dc509f03e =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[44] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[45] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[46] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[47] +
                                                0;
wire [3-1:0] Ibc8dac38b9f2fef1a593e9ea01a6b056909912b0d7fca6f4bd9a4a6a78ecedba;
            assign Ibc8dac38b9f2fef1a593e9ea01a6b056909912b0d7fca6f4bd9a4a6a78ecedba =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[48] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[49] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[50] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[51] +
                                                0;
wire [3-1:0] I98fe489c4ca3d321ad8fe7da1c9e91258367cde5794daab39249ba76744ec570;
            assign I98fe489c4ca3d321ad8fe7da1c9e91258367cde5794daab39249ba76744ec570 =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[52] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[53] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[54] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[55] +
                                                0;
wire [3-1:0] I379578f81074dcd51f23a8d4ba6cf0092993c26b8f0d4eea75dbd7f24c30aae1;
            assign I379578f81074dcd51f23a8d4ba6cf0092993c26b8f0d4eea75dbd7f24c30aae1 =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[56] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[57] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[58] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[59] +
                                                0;
wire [3-1:0] I03b75ee59fc3ad0aa7fea65d6a1f859e64560ea32bd430db518c94aea3242cf5;
            assign I03b75ee59fc3ad0aa7fea65d6a1f859e64560ea32bd430db518c94aea3242cf5 =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[60] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[61] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[62] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[63] +
                                                0;
wire [3-1:0] I3990d279646d68ef73d997cef6b27bd26a135e91cfebcc7a985fcb2f5cf954e0;
            assign I3990d279646d68ef73d997cef6b27bd26a135e91cfebcc7a985fcb2f5cf954e0 =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[64] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[65] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[66] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[67] +
                                                0;
wire [3-1:0] I40d29544ccebef7ebeebe1f36fc74248ea40136e22edbc2e02210ebdcb9adee6;
            assign I40d29544ccebef7ebeebe1f36fc74248ea40136e22edbc2e02210ebdcb9adee6 =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[68] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[69] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[70] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[71] +
                                                0;
wire [3-1:0] I27eca33c273a568e629e142f7aa368cc2bd0a123c2fbb420a160df42fc952f86;
            assign I27eca33c273a568e629e142f7aa368cc2bd0a123c2fbb420a160df42fc952f86 =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[72] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[73] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[74] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[75] +
                                                0;
wire [3-1:0] I4d0232bcffb0d85cc00f06ed58f90aaded6f73f678f05dcd8693a466bce94934;
            assign I4d0232bcffb0d85cc00f06ed58f90aaded6f73f678f05dcd8693a466bce94934 =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[76] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[77] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[78] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[79] +
                                                0;
wire [3-1:0] Ic23eb7e5f040413bf0572a87b07c11af5fba085089794d3bf84857a4490ff2f8;
            assign Ic23eb7e5f040413bf0572a87b07c11af5fba085089794d3bf84857a4490ff2f8 =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[80] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[81] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[82] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[83] +
                                                0;
wire [3-1:0] I6f2e83d126bcd76ea0eb4a4c7b90c4be34d25f8b809ff2c4a6c54c1749a05593;
            assign I6f2e83d126bcd76ea0eb4a4c7b90c4be34d25f8b809ff2c4a6c54c1749a05593 =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[84] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[85] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[86] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[87] +
                                                0;
wire [3-1:0] Ic33d190da2d5120cc4b7ee4c677d091adafdecc9f0f54b1ceaf3c9e22a0f204a;
            assign Ic33d190da2d5120cc4b7ee4c677d091adafdecc9f0f54b1ceaf3c9e22a0f204a =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[88] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[89] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[90] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[91] +
                                                0;
wire [3-1:0] Icfa3d5a05dfa45e86474c759aa04152445c0272f3cafae493aac36ccc848bfb6;
            assign Icfa3d5a05dfa45e86474c759aa04152445c0272f3cafae493aac36ccc848bfb6 =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[92] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[93] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[94] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[95] +
                                                0;
wire [3-1:0] Ia33b424c118f84dd02fc1130a0e577da602883af6988e0402a5342b8e2c1ff57;
            assign Ia33b424c118f84dd02fc1130a0e577da602883af6988e0402a5342b8e2c1ff57 =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[96] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[97] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[98] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[99] +
                                                0;
wire [3-1:0] I9afe770a10eb445d0644c69016263771e6709cd38e816997b92ff31376d7ecdf;
            assign I9afe770a10eb445d0644c69016263771e6709cd38e816997b92ff31376d7ecdf =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[100] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[101] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[102] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[103] +
                                                0;
wire [3-1:0] Idc27cacedbaa5fea4028024f3e7a02548000ed9c77731acb65f5f87727d6b13d;
            assign Idc27cacedbaa5fea4028024f3e7a02548000ed9c77731acb65f5f87727d6b13d =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[104] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[105] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[106] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[107] +
                                                0;
wire [3-1:0] Ida5f4ac896d3fefa909bc7714d17c74e645262d648c58a0e32a5687e1122c37b;
            assign Ida5f4ac896d3fefa909bc7714d17c74e645262d648c58a0e32a5687e1122c37b =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[108] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[109] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[110] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[111] +
                                                0;
wire [3-1:0] Iaed16423a55746841a2541db0f40cdfc54c2616e30a6363f48da4af6c5d3d581;
            assign Iaed16423a55746841a2541db0f40cdfc54c2616e30a6363f48da4af6c5d3d581 =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[112] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[113] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[114] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[115] +
                                                0;
wire [3-1:0] I92bb1c56abdd696f780757ba21c0bcd62ad5957ad3214e0230b0a2ffa91d0591;
            assign I92bb1c56abdd696f780757ba21c0bcd62ad5957ad3214e0230b0a2ffa91d0591 =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[116] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[117] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[118] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[119] +
                                                0;
wire [3-1:0] If98975980e19197790888665ab6d1cabbf2cb08fb50dbb3e7abc103e729a8e3e;
            assign If98975980e19197790888665ab6d1cabbf2cb08fb50dbb3e7abc103e729a8e3e =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[120] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[121] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[122] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[123] +
                                                0;
wire [3-1:0] Icf5371b8dce23de626277fef7c0621d3abfdf509a0c5caedb7185fb8de66de6c;
            assign Icf5371b8dce23de626277fef7c0621d3abfdf509a0c5caedb7185fb8de66de6c =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[124] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[125] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[126] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[127] +
                                                0;
wire [3-1:0] I4b9052836925b80d7cd73d27dfea63d073ef22925e4c08af155054d2615059d4;
            assign I4b9052836925b80d7cd73d27dfea63d073ef22925e4c08af155054d2615059d4 =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[128] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[129] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[130] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[131] +
                                                0;
wire [3-1:0] I7213b5da067a4cf0fa9dbbcb9a243d8c087a46e5e5e1ed591a476ce5deb3a3be;
            assign I7213b5da067a4cf0fa9dbbcb9a243d8c087a46e5e5e1ed591a476ce5deb3a3be =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[132] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[133] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[134] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[135] +
                                                0;
wire [3-1:0] I00a71d54b5f9cd5d79695a089753efce7c73de17456f397d5a50031e3e53f8ed;
            assign I00a71d54b5f9cd5d79695a089753efce7c73de17456f397d5a50031e3e53f8ed =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[136] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[137] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[138] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[139] +
                                                0;
wire [3-1:0] I99a81679d66bdb8271d2c90dc227a8d7815feaf562bc2882f95a767959a476f0;
            assign I99a81679d66bdb8271d2c90dc227a8d7815feaf562bc2882f95a767959a476f0 =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[140] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[141] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[142] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[143] +
                                                0;
wire [3-1:0] I99cf8aa9f971165076a33d633cab8a3677c745ea863ebef88c100240e68375c5;
            assign I99cf8aa9f971165076a33d633cab8a3677c745ea863ebef88c100240e68375c5 =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[144] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[145] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[146] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[147] +
                                                0;
wire [3-1:0] I71c92468bead01c807e245fcfffa56a323af641d656d3cf3f4021d9b48371cdd;
            assign I71c92468bead01c807e245fcfffa56a323af641d656d3cf3f4021d9b48371cdd =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[148] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[149] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[150] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[151] +
                                                0;
wire [3-1:0] I231fbdd5cdcd478b0599b9c2b024f989e68738c9ecf89dc0344261e7e1f7420e;
            assign I231fbdd5cdcd478b0599b9c2b024f989e68738c9ecf89dc0344261e7e1f7420e =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[152] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[153] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[154] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[155] +
                                                0;
wire [3-1:0] If7265544cf5d4d7e524a99fbc445bf2ce46aaa08fcff9c101d7003b83ae84aa6;
            assign If7265544cf5d4d7e524a99fbc445bf2ce46aaa08fcff9c101d7003b83ae84aa6 =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[156] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[157] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[158] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[159] +
                                                0;
wire [3-1:0] I28f49a0531b318ea6e3567665b90bf09c7e5c8974ef250e20f4dbfd8d17cb50b;
            assign I28f49a0531b318ea6e3567665b90bf09c7e5c8974ef250e20f4dbfd8d17cb50b =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[160] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[161] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[162] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[163] +
                                                0;
wire [3-1:0] I472015fa50db0b97d7634fc9d1c8a86b2ae61b5afcc6e655e57640b36123b256;
            assign I472015fa50db0b97d7634fc9d1c8a86b2ae61b5afcc6e655e57640b36123b256 =
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[164] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[165] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[166] +
                                                     Ic614281386cda8887a253dfbc2a7e2ea3029cc9dbd74450caeb2661feaab6e8e[167] +
                                                0;

// 42 : LEN
wire [5-1:0] Id872257e09ad72adae3049b08be33b2cc608120b23fd969f76d811478b5a969e;
                              assign Id872257e09ad72adae3049b08be33b2cc608120b23fd969f76d811478b5a969e =
                                                     I944779deeb85d7d8a0dba4d680192b22dbfb7a08a0577860a8d76104eaeb23a0 +
                                                     I30ae112f8fb5e53f74e3988bc61fa8ea49accfe350f847a0ae85c922bd66aa3c +
                                                     Ib0dcc7e27183fc209f5592897dda4d6e12e66396484354bf7ff51ab939d5a3dd +
                                                     I681e8f930bdf6be123094f5e6096415a9ee6b6d5615ba550505b413202be2e35 ;
wire [5-1:0] Id5f810559af335642435a2fd85f43f38c0b6c2d438b880fb1e5a2b5aa1cba29d;
                              assign Id5f810559af335642435a2fd85f43f38c0b6c2d438b880fb1e5a2b5aa1cba29d =
                                                     I9b264334cf0f94f12d345114acfc1fcae739be55ce0050e4d9064477aa338002 +
                                                     If58eeaaf40ddd66bded568d044d3cbbcab3bf8f1d7bd52684093db555b679d53 +
                                                     I6f7e327d05991e592e81d9b7886844896adb5bc0d28a98830f1e3173c96b49ae +
                                                     Iadc65eb532b959fb535efab73abbd460fc9ad3c6de17d9b767f41f23c97831e2 ;
wire [5-1:0] Ia4cbc49fa8bcd6f8d1c8f963b8b6c208a97811cc3fee7a5888f552b31762c3ae;
                              assign Ia4cbc49fa8bcd6f8d1c8f963b8b6c208a97811cc3fee7a5888f552b31762c3ae =
                                                     Idef1287e81d9b31855e0107e1f1fd5c155db49f96de751047ffde3ac6a8d303d +
                                                     I534b3818e2a9a99d41f89a2aa87b790cd94bb3deeac1eae7cbe0bffcc5886173 +
                                                     I301afb5269dbacefd4c6a29e4e98eb3e8451091965013943d6892e582e25a18e +
                                                     I8ffa56f768dd4ab0019c8b9b4b308eb832d2dfb97fe3b3f810fdc39dc509f03e ;
wire [5-1:0] Ib4f35d051c3f92b956d064e7022e3ca504a6f6834cc8f08aac8ee98b84627e79;
                              assign Ib4f35d051c3f92b956d064e7022e3ca504a6f6834cc8f08aac8ee98b84627e79 =
                                                     Ibc8dac38b9f2fef1a593e9ea01a6b056909912b0d7fca6f4bd9a4a6a78ecedba +
                                                     I98fe489c4ca3d321ad8fe7da1c9e91258367cde5794daab39249ba76744ec570 +
                                                     I379578f81074dcd51f23a8d4ba6cf0092993c26b8f0d4eea75dbd7f24c30aae1 +
                                                     I03b75ee59fc3ad0aa7fea65d6a1f859e64560ea32bd430db518c94aea3242cf5 ;
wire [5-1:0] I5b2d9adcfd821b7f95d25f10c5e3cee9b2477c0e8c49fc8e56cc36dc2d503de7;
                              assign I5b2d9adcfd821b7f95d25f10c5e3cee9b2477c0e8c49fc8e56cc36dc2d503de7 =
                                                     I3990d279646d68ef73d997cef6b27bd26a135e91cfebcc7a985fcb2f5cf954e0 +
                                                     I40d29544ccebef7ebeebe1f36fc74248ea40136e22edbc2e02210ebdcb9adee6 +
                                                     I27eca33c273a568e629e142f7aa368cc2bd0a123c2fbb420a160df42fc952f86 +
                                                     I4d0232bcffb0d85cc00f06ed58f90aaded6f73f678f05dcd8693a466bce94934 ;
wire [5-1:0] I761b25fd3957bda2e126a3c7be9803247eee75a759a51e2dc1c014020439c90b;
                              assign I761b25fd3957bda2e126a3c7be9803247eee75a759a51e2dc1c014020439c90b =
                                                     Ic23eb7e5f040413bf0572a87b07c11af5fba085089794d3bf84857a4490ff2f8 +
                                                     I6f2e83d126bcd76ea0eb4a4c7b90c4be34d25f8b809ff2c4a6c54c1749a05593 +
                                                     Ic33d190da2d5120cc4b7ee4c677d091adafdecc9f0f54b1ceaf3c9e22a0f204a +
                                                     Icfa3d5a05dfa45e86474c759aa04152445c0272f3cafae493aac36ccc848bfb6 ;
wire [5-1:0] I632b16934db0ca8390bf04f37a882a6a199e4bffea5f5ef3cd4b29b27fabe8a9;
                              assign I632b16934db0ca8390bf04f37a882a6a199e4bffea5f5ef3cd4b29b27fabe8a9 =
                                                     Ia33b424c118f84dd02fc1130a0e577da602883af6988e0402a5342b8e2c1ff57 +
                                                     I9afe770a10eb445d0644c69016263771e6709cd38e816997b92ff31376d7ecdf +
                                                     Idc27cacedbaa5fea4028024f3e7a02548000ed9c77731acb65f5f87727d6b13d +
                                                     Ida5f4ac896d3fefa909bc7714d17c74e645262d648c58a0e32a5687e1122c37b ;
wire [5-1:0] Ica0df511966bf0e4843f0ec06a57111d918af0db048b8c20d90f7c625e269667;
                              assign Ica0df511966bf0e4843f0ec06a57111d918af0db048b8c20d90f7c625e269667 =
                                                     Iaed16423a55746841a2541db0f40cdfc54c2616e30a6363f48da4af6c5d3d581 +
                                                     I92bb1c56abdd696f780757ba21c0bcd62ad5957ad3214e0230b0a2ffa91d0591 +
                                                     If98975980e19197790888665ab6d1cabbf2cb08fb50dbb3e7abc103e729a8e3e +
                                                     Icf5371b8dce23de626277fef7c0621d3abfdf509a0c5caedb7185fb8de66de6c ;
wire [5-1:0] I220b6e7689b6773fe7147e42a9a952d6746995a7a93b8bcb08bee07853258dac;
                              assign I220b6e7689b6773fe7147e42a9a952d6746995a7a93b8bcb08bee07853258dac =
                                                     I4b9052836925b80d7cd73d27dfea63d073ef22925e4c08af155054d2615059d4 +
                                                     I7213b5da067a4cf0fa9dbbcb9a243d8c087a46e5e5e1ed591a476ce5deb3a3be +
                                                     I00a71d54b5f9cd5d79695a089753efce7c73de17456f397d5a50031e3e53f8ed +
                                                     I99a81679d66bdb8271d2c90dc227a8d7815feaf562bc2882f95a767959a476f0 ;
wire [5-1:0] I933fb93f939f4930a0b36a15a438d2fcbaa31c7a715c22dea89729331a6feb02;
                              assign I933fb93f939f4930a0b36a15a438d2fcbaa31c7a715c22dea89729331a6feb02 =
                                                     I99cf8aa9f971165076a33d633cab8a3677c745ea863ebef88c100240e68375c5 +
                                                     I71c92468bead01c807e245fcfffa56a323af641d656d3cf3f4021d9b48371cdd +
                                                     I231fbdd5cdcd478b0599b9c2b024f989e68738c9ecf89dc0344261e7e1f7420e +
                                                     If7265544cf5d4d7e524a99fbc445bf2ce46aaa08fcff9c101d7003b83ae84aa6 ;
wire [5-1:0] I7cde0d224f7434d846208a3e66c9bfff5a857203bd4c67a203bab91e7fd144b9;
                              assign I7cde0d224f7434d846208a3e66c9bfff5a857203bd4c67a203bab91e7fd144b9 =
                                                     I28f49a0531b318ea6e3567665b90bf09c7e5c8974ef250e20f4dbfd8d17cb50b +
                                                     I472015fa50db0b97d7634fc9d1c8a86b2ae61b5afcc6e655e57640b36123b256 ;
// 11 : LEN
wire [7-1:0] I17850decf33052d6ee448d09a79ba5ec643b93cda252a7c1b69b8426051964c7;
                              assign I17850decf33052d6ee448d09a79ba5ec643b93cda252a7c1b69b8426051964c7 =
                                                     Id872257e09ad72adae3049b08be33b2cc608120b23fd969f76d811478b5a969e +
                                                     Id5f810559af335642435a2fd85f43f38c0b6c2d438b880fb1e5a2b5aa1cba29d +
                                                     Ia4cbc49fa8bcd6f8d1c8f963b8b6c208a97811cc3fee7a5888f552b31762c3ae +
                                                     Ib4f35d051c3f92b956d064e7022e3ca504a6f6834cc8f08aac8ee98b84627e79 ;
wire [7-1:0] Ie11385a61ce8515a354afedae70f4030bfb1f8a8064c7a537caae2669a79db18;
                              assign Ie11385a61ce8515a354afedae70f4030bfb1f8a8064c7a537caae2669a79db18 =
                                                     I5b2d9adcfd821b7f95d25f10c5e3cee9b2477c0e8c49fc8e56cc36dc2d503de7 +
                                                     I761b25fd3957bda2e126a3c7be9803247eee75a759a51e2dc1c014020439c90b +
                                                     I632b16934db0ca8390bf04f37a882a6a199e4bffea5f5ef3cd4b29b27fabe8a9 +
                                                     Ica0df511966bf0e4843f0ec06a57111d918af0db048b8c20d90f7c625e269667 ;
wire [7-1:0] I0eaf99572db3b5e62bc183d9eb559fc01e158b08f6bdeb776d92ae0d7688d44d;
                              assign I0eaf99572db3b5e62bc183d9eb559fc01e158b08f6bdeb776d92ae0d7688d44d =
                                                     I220b6e7689b6773fe7147e42a9a952d6746995a7a93b8bcb08bee07853258dac +
                                                     I933fb93f939f4930a0b36a15a438d2fcbaa31c7a715c22dea89729331a6feb02 +
                                                     I7cde0d224f7434d846208a3e66c9bfff5a857203bd4c67a203bab91e7fd144b9 ;
// 3 : LEN
wire [9-1:0] I10d6ebc64d85d0e02df2ff807063c1da6668a6b4eabc82186ca190fdfb864e4f;
                              assign I10d6ebc64d85d0e02df2ff807063c1da6668a6b4eabc82186ca190fdfb864e4f =
                                                     I17850decf33052d6ee448d09a79ba5ec643b93cda252a7c1b69b8426051964c7 +
                                                     Ie11385a61ce8515a354afedae70f4030bfb1f8a8064c7a537caae2669a79db18 +
                                                     I0eaf99572db3b5e62bc183d9eb559fc01e158b08f6bdeb776d92ae0d7688d44d ;
assign sum_mm = I10d6ebc64d85d0e02df2ff807063c1da6668a6b4eabc82186ca190fdfb864e4f;


`ifdef ENCRYPT
`endif

endmodule

