//`include "GF2_LDPC_flogtanh_0x00004_assign_inc.sv"
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00000] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00000] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00001] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00001] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00002] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00003] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00002] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00004] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00005] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00003] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00006] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00007] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00004] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00008] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00009] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00005] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0000a] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0000b] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00006] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0000c] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0000d] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00007] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0000e] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0000f] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00008] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00010] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00011] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00009] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00012] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00013] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0000a] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00014] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00015] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0000b] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00016] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00017] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0000c] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00018] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00019] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0000d] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0001a] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0001b] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0000e] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0001c] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0001d] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0000f] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0001e] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0001f] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00010] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00020] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00021] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00011] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00022] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00023] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00012] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00024] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00025] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00013] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00026] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00027] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00014] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00028] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00029] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00015] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0002a] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0002b] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00016] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0002c] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0002d] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00017] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0002e] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0002f] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00018] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00030] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00031] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00019] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00032] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00033] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0001a] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00034] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00035] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0001b] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00036] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00037] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0001c] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00038] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00039] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0001d] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0003a] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0003b] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0001e] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0003c] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0003d] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0001f] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0003e] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0003f] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00020] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00040] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00041] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00021] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00042] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00043] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00022] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00044] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00045] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00023] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00046] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00047] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00024] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00048] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00049] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00025] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0004a] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0004b] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00026] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0004c] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0004d] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00027] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0004e] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0004f] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00028] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00050] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00051] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00029] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00052] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00053] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0002a] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00054] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00055] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0002b] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00056] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00057] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0002c] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00058] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00059] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0002d] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0005a] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0005b] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0002e] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0005c] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0005d] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0002f] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0005e] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0005f] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00030] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00060] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00061] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00031] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00062] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00063] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00032] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00064] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00065] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00033] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00066] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00067] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00034] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00068] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00069] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00035] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0006a] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0006b] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00036] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0006c] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0006d] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00037] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0006e] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0006f] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00038] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00070] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00071] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00039] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00072] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00073] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0003a] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00074] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00075] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0003b] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00076] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00077] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0003c] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00078] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00079] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0003d] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0007a] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0007b] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0003e] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0007c] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0007d] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0003f] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0007e] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0007f] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00040] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00080] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00081] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00041] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00082] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00083] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00042] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00084] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00085] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00043] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00086] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00087] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00044] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00088] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00089] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00045] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0008a] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0008b] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00046] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0008c] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0008d] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00047] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0008e] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0008f] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00048] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00090] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00091] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00049] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00092] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00093] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0004a] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00094] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00095] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0004b] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00096] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00097] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0004c] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00098] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00099] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0004d] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0009a] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0009b] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0004e] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0009c] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0009d] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0004f] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0009e] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0009f] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00050] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000a0] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000a1] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00051] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000a2] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000a3] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00052] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000a4] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000a5] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00053] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000a6] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000a7] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00054] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000a8] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000a9] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00055] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000aa] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000ab] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00056] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000ac] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000ad] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00057] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000ae] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000af] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00058] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000b0] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000b1] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00059] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000b2] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000b3] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0005a] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000b4] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000b5] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0005b] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000b6] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000b7] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0005c] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000b8] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000b9] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0005d] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000ba] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000bb] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0005e] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000bc] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000bd] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0005f] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000be] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000bf] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00060] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000c0] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000c1] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00061] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000c2] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000c3] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00062] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000c4] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000c5] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00063] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000c6] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000c7] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00064] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000c8] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000c9] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00065] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000ca] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000cb] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00066] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000cc] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000cd] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00067] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000ce] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000cf] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00068] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000d0] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000d1] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00069] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000d2] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000d3] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0006a] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000d4] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000d5] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0006b] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000d6] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000d7] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0006c] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000d8] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000d9] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0006d] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000da] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000db] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0006e] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000dc] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000dd] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0006f] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000de] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000df] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00070] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000e0] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000e1] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00071] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000e2] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000e3] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00072] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000e4] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000e5] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00073] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000e6] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000e7] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00074] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000e8] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000e9] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00075] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000ea] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000eb] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00076] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000ec] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000ed] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00077] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000ee] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000ef] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00078] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000f0] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000f1] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00079] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000f2] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000f3] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0007a] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000f4] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000f5] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0007b] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000f6] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000f7] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0007c] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000f8] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000f9] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0007d] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000fa] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000fb] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0007e] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000fc] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000fd] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0007f] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h000fe] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h000ff] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00080] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00100] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00101] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00081] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00102] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00103] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00082] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00104] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00105] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00083] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00106] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00107] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00084] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00108] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00109] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00085] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0010a] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0010b] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00086] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0010c] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0010d] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00087] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0010e] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0010f] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00088] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00110] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00111] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00089] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00112] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00113] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0008a] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00114] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00115] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0008b] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00116] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00117] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0008c] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00118] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00119] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0008d] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0011a] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0011b] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0008e] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0011c] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0011d] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0008f] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0011e] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0011f] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00090] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00120] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00121] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00091] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00122] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00123] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00092] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00124] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00125] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00093] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00126] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00127] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00094] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00128] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00129] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00095] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0012a] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0012b] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00096] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0012c] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0012d] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00097] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0012e] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0012f] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00098] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00130] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00131] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00099] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00132] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00133] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0009a] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00134] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00135] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0009b] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00136] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00137] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0009c] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00138] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00139] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0009d] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0013a] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0013b] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0009e] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0013c] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0013d] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0009f] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0013e] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0013f] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000a0] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00140] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00141] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000a1] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00142] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00143] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000a2] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00144] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00145] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000a3] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00146] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00147] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000a4] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00148] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00149] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000a5] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0014a] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0014b] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000a6] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0014c] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0014d] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000a7] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0014e] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0014f] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000a8] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00150] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00151] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000a9] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00152] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00153] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000aa] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00154] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00155] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000ab] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00156] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00157] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000ac] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00158] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00159] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000ad] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0015a] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0015b] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000ae] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0015c] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0015d] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000af] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0015e] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0015f] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000b0] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00160] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00161] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000b1] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00162] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00163] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000b2] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00164] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00165] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000b3] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00166] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00167] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000b4] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00168] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00169] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000b5] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0016a] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0016b] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000b6] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0016c] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0016d] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000b7] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0016e] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0016f] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000b8] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00170] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00171] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000b9] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00172] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00173] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000ba] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00174] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00175] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000bb] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00176] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00177] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000bc] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00178] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00179] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000bd] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0017a] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0017b] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000be] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0017c] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0017d] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000bf] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0017e] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0017f] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000c0] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00180] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00181] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000c1] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00182] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00183] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000c2] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00184] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00185] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000c3] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00186] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00187] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000c4] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00188] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00189] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000c5] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0018a] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0018b] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000c6] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0018c] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0018d] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000c7] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0018e] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0018f] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000c8] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00190] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00191] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000c9] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00192] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00193] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000ca] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00194] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00195] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000cb] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00196] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00197] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000cc] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00198] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00199] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000cd] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0019a] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0019b] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000ce] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0019c] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0019d] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000cf] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0019e] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0019f] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000d0] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001a0] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001a1] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000d1] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001a2] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001a3] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000d2] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001a4] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001a5] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000d3] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001a6] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001a7] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000d4] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001a8] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001a9] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000d5] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001aa] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001ab] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000d6] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001ac] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001ad] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000d7] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001ae] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001af] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000d8] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001b0] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001b1] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000d9] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001b2] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001b3] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000da] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001b4] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001b5] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000db] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001b6] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001b7] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000dc] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001b8] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001b9] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000dd] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001ba] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001bb] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000de] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001bc] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001bd] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000df] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001be] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001bf] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000e0] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001c0] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001c1] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000e1] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001c2] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001c3] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000e2] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001c4] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001c5] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000e3] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001c6] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001c7] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000e4] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001c8] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001c9] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000e5] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001ca] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001cb] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000e6] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001cc] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001cd] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000e7] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001ce] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001cf] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000e8] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001d0] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001d1] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000e9] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001d2] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001d3] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000ea] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001d4] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001d5] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000eb] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001d6] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001d7] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000ec] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001d8] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001d9] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000ed] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001da] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001db] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000ee] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001dc] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001dd] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000ef] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001de] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001df] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000f0] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001e0] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001e1] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000f1] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001e2] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001e3] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000f2] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001e4] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001e5] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000f3] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001e6] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001e7] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000f4] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001e8] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001e9] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000f5] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001ea] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001eb] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000f6] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001ec] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001ed] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000f7] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001ee] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001ef] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000f8] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001f0] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001f1] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000f9] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001f2] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001f3] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000fa] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001f4] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001f5] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000fb] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001f6] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001f7] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000fc] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001f8] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001f9] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000fd] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001fa] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001fb] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000fe] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001fc] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001fd] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h000ff] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h001fe] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h001ff] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00100] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00200] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00201] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00101] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00202] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00203] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00102] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00204] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00205] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00103] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00206] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00207] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00104] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00208] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00209] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00105] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0020a] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0020b] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00106] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0020c] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0020d] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00107] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0020e] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0020f] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00108] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00210] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00211] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00109] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00212] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00213] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0010a] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00214] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00215] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0010b] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00216] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00217] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0010c] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00218] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00219] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0010d] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0021a] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0021b] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0010e] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0021c] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0021d] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0010f] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0021e] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0021f] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00110] =  I8a0037ad2845a3fbba9da380a8b8a576['h00220] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00111] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00222] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00223] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00112] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00224] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00225] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00113] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00226] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00227] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00114] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00228] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00229] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00115] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0022a] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0022b] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00116] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0022c] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0022d] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00117] =  I8a0037ad2845a3fbba9da380a8b8a576['h0022e] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00118] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00230] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00231] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00119] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00232] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00233] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0011a] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00234] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00235] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0011b] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00236] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00237] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0011c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00238] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0011d] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0023a] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0023b] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0011e] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0023c] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0023d] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0011f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0023e] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00120] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00240] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00241] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00121] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00242] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00243] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00122] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00244] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00245] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00123] =  I8a0037ad2845a3fbba9da380a8b8a576['h00246] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00124] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00248] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00249] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00125] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0024a] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0024b] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00126] =  I8a0037ad2845a3fbba9da380a8b8a576['h0024c] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00127] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0024e] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0024f] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00128] =  I8a0037ad2845a3fbba9da380a8b8a576['h00250] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00129] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00252] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00253] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0012a] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00254] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00255] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0012b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00256] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0012c] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00258] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00259] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0012d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0025a] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0012e] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0025c] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0025d] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0012f] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0025e] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0025f] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00130] =  I8a0037ad2845a3fbba9da380a8b8a576['h00260] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00131] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00262] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00263] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00132] =  I8a0037ad2845a3fbba9da380a8b8a576['h00264] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00133] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00266] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00267] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00134] =  I8a0037ad2845a3fbba9da380a8b8a576['h00268] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00135] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0026a] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0026b] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00136] =  I8a0037ad2845a3fbba9da380a8b8a576['h0026c] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00137] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0026e] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0026f] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00138] =  I8a0037ad2845a3fbba9da380a8b8a576['h00270] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00139] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00272] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00273] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0013a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00274] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0013b] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00276] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00277] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0013c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00278] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0013d] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0027a] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0027b] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0013e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0027c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0013f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0027e] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00140] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00280] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00281] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00141] =  I8a0037ad2845a3fbba9da380a8b8a576['h00282] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00142] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00284] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00285] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00143] =  I8a0037ad2845a3fbba9da380a8b8a576['h00286] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00144] =  I8a0037ad2845a3fbba9da380a8b8a576['h00288] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00145] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0028a] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0028b] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00146] =  I8a0037ad2845a3fbba9da380a8b8a576['h0028c] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00147] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0028e] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0028f] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00148] =  I8a0037ad2845a3fbba9da380a8b8a576['h00290] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00149] =  I8a0037ad2845a3fbba9da380a8b8a576['h00292] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0014a] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00294] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00295] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0014b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00296] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0014c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00298] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0014d] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0029a] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0029b] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0014e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0029c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0014f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0029e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00150] =  I8a0037ad2845a3fbba9da380a8b8a576['h002a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00151] =  I8a0037ad2845a3fbba9da380a8b8a576['h002a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00152] =  I8a0037ad2845a3fbba9da380a8b8a576['h002a4] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00153] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h002a6] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h002a7] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00154] =  I8a0037ad2845a3fbba9da380a8b8a576['h002a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00155] =  I8a0037ad2845a3fbba9da380a8b8a576['h002aa] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00156] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h002ac] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h002ad] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00157] =  I8a0037ad2845a3fbba9da380a8b8a576['h002ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00158] =  I8a0037ad2845a3fbba9da380a8b8a576['h002b0] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00159] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h002b2] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h002b3] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0015a] =  I8a0037ad2845a3fbba9da380a8b8a576['h002b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0015b] =  I8a0037ad2845a3fbba9da380a8b8a576['h002b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0015c] =  I8a0037ad2845a3fbba9da380a8b8a576['h002b8] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0015d] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h002ba] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h002bb] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0015e] =  I8a0037ad2845a3fbba9da380a8b8a576['h002bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0015f] =  I8a0037ad2845a3fbba9da380a8b8a576['h002be] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00160] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h002c0] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h002c1] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00161] =  I8a0037ad2845a3fbba9da380a8b8a576['h002c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00162] =  I8a0037ad2845a3fbba9da380a8b8a576['h002c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00163] =  I8a0037ad2845a3fbba9da380a8b8a576['h002c6] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00164] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h002c8] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h002c9] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00165] =  I8a0037ad2845a3fbba9da380a8b8a576['h002ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00166] =  I8a0037ad2845a3fbba9da380a8b8a576['h002cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00167] =  I8a0037ad2845a3fbba9da380a8b8a576['h002ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00168] =  I8a0037ad2845a3fbba9da380a8b8a576['h002d0] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00169] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h002d2] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h002d3] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0016a] =  I8a0037ad2845a3fbba9da380a8b8a576['h002d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0016b] =  I8a0037ad2845a3fbba9da380a8b8a576['h002d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0016c] =  I8a0037ad2845a3fbba9da380a8b8a576['h002d8] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0016d] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h002da] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h002db] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0016e] =  I8a0037ad2845a3fbba9da380a8b8a576['h002dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0016f] =  I8a0037ad2845a3fbba9da380a8b8a576['h002de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00170] =  I8a0037ad2845a3fbba9da380a8b8a576['h002e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00171] =  I8a0037ad2845a3fbba9da380a8b8a576['h002e2] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00172] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h002e4] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h002e5] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00173] =  I8a0037ad2845a3fbba9da380a8b8a576['h002e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00174] =  I8a0037ad2845a3fbba9da380a8b8a576['h002e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00175] =  I8a0037ad2845a3fbba9da380a8b8a576['h002ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00176] =  I8a0037ad2845a3fbba9da380a8b8a576['h002ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00177] =  I8a0037ad2845a3fbba9da380a8b8a576['h002ee] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00178] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h002f0] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h002f1] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00179] =  I8a0037ad2845a3fbba9da380a8b8a576['h002f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0017a] =  I8a0037ad2845a3fbba9da380a8b8a576['h002f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0017b] =  I8a0037ad2845a3fbba9da380a8b8a576['h002f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0017c] =  I8a0037ad2845a3fbba9da380a8b8a576['h002f8] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0017d] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h002fa] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h002fb] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0017e] =  I8a0037ad2845a3fbba9da380a8b8a576['h002fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0017f] =  I8a0037ad2845a3fbba9da380a8b8a576['h002fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00180] =  I8a0037ad2845a3fbba9da380a8b8a576['h00300] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00181] =  I8a0037ad2845a3fbba9da380a8b8a576['h00302] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00182] =  I8a0037ad2845a3fbba9da380a8b8a576['h00304] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00183] =  I8a0037ad2845a3fbba9da380a8b8a576['h00306] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00184] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00308] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00309] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00185] =  I8a0037ad2845a3fbba9da380a8b8a576['h0030a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00186] =  I8a0037ad2845a3fbba9da380a8b8a576['h0030c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00187] =  I8a0037ad2845a3fbba9da380a8b8a576['h0030e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00188] =  I8a0037ad2845a3fbba9da380a8b8a576['h00310] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00189] =  I8a0037ad2845a3fbba9da380a8b8a576['h00312] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0018a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00314] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0018b] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00316] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00317] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0018c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00318] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0018d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0031a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0018e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0031c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0018f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0031e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00190] =  I8a0037ad2845a3fbba9da380a8b8a576['h00320] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00191] =  I8a0037ad2845a3fbba9da380a8b8a576['h00322] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00192] =  I8a0037ad2845a3fbba9da380a8b8a576['h00324] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00193] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00326] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00327] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00194] =  I8a0037ad2845a3fbba9da380a8b8a576['h00328] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00195] =  I8a0037ad2845a3fbba9da380a8b8a576['h0032a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00196] =  I8a0037ad2845a3fbba9da380a8b8a576['h0032c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00197] =  I8a0037ad2845a3fbba9da380a8b8a576['h0032e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00198] =  I8a0037ad2845a3fbba9da380a8b8a576['h00330] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00199] =  I8a0037ad2845a3fbba9da380a8b8a576['h00332] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0019a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00334] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0019b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00336] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h0019c] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00338] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00339] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0019d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0033a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0019e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0033c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0019f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0033e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h00340] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h00342] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h00344] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h00346] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h00348] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0034a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0034c] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h001a7] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h0034e] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h0034f] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h00350] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h00352] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h00354] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h00356] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h00358] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0035a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0035c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001af] =  I8a0037ad2845a3fbba9da380a8b8a576['h0035e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h00360] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h00362] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h00364] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h00366] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h001b4] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00368] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00369] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0036a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0036c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0036e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h00370] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h00372] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h00374] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h00376] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h00378] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0037a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001be] =  I8a0037ad2845a3fbba9da380a8b8a576['h0037c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0037e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h00380] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h00382] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h00384] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h00386] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h001c4] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00388] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00389] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0038a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0038c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0038e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h00390] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h00392] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h00394] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h00396] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h00398] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0039a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0039c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0039e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h003a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h003a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h003a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h003a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h003a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h003aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h003ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h003ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h003b0] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h001d9] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h003b2] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h003b3] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001da] =  I8a0037ad2845a3fbba9da380a8b8a576['h003b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001db] =  I8a0037ad2845a3fbba9da380a8b8a576['h003b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h003b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h003ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001de] =  I8a0037ad2845a3fbba9da380a8b8a576['h003bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001df] =  I8a0037ad2845a3fbba9da380a8b8a576['h003be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h003c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h003c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h003c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h003c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h003c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h003ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h003cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h003ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h003d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h003d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h003d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h003d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h003d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h003da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h003dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h003de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h003e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h003e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h003e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h003e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h003e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h003ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h003ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h003ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h003f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h003f2] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h001fa] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h003f4] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h003f5] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h003f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h003f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h003fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h003fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h001ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h003fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00200] =  I8a0037ad2845a3fbba9da380a8b8a576['h00400] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00201] =  I8a0037ad2845a3fbba9da380a8b8a576['h00402] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00202] =  I8a0037ad2845a3fbba9da380a8b8a576['h00404] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00203] =  I8a0037ad2845a3fbba9da380a8b8a576['h00406] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00204] =  I8a0037ad2845a3fbba9da380a8b8a576['h00408] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00205] =  I8a0037ad2845a3fbba9da380a8b8a576['h0040a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00206] =  I8a0037ad2845a3fbba9da380a8b8a576['h0040c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00207] =  I8a0037ad2845a3fbba9da380a8b8a576['h0040e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00208] =  I8a0037ad2845a3fbba9da380a8b8a576['h00410] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00209] =  I8a0037ad2845a3fbba9da380a8b8a576['h00412] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0020a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00414] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0020b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00416] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0020c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00418] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0020d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0041a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0020e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0041c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0020f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0041e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00210] =  I8a0037ad2845a3fbba9da380a8b8a576['h00420] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00211] =  I8a0037ad2845a3fbba9da380a8b8a576['h00422] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00212] =  I8a0037ad2845a3fbba9da380a8b8a576['h00424] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00213] =  I8a0037ad2845a3fbba9da380a8b8a576['h00426] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00214] =  I8a0037ad2845a3fbba9da380a8b8a576['h00428] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00215] =  I8a0037ad2845a3fbba9da380a8b8a576['h0042a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00216] =  I8a0037ad2845a3fbba9da380a8b8a576['h0042c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00217] =  I8a0037ad2845a3fbba9da380a8b8a576['h0042e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00218] =  I8a0037ad2845a3fbba9da380a8b8a576['h00430] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00219] =  I8a0037ad2845a3fbba9da380a8b8a576['h00432] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0021a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00434] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0021b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00436] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0021c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00438] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0021d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0043a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0021e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0043c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0021f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0043e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00220] =  I8a0037ad2845a3fbba9da380a8b8a576['h00440] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00221] =  I8a0037ad2845a3fbba9da380a8b8a576['h00442] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00222] =  I8a0037ad2845a3fbba9da380a8b8a576['h00444] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00223] =  I8a0037ad2845a3fbba9da380a8b8a576['h00446] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00224] =  I8a0037ad2845a3fbba9da380a8b8a576['h00448] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00225] =  I8a0037ad2845a3fbba9da380a8b8a576['h0044a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00226] =  I8a0037ad2845a3fbba9da380a8b8a576['h0044c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00227] =  I8a0037ad2845a3fbba9da380a8b8a576['h0044e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00228] =  I8a0037ad2845a3fbba9da380a8b8a576['h00450] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00229] =  I8a0037ad2845a3fbba9da380a8b8a576['h00452] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0022a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00454] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0022b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00456] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0022c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00458] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0022d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0045a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0022e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0045c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0022f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0045e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00230] =  I8a0037ad2845a3fbba9da380a8b8a576['h00460] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00231] =  I8a0037ad2845a3fbba9da380a8b8a576['h00462] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00232] =  I8a0037ad2845a3fbba9da380a8b8a576['h00464] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00233] =  I8a0037ad2845a3fbba9da380a8b8a576['h00466] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00234] =  I8a0037ad2845a3fbba9da380a8b8a576['h00468] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00235] =  I8a0037ad2845a3fbba9da380a8b8a576['h0046a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00236] =  I8a0037ad2845a3fbba9da380a8b8a576['h0046c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00237] =  I8a0037ad2845a3fbba9da380a8b8a576['h0046e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00238] =  I8a0037ad2845a3fbba9da380a8b8a576['h00470] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00239] =  I8a0037ad2845a3fbba9da380a8b8a576['h00472] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0023a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00474] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0023b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00476] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0023c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00478] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0023d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0047a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0023e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0047c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0023f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0047e] ;
//end
//always_comb begin
              I0310077d53ae4ed9904df42e3f81c634['h00240] = 
          (!flogtanh_sel['h00004]) ? 
                       I8a0037ad2845a3fbba9da380a8b8a576['h00480] : //%
                       I8a0037ad2845a3fbba9da380a8b8a576['h00481] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00241] =  I8a0037ad2845a3fbba9da380a8b8a576['h00482] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00242] =  I8a0037ad2845a3fbba9da380a8b8a576['h00484] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00243] =  I8a0037ad2845a3fbba9da380a8b8a576['h00486] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00244] =  I8a0037ad2845a3fbba9da380a8b8a576['h00488] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00245] =  I8a0037ad2845a3fbba9da380a8b8a576['h0048a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00246] =  I8a0037ad2845a3fbba9da380a8b8a576['h0048c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00247] =  I8a0037ad2845a3fbba9da380a8b8a576['h0048e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00248] =  I8a0037ad2845a3fbba9da380a8b8a576['h00490] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00249] =  I8a0037ad2845a3fbba9da380a8b8a576['h00492] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0024a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00494] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0024b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00496] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0024c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00498] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0024d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0049a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0024e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0049c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0024f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0049e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00250] =  I8a0037ad2845a3fbba9da380a8b8a576['h004a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00251] =  I8a0037ad2845a3fbba9da380a8b8a576['h004a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00252] =  I8a0037ad2845a3fbba9da380a8b8a576['h004a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00253] =  I8a0037ad2845a3fbba9da380a8b8a576['h004a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00254] =  I8a0037ad2845a3fbba9da380a8b8a576['h004a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00255] =  I8a0037ad2845a3fbba9da380a8b8a576['h004aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00256] =  I8a0037ad2845a3fbba9da380a8b8a576['h004ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00257] =  I8a0037ad2845a3fbba9da380a8b8a576['h004ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00258] =  I8a0037ad2845a3fbba9da380a8b8a576['h004b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00259] =  I8a0037ad2845a3fbba9da380a8b8a576['h004b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0025a] =  I8a0037ad2845a3fbba9da380a8b8a576['h004b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0025b] =  I8a0037ad2845a3fbba9da380a8b8a576['h004b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0025c] =  I8a0037ad2845a3fbba9da380a8b8a576['h004b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0025d] =  I8a0037ad2845a3fbba9da380a8b8a576['h004ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0025e] =  I8a0037ad2845a3fbba9da380a8b8a576['h004bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0025f] =  I8a0037ad2845a3fbba9da380a8b8a576['h004be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00260] =  I8a0037ad2845a3fbba9da380a8b8a576['h004c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00261] =  I8a0037ad2845a3fbba9da380a8b8a576['h004c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00262] =  I8a0037ad2845a3fbba9da380a8b8a576['h004c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00263] =  I8a0037ad2845a3fbba9da380a8b8a576['h004c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00264] =  I8a0037ad2845a3fbba9da380a8b8a576['h004c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00265] =  I8a0037ad2845a3fbba9da380a8b8a576['h004ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00266] =  I8a0037ad2845a3fbba9da380a8b8a576['h004cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00267] =  I8a0037ad2845a3fbba9da380a8b8a576['h004ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00268] =  I8a0037ad2845a3fbba9da380a8b8a576['h004d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00269] =  I8a0037ad2845a3fbba9da380a8b8a576['h004d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0026a] =  I8a0037ad2845a3fbba9da380a8b8a576['h004d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0026b] =  I8a0037ad2845a3fbba9da380a8b8a576['h004d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0026c] =  I8a0037ad2845a3fbba9da380a8b8a576['h004d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0026d] =  I8a0037ad2845a3fbba9da380a8b8a576['h004da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0026e] =  I8a0037ad2845a3fbba9da380a8b8a576['h004dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0026f] =  I8a0037ad2845a3fbba9da380a8b8a576['h004de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00270] =  I8a0037ad2845a3fbba9da380a8b8a576['h004e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00271] =  I8a0037ad2845a3fbba9da380a8b8a576['h004e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00272] =  I8a0037ad2845a3fbba9da380a8b8a576['h004e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00273] =  I8a0037ad2845a3fbba9da380a8b8a576['h004e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00274] =  I8a0037ad2845a3fbba9da380a8b8a576['h004e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00275] =  I8a0037ad2845a3fbba9da380a8b8a576['h004ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00276] =  I8a0037ad2845a3fbba9da380a8b8a576['h004ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00277] =  I8a0037ad2845a3fbba9da380a8b8a576['h004ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00278] =  I8a0037ad2845a3fbba9da380a8b8a576['h004f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00279] =  I8a0037ad2845a3fbba9da380a8b8a576['h004f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0027a] =  I8a0037ad2845a3fbba9da380a8b8a576['h004f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0027b] =  I8a0037ad2845a3fbba9da380a8b8a576['h004f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0027c] =  I8a0037ad2845a3fbba9da380a8b8a576['h004f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0027d] =  I8a0037ad2845a3fbba9da380a8b8a576['h004fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0027e] =  I8a0037ad2845a3fbba9da380a8b8a576['h004fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0027f] =  I8a0037ad2845a3fbba9da380a8b8a576['h004fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00280] =  I8a0037ad2845a3fbba9da380a8b8a576['h00500] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00281] =  I8a0037ad2845a3fbba9da380a8b8a576['h00502] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00282] =  I8a0037ad2845a3fbba9da380a8b8a576['h00504] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00283] =  I8a0037ad2845a3fbba9da380a8b8a576['h00506] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00284] =  I8a0037ad2845a3fbba9da380a8b8a576['h00508] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00285] =  I8a0037ad2845a3fbba9da380a8b8a576['h0050a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00286] =  I8a0037ad2845a3fbba9da380a8b8a576['h0050c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00287] =  I8a0037ad2845a3fbba9da380a8b8a576['h0050e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00288] =  I8a0037ad2845a3fbba9da380a8b8a576['h00510] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00289] =  I8a0037ad2845a3fbba9da380a8b8a576['h00512] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0028a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00514] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0028b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00516] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0028c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00518] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0028d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0051a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0028e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0051c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0028f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0051e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00290] =  I8a0037ad2845a3fbba9da380a8b8a576['h00520] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00291] =  I8a0037ad2845a3fbba9da380a8b8a576['h00522] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00292] =  I8a0037ad2845a3fbba9da380a8b8a576['h00524] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00293] =  I8a0037ad2845a3fbba9da380a8b8a576['h00526] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00294] =  I8a0037ad2845a3fbba9da380a8b8a576['h00528] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00295] =  I8a0037ad2845a3fbba9da380a8b8a576['h0052a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00296] =  I8a0037ad2845a3fbba9da380a8b8a576['h0052c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00297] =  I8a0037ad2845a3fbba9da380a8b8a576['h0052e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00298] =  I8a0037ad2845a3fbba9da380a8b8a576['h00530] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00299] =  I8a0037ad2845a3fbba9da380a8b8a576['h00532] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0029a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00534] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0029b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00536] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0029c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00538] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0029d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0053a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0029e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0053c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0029f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0053e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h00540] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h00542] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h00544] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h00546] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h00548] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0054a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0054c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0054e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h00550] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h00552] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h00554] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h00556] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h00558] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0055a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0055c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002af] =  I8a0037ad2845a3fbba9da380a8b8a576['h0055e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h00560] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h00562] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h00564] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h00566] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h00568] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0056a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0056c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0056e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h00570] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h00572] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h00574] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h00576] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h00578] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0057a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002be] =  I8a0037ad2845a3fbba9da380a8b8a576['h0057c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0057e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h00580] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h00582] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h00584] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h00586] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h00588] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0058a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0058c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0058e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h00590] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h00592] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h00594] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h00596] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h00598] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0059a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0059c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0059e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h005a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h005a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h005a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h005a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h005a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h005aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h005ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h005ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h005b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h005b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002da] =  I8a0037ad2845a3fbba9da380a8b8a576['h005b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002db] =  I8a0037ad2845a3fbba9da380a8b8a576['h005b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h005b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h005ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002de] =  I8a0037ad2845a3fbba9da380a8b8a576['h005bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002df] =  I8a0037ad2845a3fbba9da380a8b8a576['h005be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h005c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h005c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h005c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h005c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h005c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h005ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h005cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h005ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h005d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h005d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h005d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h005d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h005d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h005da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h005dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h005de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h005e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h005e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h005e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h005e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h005e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h005ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h005ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h005ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h005f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h005f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h005f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h005f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h005f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h005fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h005fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h002ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h005fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00300] =  I8a0037ad2845a3fbba9da380a8b8a576['h00600] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00301] =  I8a0037ad2845a3fbba9da380a8b8a576['h00602] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00302] =  I8a0037ad2845a3fbba9da380a8b8a576['h00604] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00303] =  I8a0037ad2845a3fbba9da380a8b8a576['h00606] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00304] =  I8a0037ad2845a3fbba9da380a8b8a576['h00608] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00305] =  I8a0037ad2845a3fbba9da380a8b8a576['h0060a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00306] =  I8a0037ad2845a3fbba9da380a8b8a576['h0060c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00307] =  I8a0037ad2845a3fbba9da380a8b8a576['h0060e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00308] =  I8a0037ad2845a3fbba9da380a8b8a576['h00610] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00309] =  I8a0037ad2845a3fbba9da380a8b8a576['h00612] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0030a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00614] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0030b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00616] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0030c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00618] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0030d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0061a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0030e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0061c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0030f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0061e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00310] =  I8a0037ad2845a3fbba9da380a8b8a576['h00620] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00311] =  I8a0037ad2845a3fbba9da380a8b8a576['h00622] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00312] =  I8a0037ad2845a3fbba9da380a8b8a576['h00624] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00313] =  I8a0037ad2845a3fbba9da380a8b8a576['h00626] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00314] =  I8a0037ad2845a3fbba9da380a8b8a576['h00628] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00315] =  I8a0037ad2845a3fbba9da380a8b8a576['h0062a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00316] =  I8a0037ad2845a3fbba9da380a8b8a576['h0062c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00317] =  I8a0037ad2845a3fbba9da380a8b8a576['h0062e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00318] =  I8a0037ad2845a3fbba9da380a8b8a576['h00630] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00319] =  I8a0037ad2845a3fbba9da380a8b8a576['h00632] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0031a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00634] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0031b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00636] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0031c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00638] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0031d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0063a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0031e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0063c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0031f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0063e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00320] =  I8a0037ad2845a3fbba9da380a8b8a576['h00640] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00321] =  I8a0037ad2845a3fbba9da380a8b8a576['h00642] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00322] =  I8a0037ad2845a3fbba9da380a8b8a576['h00644] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00323] =  I8a0037ad2845a3fbba9da380a8b8a576['h00646] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00324] =  I8a0037ad2845a3fbba9da380a8b8a576['h00648] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00325] =  I8a0037ad2845a3fbba9da380a8b8a576['h0064a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00326] =  I8a0037ad2845a3fbba9da380a8b8a576['h0064c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00327] =  I8a0037ad2845a3fbba9da380a8b8a576['h0064e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00328] =  I8a0037ad2845a3fbba9da380a8b8a576['h00650] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00329] =  I8a0037ad2845a3fbba9da380a8b8a576['h00652] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0032a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00654] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0032b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00656] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0032c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00658] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0032d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0065a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0032e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0065c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0032f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0065e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00330] =  I8a0037ad2845a3fbba9da380a8b8a576['h00660] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00331] =  I8a0037ad2845a3fbba9da380a8b8a576['h00662] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00332] =  I8a0037ad2845a3fbba9da380a8b8a576['h00664] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00333] =  I8a0037ad2845a3fbba9da380a8b8a576['h00666] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00334] =  I8a0037ad2845a3fbba9da380a8b8a576['h00668] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00335] =  I8a0037ad2845a3fbba9da380a8b8a576['h0066a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00336] =  I8a0037ad2845a3fbba9da380a8b8a576['h0066c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00337] =  I8a0037ad2845a3fbba9da380a8b8a576['h0066e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00338] =  I8a0037ad2845a3fbba9da380a8b8a576['h00670] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00339] =  I8a0037ad2845a3fbba9da380a8b8a576['h00672] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0033a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00674] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0033b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00676] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0033c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00678] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0033d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0067a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0033e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0067c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0033f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0067e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00340] =  I8a0037ad2845a3fbba9da380a8b8a576['h00680] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00341] =  I8a0037ad2845a3fbba9da380a8b8a576['h00682] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00342] =  I8a0037ad2845a3fbba9da380a8b8a576['h00684] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00343] =  I8a0037ad2845a3fbba9da380a8b8a576['h00686] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00344] =  I8a0037ad2845a3fbba9da380a8b8a576['h00688] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00345] =  I8a0037ad2845a3fbba9da380a8b8a576['h0068a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00346] =  I8a0037ad2845a3fbba9da380a8b8a576['h0068c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00347] =  I8a0037ad2845a3fbba9da380a8b8a576['h0068e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00348] =  I8a0037ad2845a3fbba9da380a8b8a576['h00690] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00349] =  I8a0037ad2845a3fbba9da380a8b8a576['h00692] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0034a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00694] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0034b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00696] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0034c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00698] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0034d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0069a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0034e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0069c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0034f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0069e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00350] =  I8a0037ad2845a3fbba9da380a8b8a576['h006a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00351] =  I8a0037ad2845a3fbba9da380a8b8a576['h006a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00352] =  I8a0037ad2845a3fbba9da380a8b8a576['h006a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00353] =  I8a0037ad2845a3fbba9da380a8b8a576['h006a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00354] =  I8a0037ad2845a3fbba9da380a8b8a576['h006a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00355] =  I8a0037ad2845a3fbba9da380a8b8a576['h006aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00356] =  I8a0037ad2845a3fbba9da380a8b8a576['h006ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00357] =  I8a0037ad2845a3fbba9da380a8b8a576['h006ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00358] =  I8a0037ad2845a3fbba9da380a8b8a576['h006b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00359] =  I8a0037ad2845a3fbba9da380a8b8a576['h006b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0035a] =  I8a0037ad2845a3fbba9da380a8b8a576['h006b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0035b] =  I8a0037ad2845a3fbba9da380a8b8a576['h006b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0035c] =  I8a0037ad2845a3fbba9da380a8b8a576['h006b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0035d] =  I8a0037ad2845a3fbba9da380a8b8a576['h006ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0035e] =  I8a0037ad2845a3fbba9da380a8b8a576['h006bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0035f] =  I8a0037ad2845a3fbba9da380a8b8a576['h006be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00360] =  I8a0037ad2845a3fbba9da380a8b8a576['h006c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00361] =  I8a0037ad2845a3fbba9da380a8b8a576['h006c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00362] =  I8a0037ad2845a3fbba9da380a8b8a576['h006c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00363] =  I8a0037ad2845a3fbba9da380a8b8a576['h006c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00364] =  I8a0037ad2845a3fbba9da380a8b8a576['h006c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00365] =  I8a0037ad2845a3fbba9da380a8b8a576['h006ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00366] =  I8a0037ad2845a3fbba9da380a8b8a576['h006cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00367] =  I8a0037ad2845a3fbba9da380a8b8a576['h006ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00368] =  I8a0037ad2845a3fbba9da380a8b8a576['h006d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00369] =  I8a0037ad2845a3fbba9da380a8b8a576['h006d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0036a] =  I8a0037ad2845a3fbba9da380a8b8a576['h006d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0036b] =  I8a0037ad2845a3fbba9da380a8b8a576['h006d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0036c] =  I8a0037ad2845a3fbba9da380a8b8a576['h006d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0036d] =  I8a0037ad2845a3fbba9da380a8b8a576['h006da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0036e] =  I8a0037ad2845a3fbba9da380a8b8a576['h006dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0036f] =  I8a0037ad2845a3fbba9da380a8b8a576['h006de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00370] =  I8a0037ad2845a3fbba9da380a8b8a576['h006e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00371] =  I8a0037ad2845a3fbba9da380a8b8a576['h006e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00372] =  I8a0037ad2845a3fbba9da380a8b8a576['h006e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00373] =  I8a0037ad2845a3fbba9da380a8b8a576['h006e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00374] =  I8a0037ad2845a3fbba9da380a8b8a576['h006e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00375] =  I8a0037ad2845a3fbba9da380a8b8a576['h006ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00376] =  I8a0037ad2845a3fbba9da380a8b8a576['h006ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00377] =  I8a0037ad2845a3fbba9da380a8b8a576['h006ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00378] =  I8a0037ad2845a3fbba9da380a8b8a576['h006f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00379] =  I8a0037ad2845a3fbba9da380a8b8a576['h006f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0037a] =  I8a0037ad2845a3fbba9da380a8b8a576['h006f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0037b] =  I8a0037ad2845a3fbba9da380a8b8a576['h006f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0037c] =  I8a0037ad2845a3fbba9da380a8b8a576['h006f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0037d] =  I8a0037ad2845a3fbba9da380a8b8a576['h006fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0037e] =  I8a0037ad2845a3fbba9da380a8b8a576['h006fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0037f] =  I8a0037ad2845a3fbba9da380a8b8a576['h006fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00380] =  I8a0037ad2845a3fbba9da380a8b8a576['h00700] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00381] =  I8a0037ad2845a3fbba9da380a8b8a576['h00702] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00382] =  I8a0037ad2845a3fbba9da380a8b8a576['h00704] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00383] =  I8a0037ad2845a3fbba9da380a8b8a576['h00706] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00384] =  I8a0037ad2845a3fbba9da380a8b8a576['h00708] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00385] =  I8a0037ad2845a3fbba9da380a8b8a576['h0070a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00386] =  I8a0037ad2845a3fbba9da380a8b8a576['h0070c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00387] =  I8a0037ad2845a3fbba9da380a8b8a576['h0070e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00388] =  I8a0037ad2845a3fbba9da380a8b8a576['h00710] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00389] =  I8a0037ad2845a3fbba9da380a8b8a576['h00712] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0038a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00714] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0038b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00716] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0038c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00718] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0038d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0071a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0038e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0071c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0038f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0071e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00390] =  I8a0037ad2845a3fbba9da380a8b8a576['h00720] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00391] =  I8a0037ad2845a3fbba9da380a8b8a576['h00722] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00392] =  I8a0037ad2845a3fbba9da380a8b8a576['h00724] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00393] =  I8a0037ad2845a3fbba9da380a8b8a576['h00726] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00394] =  I8a0037ad2845a3fbba9da380a8b8a576['h00728] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00395] =  I8a0037ad2845a3fbba9da380a8b8a576['h0072a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00396] =  I8a0037ad2845a3fbba9da380a8b8a576['h0072c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00397] =  I8a0037ad2845a3fbba9da380a8b8a576['h0072e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00398] =  I8a0037ad2845a3fbba9da380a8b8a576['h00730] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00399] =  I8a0037ad2845a3fbba9da380a8b8a576['h00732] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0039a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00734] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0039b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00736] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0039c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00738] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0039d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0073a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0039e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0073c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0039f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0073e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h00740] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h00742] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h00744] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h00746] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h00748] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0074a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0074c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0074e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h00750] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h00752] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h00754] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h00756] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h00758] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0075a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0075c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003af] =  I8a0037ad2845a3fbba9da380a8b8a576['h0075e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h00760] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h00762] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h00764] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h00766] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h00768] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0076a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0076c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0076e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h00770] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h00772] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h00774] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h00776] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h00778] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0077a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003be] =  I8a0037ad2845a3fbba9da380a8b8a576['h0077c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0077e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h00780] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h00782] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h00784] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h00786] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h00788] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0078a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0078c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0078e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h00790] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h00792] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h00794] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h00796] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h00798] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0079a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0079c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0079e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h007a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h007a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h007a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h007a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h007a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h007aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h007ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h007ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h007b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h007b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003da] =  I8a0037ad2845a3fbba9da380a8b8a576['h007b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003db] =  I8a0037ad2845a3fbba9da380a8b8a576['h007b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h007b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h007ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003de] =  I8a0037ad2845a3fbba9da380a8b8a576['h007bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003df] =  I8a0037ad2845a3fbba9da380a8b8a576['h007be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h007c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h007c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h007c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h007c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h007c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h007ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h007cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h007ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h007d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h007d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h007d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h007d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h007d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h007da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h007dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h007de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h007e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h007e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h007e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h007e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h007e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h007ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h007ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h007ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h007f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h007f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h007f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h007f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h007f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h007fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h007fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h003ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h007fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00400] =  I8a0037ad2845a3fbba9da380a8b8a576['h00800] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00401] =  I8a0037ad2845a3fbba9da380a8b8a576['h00802] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00402] =  I8a0037ad2845a3fbba9da380a8b8a576['h00804] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00403] =  I8a0037ad2845a3fbba9da380a8b8a576['h00806] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00404] =  I8a0037ad2845a3fbba9da380a8b8a576['h00808] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00405] =  I8a0037ad2845a3fbba9da380a8b8a576['h0080a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00406] =  I8a0037ad2845a3fbba9da380a8b8a576['h0080c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00407] =  I8a0037ad2845a3fbba9da380a8b8a576['h0080e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00408] =  I8a0037ad2845a3fbba9da380a8b8a576['h00810] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00409] =  I8a0037ad2845a3fbba9da380a8b8a576['h00812] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0040a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00814] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0040b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00816] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0040c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00818] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0040d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0081a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0040e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0081c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0040f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0081e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00410] =  I8a0037ad2845a3fbba9da380a8b8a576['h00820] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00411] =  I8a0037ad2845a3fbba9da380a8b8a576['h00822] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00412] =  I8a0037ad2845a3fbba9da380a8b8a576['h00824] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00413] =  I8a0037ad2845a3fbba9da380a8b8a576['h00826] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00414] =  I8a0037ad2845a3fbba9da380a8b8a576['h00828] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00415] =  I8a0037ad2845a3fbba9da380a8b8a576['h0082a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00416] =  I8a0037ad2845a3fbba9da380a8b8a576['h0082c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00417] =  I8a0037ad2845a3fbba9da380a8b8a576['h0082e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00418] =  I8a0037ad2845a3fbba9da380a8b8a576['h00830] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00419] =  I8a0037ad2845a3fbba9da380a8b8a576['h00832] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0041a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00834] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0041b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00836] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0041c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00838] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0041d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0083a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0041e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0083c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0041f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0083e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00420] =  I8a0037ad2845a3fbba9da380a8b8a576['h00840] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00421] =  I8a0037ad2845a3fbba9da380a8b8a576['h00842] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00422] =  I8a0037ad2845a3fbba9da380a8b8a576['h00844] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00423] =  I8a0037ad2845a3fbba9da380a8b8a576['h00846] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00424] =  I8a0037ad2845a3fbba9da380a8b8a576['h00848] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00425] =  I8a0037ad2845a3fbba9da380a8b8a576['h0084a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00426] =  I8a0037ad2845a3fbba9da380a8b8a576['h0084c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00427] =  I8a0037ad2845a3fbba9da380a8b8a576['h0084e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00428] =  I8a0037ad2845a3fbba9da380a8b8a576['h00850] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00429] =  I8a0037ad2845a3fbba9da380a8b8a576['h00852] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0042a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00854] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0042b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00856] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0042c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00858] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0042d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0085a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0042e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0085c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0042f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0085e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00430] =  I8a0037ad2845a3fbba9da380a8b8a576['h00860] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00431] =  I8a0037ad2845a3fbba9da380a8b8a576['h00862] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00432] =  I8a0037ad2845a3fbba9da380a8b8a576['h00864] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00433] =  I8a0037ad2845a3fbba9da380a8b8a576['h00866] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00434] =  I8a0037ad2845a3fbba9da380a8b8a576['h00868] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00435] =  I8a0037ad2845a3fbba9da380a8b8a576['h0086a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00436] =  I8a0037ad2845a3fbba9da380a8b8a576['h0086c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00437] =  I8a0037ad2845a3fbba9da380a8b8a576['h0086e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00438] =  I8a0037ad2845a3fbba9da380a8b8a576['h00870] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00439] =  I8a0037ad2845a3fbba9da380a8b8a576['h00872] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0043a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00874] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0043b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00876] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0043c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00878] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0043d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0087a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0043e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0087c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0043f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0087e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00440] =  I8a0037ad2845a3fbba9da380a8b8a576['h00880] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00441] =  I8a0037ad2845a3fbba9da380a8b8a576['h00882] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00442] =  I8a0037ad2845a3fbba9da380a8b8a576['h00884] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00443] =  I8a0037ad2845a3fbba9da380a8b8a576['h00886] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00444] =  I8a0037ad2845a3fbba9da380a8b8a576['h00888] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00445] =  I8a0037ad2845a3fbba9da380a8b8a576['h0088a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00446] =  I8a0037ad2845a3fbba9da380a8b8a576['h0088c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00447] =  I8a0037ad2845a3fbba9da380a8b8a576['h0088e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00448] =  I8a0037ad2845a3fbba9da380a8b8a576['h00890] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00449] =  I8a0037ad2845a3fbba9da380a8b8a576['h00892] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0044a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00894] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0044b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00896] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0044c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00898] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0044d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0089a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0044e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0089c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0044f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0089e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00450] =  I8a0037ad2845a3fbba9da380a8b8a576['h008a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00451] =  I8a0037ad2845a3fbba9da380a8b8a576['h008a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00452] =  I8a0037ad2845a3fbba9da380a8b8a576['h008a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00453] =  I8a0037ad2845a3fbba9da380a8b8a576['h008a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00454] =  I8a0037ad2845a3fbba9da380a8b8a576['h008a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00455] =  I8a0037ad2845a3fbba9da380a8b8a576['h008aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00456] =  I8a0037ad2845a3fbba9da380a8b8a576['h008ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00457] =  I8a0037ad2845a3fbba9da380a8b8a576['h008ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00458] =  I8a0037ad2845a3fbba9da380a8b8a576['h008b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00459] =  I8a0037ad2845a3fbba9da380a8b8a576['h008b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0045a] =  I8a0037ad2845a3fbba9da380a8b8a576['h008b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0045b] =  I8a0037ad2845a3fbba9da380a8b8a576['h008b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0045c] =  I8a0037ad2845a3fbba9da380a8b8a576['h008b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0045d] =  I8a0037ad2845a3fbba9da380a8b8a576['h008ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0045e] =  I8a0037ad2845a3fbba9da380a8b8a576['h008bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0045f] =  I8a0037ad2845a3fbba9da380a8b8a576['h008be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00460] =  I8a0037ad2845a3fbba9da380a8b8a576['h008c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00461] =  I8a0037ad2845a3fbba9da380a8b8a576['h008c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00462] =  I8a0037ad2845a3fbba9da380a8b8a576['h008c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00463] =  I8a0037ad2845a3fbba9da380a8b8a576['h008c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00464] =  I8a0037ad2845a3fbba9da380a8b8a576['h008c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00465] =  I8a0037ad2845a3fbba9da380a8b8a576['h008ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00466] =  I8a0037ad2845a3fbba9da380a8b8a576['h008cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00467] =  I8a0037ad2845a3fbba9da380a8b8a576['h008ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00468] =  I8a0037ad2845a3fbba9da380a8b8a576['h008d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00469] =  I8a0037ad2845a3fbba9da380a8b8a576['h008d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0046a] =  I8a0037ad2845a3fbba9da380a8b8a576['h008d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0046b] =  I8a0037ad2845a3fbba9da380a8b8a576['h008d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0046c] =  I8a0037ad2845a3fbba9da380a8b8a576['h008d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0046d] =  I8a0037ad2845a3fbba9da380a8b8a576['h008da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0046e] =  I8a0037ad2845a3fbba9da380a8b8a576['h008dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0046f] =  I8a0037ad2845a3fbba9da380a8b8a576['h008de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00470] =  I8a0037ad2845a3fbba9da380a8b8a576['h008e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00471] =  I8a0037ad2845a3fbba9da380a8b8a576['h008e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00472] =  I8a0037ad2845a3fbba9da380a8b8a576['h008e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00473] =  I8a0037ad2845a3fbba9da380a8b8a576['h008e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00474] =  I8a0037ad2845a3fbba9da380a8b8a576['h008e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00475] =  I8a0037ad2845a3fbba9da380a8b8a576['h008ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00476] =  I8a0037ad2845a3fbba9da380a8b8a576['h008ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00477] =  I8a0037ad2845a3fbba9da380a8b8a576['h008ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00478] =  I8a0037ad2845a3fbba9da380a8b8a576['h008f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00479] =  I8a0037ad2845a3fbba9da380a8b8a576['h008f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0047a] =  I8a0037ad2845a3fbba9da380a8b8a576['h008f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0047b] =  I8a0037ad2845a3fbba9da380a8b8a576['h008f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0047c] =  I8a0037ad2845a3fbba9da380a8b8a576['h008f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0047d] =  I8a0037ad2845a3fbba9da380a8b8a576['h008fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0047e] =  I8a0037ad2845a3fbba9da380a8b8a576['h008fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0047f] =  I8a0037ad2845a3fbba9da380a8b8a576['h008fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00480] =  I8a0037ad2845a3fbba9da380a8b8a576['h00900] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00481] =  I8a0037ad2845a3fbba9da380a8b8a576['h00902] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00482] =  I8a0037ad2845a3fbba9da380a8b8a576['h00904] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00483] =  I8a0037ad2845a3fbba9da380a8b8a576['h00906] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00484] =  I8a0037ad2845a3fbba9da380a8b8a576['h00908] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00485] =  I8a0037ad2845a3fbba9da380a8b8a576['h0090a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00486] =  I8a0037ad2845a3fbba9da380a8b8a576['h0090c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00487] =  I8a0037ad2845a3fbba9da380a8b8a576['h0090e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00488] =  I8a0037ad2845a3fbba9da380a8b8a576['h00910] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00489] =  I8a0037ad2845a3fbba9da380a8b8a576['h00912] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0048a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00914] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0048b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00916] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0048c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00918] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0048d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0091a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0048e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0091c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0048f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0091e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00490] =  I8a0037ad2845a3fbba9da380a8b8a576['h00920] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00491] =  I8a0037ad2845a3fbba9da380a8b8a576['h00922] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00492] =  I8a0037ad2845a3fbba9da380a8b8a576['h00924] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00493] =  I8a0037ad2845a3fbba9da380a8b8a576['h00926] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00494] =  I8a0037ad2845a3fbba9da380a8b8a576['h00928] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00495] =  I8a0037ad2845a3fbba9da380a8b8a576['h0092a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00496] =  I8a0037ad2845a3fbba9da380a8b8a576['h0092c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00497] =  I8a0037ad2845a3fbba9da380a8b8a576['h0092e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00498] =  I8a0037ad2845a3fbba9da380a8b8a576['h00930] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00499] =  I8a0037ad2845a3fbba9da380a8b8a576['h00932] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0049a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00934] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0049b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00936] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0049c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00938] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0049d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0093a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0049e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0093c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0049f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0093e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h00940] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h00942] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h00944] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h00946] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h00948] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0094a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0094c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0094e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h00950] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h00952] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h00954] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h00956] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h00958] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0095a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0095c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004af] =  I8a0037ad2845a3fbba9da380a8b8a576['h0095e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h00960] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h00962] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h00964] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h00966] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h00968] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0096a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0096c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0096e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h00970] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h00972] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h00974] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h00976] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h00978] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0097a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004be] =  I8a0037ad2845a3fbba9da380a8b8a576['h0097c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0097e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h00980] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h00982] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h00984] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h00986] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h00988] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0098a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0098c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0098e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h00990] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h00992] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h00994] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h00996] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h00998] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0099a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0099c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0099e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h009a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h009a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h009a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h009a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h009a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h009aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h009ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h009ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h009b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h009b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004da] =  I8a0037ad2845a3fbba9da380a8b8a576['h009b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004db] =  I8a0037ad2845a3fbba9da380a8b8a576['h009b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h009b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h009ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004de] =  I8a0037ad2845a3fbba9da380a8b8a576['h009bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004df] =  I8a0037ad2845a3fbba9da380a8b8a576['h009be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h009c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h009c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h009c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h009c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h009c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h009ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h009cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h009ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h009d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h009d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h009d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h009d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h009d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h009da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h009dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h009de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h009e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h009e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h009e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h009e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h009e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h009ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h009ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h009ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h009f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h009f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h009f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h009f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h009f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h009fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h009fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h004ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h009fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00500] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00501] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00502] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00503] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00504] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00505] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00506] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00507] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00508] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00509] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0050a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0050b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0050c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0050d] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0050e] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0050f] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00510] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00511] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00512] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00513] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00514] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00515] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00516] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00517] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00518] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00519] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0051a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0051b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0051c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0051d] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0051e] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0051f] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00520] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00521] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00522] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00523] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00524] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00525] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00526] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00527] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00528] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00529] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0052a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0052b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0052c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0052d] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0052e] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0052f] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00530] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00531] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00532] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00533] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00534] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00535] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00536] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00537] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00538] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00539] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0053a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0053b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0053c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0053d] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0053e] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0053f] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00540] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00541] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00542] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00543] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00544] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00545] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00546] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00547] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00548] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00549] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0054a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0054b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0054c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0054d] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0054e] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0054f] =  I8a0037ad2845a3fbba9da380a8b8a576['h00a9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00550] =  I8a0037ad2845a3fbba9da380a8b8a576['h00aa0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00551] =  I8a0037ad2845a3fbba9da380a8b8a576['h00aa2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00552] =  I8a0037ad2845a3fbba9da380a8b8a576['h00aa4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00553] =  I8a0037ad2845a3fbba9da380a8b8a576['h00aa6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00554] =  I8a0037ad2845a3fbba9da380a8b8a576['h00aa8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00555] =  I8a0037ad2845a3fbba9da380a8b8a576['h00aaa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00556] =  I8a0037ad2845a3fbba9da380a8b8a576['h00aac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00557] =  I8a0037ad2845a3fbba9da380a8b8a576['h00aae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00558] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ab0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00559] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ab2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0055a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ab4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0055b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ab6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0055c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ab8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0055d] =  I8a0037ad2845a3fbba9da380a8b8a576['h00aba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0055e] =  I8a0037ad2845a3fbba9da380a8b8a576['h00abc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0055f] =  I8a0037ad2845a3fbba9da380a8b8a576['h00abe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00560] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ac0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00561] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ac2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00562] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ac4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00563] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ac6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00564] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ac8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00565] =  I8a0037ad2845a3fbba9da380a8b8a576['h00aca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00566] =  I8a0037ad2845a3fbba9da380a8b8a576['h00acc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00567] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ace] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00568] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ad0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00569] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ad2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0056a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ad4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0056b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ad6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0056c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ad8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0056d] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ada] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0056e] =  I8a0037ad2845a3fbba9da380a8b8a576['h00adc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0056f] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ade] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00570] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ae0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00571] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ae2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00572] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ae4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00573] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ae6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00574] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ae8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00575] =  I8a0037ad2845a3fbba9da380a8b8a576['h00aea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00576] =  I8a0037ad2845a3fbba9da380a8b8a576['h00aec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00577] =  I8a0037ad2845a3fbba9da380a8b8a576['h00aee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00578] =  I8a0037ad2845a3fbba9da380a8b8a576['h00af0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00579] =  I8a0037ad2845a3fbba9da380a8b8a576['h00af2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0057a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00af4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0057b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00af6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0057c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00af8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0057d] =  I8a0037ad2845a3fbba9da380a8b8a576['h00afa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0057e] =  I8a0037ad2845a3fbba9da380a8b8a576['h00afc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0057f] =  I8a0037ad2845a3fbba9da380a8b8a576['h00afe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00580] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00581] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00582] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00583] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00584] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00585] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00586] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00587] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00588] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00589] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0058a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0058b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0058c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0058d] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0058e] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0058f] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00590] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00591] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00592] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00593] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00594] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00595] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00596] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00597] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00598] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00599] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0059a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0059b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0059c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0059d] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0059e] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0059f] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005af] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005be] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h00b9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ba0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ba2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ba4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ba6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ba8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h00baa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005da] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005db] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005de] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005df] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bcc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bdc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h00be0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h00be2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h00be4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h00be6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h00be8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bf0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bf2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bf4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bf6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bf8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bfa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bfc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h005ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h00bfe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00600] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00601] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00602] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00603] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00604] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00605] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00606] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00607] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00608] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00609] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0060a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0060b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0060c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0060d] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0060e] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0060f] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00610] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00611] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00612] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00613] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00614] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00615] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00616] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00617] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00618] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00619] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0061a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0061b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0061c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0061d] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0061e] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0061f] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00620] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00621] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00622] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00623] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00624] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00625] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00626] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00627] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00628] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00629] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0062a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0062b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0062c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0062d] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0062e] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0062f] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00630] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00631] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00632] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00633] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00634] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00635] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00636] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00637] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00638] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00639] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0063a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0063b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0063c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0063d] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0063e] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0063f] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00640] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00641] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00642] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00643] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00644] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00645] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00646] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00647] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00648] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00649] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0064a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0064b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0064c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0064d] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0064e] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0064f] =  I8a0037ad2845a3fbba9da380a8b8a576['h00c9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00650] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ca0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00651] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ca2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00652] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ca4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00653] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ca6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00654] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ca8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00655] =  I8a0037ad2845a3fbba9da380a8b8a576['h00caa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00656] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00657] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00658] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00659] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0065a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0065b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0065c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0065d] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0065e] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0065f] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00660] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00661] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00662] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00663] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00664] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00665] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00666] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ccc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00667] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00668] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00669] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0066a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0066b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0066c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0066d] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0066e] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cdc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0066f] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00670] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ce0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00671] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ce2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00672] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ce4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00673] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ce6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00674] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ce8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00675] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00676] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00677] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00678] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cf0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00679] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cf2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0067a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cf4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0067b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cf6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0067c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cf8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0067d] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cfa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0067e] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cfc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0067f] =  I8a0037ad2845a3fbba9da380a8b8a576['h00cfe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00680] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00681] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00682] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00683] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00684] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00685] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00686] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00687] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00688] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00689] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0068a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0068b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0068c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0068d] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0068e] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0068f] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00690] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00691] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00692] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00693] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00694] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00695] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00696] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00697] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00698] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00699] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0069a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0069b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0069c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0069d] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0069e] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0069f] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006af] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006be] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h00d9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h00da0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h00da2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h00da4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h00da6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h00da8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h00daa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h00dac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h00dae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h00db0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h00db2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006da] =  I8a0037ad2845a3fbba9da380a8b8a576['h00db4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006db] =  I8a0037ad2845a3fbba9da380a8b8a576['h00db6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h00db8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h00dba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006de] =  I8a0037ad2845a3fbba9da380a8b8a576['h00dbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006df] =  I8a0037ad2845a3fbba9da380a8b8a576['h00dbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h00dc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h00dc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h00dc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h00dc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h00dc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h00dca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h00dcc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h00dce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h00dd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h00dd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h00dd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h00dd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h00dd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h00dda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ddc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h00dde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h00de0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h00de2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h00de4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h00de6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h00de8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h00dea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h00dec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h00dee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h00df0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h00df2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h00df4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h00df6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h00df8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h00dfa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h00dfc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h006ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h00dfe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00700] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00701] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00702] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00703] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00704] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00705] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00706] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00707] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00708] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00709] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0070a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0070b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0070c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0070d] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0070e] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0070f] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00710] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00711] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00712] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00713] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00714] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00715] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00716] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00717] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00718] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00719] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0071a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0071b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0071c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0071d] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0071e] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0071f] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00720] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00721] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00722] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00723] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00724] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00725] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00726] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00727] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00728] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00729] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0072a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0072b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0072c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0072d] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0072e] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0072f] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00730] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00731] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00732] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00733] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00734] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00735] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00736] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00737] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00738] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00739] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0073a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0073b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0073c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0073d] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0073e] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0073f] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00740] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00741] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00742] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00743] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00744] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00745] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00746] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00747] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00748] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00749] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0074a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0074b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0074c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0074d] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0074e] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0074f] =  I8a0037ad2845a3fbba9da380a8b8a576['h00e9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00750] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ea0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00751] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ea2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00752] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ea4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00753] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ea6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00754] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ea8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00755] =  I8a0037ad2845a3fbba9da380a8b8a576['h00eaa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00756] =  I8a0037ad2845a3fbba9da380a8b8a576['h00eac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00757] =  I8a0037ad2845a3fbba9da380a8b8a576['h00eae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00758] =  I8a0037ad2845a3fbba9da380a8b8a576['h00eb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00759] =  I8a0037ad2845a3fbba9da380a8b8a576['h00eb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0075a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00eb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0075b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00eb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0075c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00eb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0075d] =  I8a0037ad2845a3fbba9da380a8b8a576['h00eba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0075e] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ebc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0075f] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ebe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00760] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ec0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00761] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ec2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00762] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ec4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00763] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ec6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00764] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ec8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00765] =  I8a0037ad2845a3fbba9da380a8b8a576['h00eca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00766] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ecc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00767] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ece] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00768] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ed0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00769] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ed2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0076a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ed4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0076b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ed6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0076c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ed8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0076d] =  I8a0037ad2845a3fbba9da380a8b8a576['h00eda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0076e] =  I8a0037ad2845a3fbba9da380a8b8a576['h00edc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0076f] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ede] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00770] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ee0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00771] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ee2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00772] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ee4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00773] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ee6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00774] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ee8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00775] =  I8a0037ad2845a3fbba9da380a8b8a576['h00eea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00776] =  I8a0037ad2845a3fbba9da380a8b8a576['h00eec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00777] =  I8a0037ad2845a3fbba9da380a8b8a576['h00eee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00778] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ef0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00779] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ef2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0077a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ef4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0077b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ef6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0077c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ef8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0077d] =  I8a0037ad2845a3fbba9da380a8b8a576['h00efa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0077e] =  I8a0037ad2845a3fbba9da380a8b8a576['h00efc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0077f] =  I8a0037ad2845a3fbba9da380a8b8a576['h00efe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00780] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00781] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00782] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00783] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00784] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00785] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00786] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00787] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00788] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00789] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0078a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0078b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0078c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0078d] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0078e] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0078f] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00790] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00791] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00792] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00793] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00794] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00795] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00796] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00797] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00798] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00799] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0079a] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0079b] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0079c] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0079d] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0079e] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0079f] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007af] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007be] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h00f9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fa0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fa2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fa4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fa6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fa8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h00faa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007da] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007db] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007de] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007df] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fcc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fdc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fe0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fe2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fe4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fe6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fe8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h00fee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ff0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ff2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ff4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ff6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ff8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ffa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ffc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h007ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h00ffe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00800] =  I8a0037ad2845a3fbba9da380a8b8a576['h01000] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00801] =  I8a0037ad2845a3fbba9da380a8b8a576['h01002] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00802] =  I8a0037ad2845a3fbba9da380a8b8a576['h01004] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00803] =  I8a0037ad2845a3fbba9da380a8b8a576['h01006] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00804] =  I8a0037ad2845a3fbba9da380a8b8a576['h01008] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00805] =  I8a0037ad2845a3fbba9da380a8b8a576['h0100a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00806] =  I8a0037ad2845a3fbba9da380a8b8a576['h0100c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00807] =  I8a0037ad2845a3fbba9da380a8b8a576['h0100e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00808] =  I8a0037ad2845a3fbba9da380a8b8a576['h01010] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00809] =  I8a0037ad2845a3fbba9da380a8b8a576['h01012] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0080a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01014] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0080b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01016] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0080c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01018] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0080d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0101a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0080e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0101c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0080f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0101e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00810] =  I8a0037ad2845a3fbba9da380a8b8a576['h01020] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00811] =  I8a0037ad2845a3fbba9da380a8b8a576['h01022] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00812] =  I8a0037ad2845a3fbba9da380a8b8a576['h01024] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00813] =  I8a0037ad2845a3fbba9da380a8b8a576['h01026] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00814] =  I8a0037ad2845a3fbba9da380a8b8a576['h01028] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00815] =  I8a0037ad2845a3fbba9da380a8b8a576['h0102a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00816] =  I8a0037ad2845a3fbba9da380a8b8a576['h0102c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00817] =  I8a0037ad2845a3fbba9da380a8b8a576['h0102e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00818] =  I8a0037ad2845a3fbba9da380a8b8a576['h01030] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00819] =  I8a0037ad2845a3fbba9da380a8b8a576['h01032] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0081a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01034] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0081b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01036] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0081c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01038] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0081d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0103a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0081e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0103c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0081f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0103e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00820] =  I8a0037ad2845a3fbba9da380a8b8a576['h01040] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00821] =  I8a0037ad2845a3fbba9da380a8b8a576['h01042] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00822] =  I8a0037ad2845a3fbba9da380a8b8a576['h01044] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00823] =  I8a0037ad2845a3fbba9da380a8b8a576['h01046] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00824] =  I8a0037ad2845a3fbba9da380a8b8a576['h01048] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00825] =  I8a0037ad2845a3fbba9da380a8b8a576['h0104a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00826] =  I8a0037ad2845a3fbba9da380a8b8a576['h0104c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00827] =  I8a0037ad2845a3fbba9da380a8b8a576['h0104e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00828] =  I8a0037ad2845a3fbba9da380a8b8a576['h01050] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00829] =  I8a0037ad2845a3fbba9da380a8b8a576['h01052] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0082a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01054] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0082b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01056] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0082c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01058] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0082d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0105a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0082e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0105c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0082f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0105e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00830] =  I8a0037ad2845a3fbba9da380a8b8a576['h01060] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00831] =  I8a0037ad2845a3fbba9da380a8b8a576['h01062] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00832] =  I8a0037ad2845a3fbba9da380a8b8a576['h01064] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00833] =  I8a0037ad2845a3fbba9da380a8b8a576['h01066] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00834] =  I8a0037ad2845a3fbba9da380a8b8a576['h01068] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00835] =  I8a0037ad2845a3fbba9da380a8b8a576['h0106a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00836] =  I8a0037ad2845a3fbba9da380a8b8a576['h0106c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00837] =  I8a0037ad2845a3fbba9da380a8b8a576['h0106e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00838] =  I8a0037ad2845a3fbba9da380a8b8a576['h01070] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00839] =  I8a0037ad2845a3fbba9da380a8b8a576['h01072] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0083a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01074] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0083b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01076] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0083c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01078] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0083d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0107a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0083e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0107c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0083f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0107e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00840] =  I8a0037ad2845a3fbba9da380a8b8a576['h01080] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00841] =  I8a0037ad2845a3fbba9da380a8b8a576['h01082] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00842] =  I8a0037ad2845a3fbba9da380a8b8a576['h01084] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00843] =  I8a0037ad2845a3fbba9da380a8b8a576['h01086] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00844] =  I8a0037ad2845a3fbba9da380a8b8a576['h01088] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00845] =  I8a0037ad2845a3fbba9da380a8b8a576['h0108a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00846] =  I8a0037ad2845a3fbba9da380a8b8a576['h0108c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00847] =  I8a0037ad2845a3fbba9da380a8b8a576['h0108e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00848] =  I8a0037ad2845a3fbba9da380a8b8a576['h01090] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00849] =  I8a0037ad2845a3fbba9da380a8b8a576['h01092] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0084a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01094] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0084b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01096] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0084c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01098] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0084d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0109a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0084e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0109c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0084f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0109e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00850] =  I8a0037ad2845a3fbba9da380a8b8a576['h010a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00851] =  I8a0037ad2845a3fbba9da380a8b8a576['h010a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00852] =  I8a0037ad2845a3fbba9da380a8b8a576['h010a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00853] =  I8a0037ad2845a3fbba9da380a8b8a576['h010a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00854] =  I8a0037ad2845a3fbba9da380a8b8a576['h010a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00855] =  I8a0037ad2845a3fbba9da380a8b8a576['h010aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00856] =  I8a0037ad2845a3fbba9da380a8b8a576['h010ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00857] =  I8a0037ad2845a3fbba9da380a8b8a576['h010ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00858] =  I8a0037ad2845a3fbba9da380a8b8a576['h010b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00859] =  I8a0037ad2845a3fbba9da380a8b8a576['h010b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0085a] =  I8a0037ad2845a3fbba9da380a8b8a576['h010b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0085b] =  I8a0037ad2845a3fbba9da380a8b8a576['h010b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0085c] =  I8a0037ad2845a3fbba9da380a8b8a576['h010b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0085d] =  I8a0037ad2845a3fbba9da380a8b8a576['h010ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0085e] =  I8a0037ad2845a3fbba9da380a8b8a576['h010bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0085f] =  I8a0037ad2845a3fbba9da380a8b8a576['h010be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00860] =  I8a0037ad2845a3fbba9da380a8b8a576['h010c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00861] =  I8a0037ad2845a3fbba9da380a8b8a576['h010c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00862] =  I8a0037ad2845a3fbba9da380a8b8a576['h010c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00863] =  I8a0037ad2845a3fbba9da380a8b8a576['h010c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00864] =  I8a0037ad2845a3fbba9da380a8b8a576['h010c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00865] =  I8a0037ad2845a3fbba9da380a8b8a576['h010ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00866] =  I8a0037ad2845a3fbba9da380a8b8a576['h010cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00867] =  I8a0037ad2845a3fbba9da380a8b8a576['h010ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00868] =  I8a0037ad2845a3fbba9da380a8b8a576['h010d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00869] =  I8a0037ad2845a3fbba9da380a8b8a576['h010d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0086a] =  I8a0037ad2845a3fbba9da380a8b8a576['h010d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0086b] =  I8a0037ad2845a3fbba9da380a8b8a576['h010d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0086c] =  I8a0037ad2845a3fbba9da380a8b8a576['h010d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0086d] =  I8a0037ad2845a3fbba9da380a8b8a576['h010da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0086e] =  I8a0037ad2845a3fbba9da380a8b8a576['h010dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0086f] =  I8a0037ad2845a3fbba9da380a8b8a576['h010de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00870] =  I8a0037ad2845a3fbba9da380a8b8a576['h010e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00871] =  I8a0037ad2845a3fbba9da380a8b8a576['h010e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00872] =  I8a0037ad2845a3fbba9da380a8b8a576['h010e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00873] =  I8a0037ad2845a3fbba9da380a8b8a576['h010e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00874] =  I8a0037ad2845a3fbba9da380a8b8a576['h010e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00875] =  I8a0037ad2845a3fbba9da380a8b8a576['h010ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00876] =  I8a0037ad2845a3fbba9da380a8b8a576['h010ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00877] =  I8a0037ad2845a3fbba9da380a8b8a576['h010ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00878] =  I8a0037ad2845a3fbba9da380a8b8a576['h010f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00879] =  I8a0037ad2845a3fbba9da380a8b8a576['h010f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0087a] =  I8a0037ad2845a3fbba9da380a8b8a576['h010f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0087b] =  I8a0037ad2845a3fbba9da380a8b8a576['h010f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0087c] =  I8a0037ad2845a3fbba9da380a8b8a576['h010f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0087d] =  I8a0037ad2845a3fbba9da380a8b8a576['h010fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0087e] =  I8a0037ad2845a3fbba9da380a8b8a576['h010fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0087f] =  I8a0037ad2845a3fbba9da380a8b8a576['h010fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00880] =  I8a0037ad2845a3fbba9da380a8b8a576['h01100] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00881] =  I8a0037ad2845a3fbba9da380a8b8a576['h01102] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00882] =  I8a0037ad2845a3fbba9da380a8b8a576['h01104] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00883] =  I8a0037ad2845a3fbba9da380a8b8a576['h01106] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00884] =  I8a0037ad2845a3fbba9da380a8b8a576['h01108] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00885] =  I8a0037ad2845a3fbba9da380a8b8a576['h0110a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00886] =  I8a0037ad2845a3fbba9da380a8b8a576['h0110c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00887] =  I8a0037ad2845a3fbba9da380a8b8a576['h0110e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00888] =  I8a0037ad2845a3fbba9da380a8b8a576['h01110] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00889] =  I8a0037ad2845a3fbba9da380a8b8a576['h01112] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0088a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01114] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0088b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01116] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0088c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01118] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0088d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0111a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0088e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0111c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0088f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0111e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00890] =  I8a0037ad2845a3fbba9da380a8b8a576['h01120] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00891] =  I8a0037ad2845a3fbba9da380a8b8a576['h01122] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00892] =  I8a0037ad2845a3fbba9da380a8b8a576['h01124] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00893] =  I8a0037ad2845a3fbba9da380a8b8a576['h01126] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00894] =  I8a0037ad2845a3fbba9da380a8b8a576['h01128] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00895] =  I8a0037ad2845a3fbba9da380a8b8a576['h0112a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00896] =  I8a0037ad2845a3fbba9da380a8b8a576['h0112c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00897] =  I8a0037ad2845a3fbba9da380a8b8a576['h0112e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00898] =  I8a0037ad2845a3fbba9da380a8b8a576['h01130] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00899] =  I8a0037ad2845a3fbba9da380a8b8a576['h01132] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0089a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01134] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0089b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01136] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0089c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01138] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0089d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0113a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0089e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0113c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0089f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0113e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01140] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01142] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01144] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01146] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01148] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0114a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0114c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0114e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01150] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01152] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h01154] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h01156] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h01158] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0115a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0115c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008af] =  I8a0037ad2845a3fbba9da380a8b8a576['h0115e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01160] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01162] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01164] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01166] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01168] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0116a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0116c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0116e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01170] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01172] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h01174] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h01176] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h01178] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0117a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008be] =  I8a0037ad2845a3fbba9da380a8b8a576['h0117c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0117e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01180] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01182] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01184] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01186] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01188] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0118a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0118c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0118e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01190] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01192] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h01194] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h01196] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h01198] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0119a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0119c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0119e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h011a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h011a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h011a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h011a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h011a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h011aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h011ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h011ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h011b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h011b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008da] =  I8a0037ad2845a3fbba9da380a8b8a576['h011b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008db] =  I8a0037ad2845a3fbba9da380a8b8a576['h011b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h011b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h011ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008de] =  I8a0037ad2845a3fbba9da380a8b8a576['h011bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008df] =  I8a0037ad2845a3fbba9da380a8b8a576['h011be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h011c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h011c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h011c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h011c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h011c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h011ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h011cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h011ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h011d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h011d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h011d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h011d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h011d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h011da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h011dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h011de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h011e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h011e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h011e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h011e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h011e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h011ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h011ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h011ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h011f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h011f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h011f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h011f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h011f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h011fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h011fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h008ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h011fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00900] =  I8a0037ad2845a3fbba9da380a8b8a576['h01200] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00901] =  I8a0037ad2845a3fbba9da380a8b8a576['h01202] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00902] =  I8a0037ad2845a3fbba9da380a8b8a576['h01204] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00903] =  I8a0037ad2845a3fbba9da380a8b8a576['h01206] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00904] =  I8a0037ad2845a3fbba9da380a8b8a576['h01208] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00905] =  I8a0037ad2845a3fbba9da380a8b8a576['h0120a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00906] =  I8a0037ad2845a3fbba9da380a8b8a576['h0120c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00907] =  I8a0037ad2845a3fbba9da380a8b8a576['h0120e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00908] =  I8a0037ad2845a3fbba9da380a8b8a576['h01210] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00909] =  I8a0037ad2845a3fbba9da380a8b8a576['h01212] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0090a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01214] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0090b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01216] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0090c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01218] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0090d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0121a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0090e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0121c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0090f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0121e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00910] =  I8a0037ad2845a3fbba9da380a8b8a576['h01220] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00911] =  I8a0037ad2845a3fbba9da380a8b8a576['h01222] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00912] =  I8a0037ad2845a3fbba9da380a8b8a576['h01224] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00913] =  I8a0037ad2845a3fbba9da380a8b8a576['h01226] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00914] =  I8a0037ad2845a3fbba9da380a8b8a576['h01228] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00915] =  I8a0037ad2845a3fbba9da380a8b8a576['h0122a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00916] =  I8a0037ad2845a3fbba9da380a8b8a576['h0122c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00917] =  I8a0037ad2845a3fbba9da380a8b8a576['h0122e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00918] =  I8a0037ad2845a3fbba9da380a8b8a576['h01230] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00919] =  I8a0037ad2845a3fbba9da380a8b8a576['h01232] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0091a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01234] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0091b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01236] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0091c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01238] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0091d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0123a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0091e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0123c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0091f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0123e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00920] =  I8a0037ad2845a3fbba9da380a8b8a576['h01240] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00921] =  I8a0037ad2845a3fbba9da380a8b8a576['h01242] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00922] =  I8a0037ad2845a3fbba9da380a8b8a576['h01244] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00923] =  I8a0037ad2845a3fbba9da380a8b8a576['h01246] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00924] =  I8a0037ad2845a3fbba9da380a8b8a576['h01248] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00925] =  I8a0037ad2845a3fbba9da380a8b8a576['h0124a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00926] =  I8a0037ad2845a3fbba9da380a8b8a576['h0124c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00927] =  I8a0037ad2845a3fbba9da380a8b8a576['h0124e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00928] =  I8a0037ad2845a3fbba9da380a8b8a576['h01250] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00929] =  I8a0037ad2845a3fbba9da380a8b8a576['h01252] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0092a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01254] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0092b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01256] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0092c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01258] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0092d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0125a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0092e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0125c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0092f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0125e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00930] =  I8a0037ad2845a3fbba9da380a8b8a576['h01260] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00931] =  I8a0037ad2845a3fbba9da380a8b8a576['h01262] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00932] =  I8a0037ad2845a3fbba9da380a8b8a576['h01264] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00933] =  I8a0037ad2845a3fbba9da380a8b8a576['h01266] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00934] =  I8a0037ad2845a3fbba9da380a8b8a576['h01268] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00935] =  I8a0037ad2845a3fbba9da380a8b8a576['h0126a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00936] =  I8a0037ad2845a3fbba9da380a8b8a576['h0126c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00937] =  I8a0037ad2845a3fbba9da380a8b8a576['h0126e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00938] =  I8a0037ad2845a3fbba9da380a8b8a576['h01270] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00939] =  I8a0037ad2845a3fbba9da380a8b8a576['h01272] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0093a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01274] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0093b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01276] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0093c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01278] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0093d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0127a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0093e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0127c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0093f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0127e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00940] =  I8a0037ad2845a3fbba9da380a8b8a576['h01280] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00941] =  I8a0037ad2845a3fbba9da380a8b8a576['h01282] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00942] =  I8a0037ad2845a3fbba9da380a8b8a576['h01284] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00943] =  I8a0037ad2845a3fbba9da380a8b8a576['h01286] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00944] =  I8a0037ad2845a3fbba9da380a8b8a576['h01288] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00945] =  I8a0037ad2845a3fbba9da380a8b8a576['h0128a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00946] =  I8a0037ad2845a3fbba9da380a8b8a576['h0128c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00947] =  I8a0037ad2845a3fbba9da380a8b8a576['h0128e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00948] =  I8a0037ad2845a3fbba9da380a8b8a576['h01290] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00949] =  I8a0037ad2845a3fbba9da380a8b8a576['h01292] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0094a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01294] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0094b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01296] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0094c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01298] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0094d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0129a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0094e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0129c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0094f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0129e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00950] =  I8a0037ad2845a3fbba9da380a8b8a576['h012a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00951] =  I8a0037ad2845a3fbba9da380a8b8a576['h012a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00952] =  I8a0037ad2845a3fbba9da380a8b8a576['h012a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00953] =  I8a0037ad2845a3fbba9da380a8b8a576['h012a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00954] =  I8a0037ad2845a3fbba9da380a8b8a576['h012a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00955] =  I8a0037ad2845a3fbba9da380a8b8a576['h012aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00956] =  I8a0037ad2845a3fbba9da380a8b8a576['h012ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00957] =  I8a0037ad2845a3fbba9da380a8b8a576['h012ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00958] =  I8a0037ad2845a3fbba9da380a8b8a576['h012b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00959] =  I8a0037ad2845a3fbba9da380a8b8a576['h012b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0095a] =  I8a0037ad2845a3fbba9da380a8b8a576['h012b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0095b] =  I8a0037ad2845a3fbba9da380a8b8a576['h012b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0095c] =  I8a0037ad2845a3fbba9da380a8b8a576['h012b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0095d] =  I8a0037ad2845a3fbba9da380a8b8a576['h012ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0095e] =  I8a0037ad2845a3fbba9da380a8b8a576['h012bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0095f] =  I8a0037ad2845a3fbba9da380a8b8a576['h012be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00960] =  I8a0037ad2845a3fbba9da380a8b8a576['h012c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00961] =  I8a0037ad2845a3fbba9da380a8b8a576['h012c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00962] =  I8a0037ad2845a3fbba9da380a8b8a576['h012c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00963] =  I8a0037ad2845a3fbba9da380a8b8a576['h012c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00964] =  I8a0037ad2845a3fbba9da380a8b8a576['h012c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00965] =  I8a0037ad2845a3fbba9da380a8b8a576['h012ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00966] =  I8a0037ad2845a3fbba9da380a8b8a576['h012cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00967] =  I8a0037ad2845a3fbba9da380a8b8a576['h012ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00968] =  I8a0037ad2845a3fbba9da380a8b8a576['h012d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00969] =  I8a0037ad2845a3fbba9da380a8b8a576['h012d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0096a] =  I8a0037ad2845a3fbba9da380a8b8a576['h012d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0096b] =  I8a0037ad2845a3fbba9da380a8b8a576['h012d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0096c] =  I8a0037ad2845a3fbba9da380a8b8a576['h012d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0096d] =  I8a0037ad2845a3fbba9da380a8b8a576['h012da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0096e] =  I8a0037ad2845a3fbba9da380a8b8a576['h012dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0096f] =  I8a0037ad2845a3fbba9da380a8b8a576['h012de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00970] =  I8a0037ad2845a3fbba9da380a8b8a576['h012e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00971] =  I8a0037ad2845a3fbba9da380a8b8a576['h012e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00972] =  I8a0037ad2845a3fbba9da380a8b8a576['h012e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00973] =  I8a0037ad2845a3fbba9da380a8b8a576['h012e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00974] =  I8a0037ad2845a3fbba9da380a8b8a576['h012e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00975] =  I8a0037ad2845a3fbba9da380a8b8a576['h012ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00976] =  I8a0037ad2845a3fbba9da380a8b8a576['h012ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00977] =  I8a0037ad2845a3fbba9da380a8b8a576['h012ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00978] =  I8a0037ad2845a3fbba9da380a8b8a576['h012f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00979] =  I8a0037ad2845a3fbba9da380a8b8a576['h012f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0097a] =  I8a0037ad2845a3fbba9da380a8b8a576['h012f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0097b] =  I8a0037ad2845a3fbba9da380a8b8a576['h012f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0097c] =  I8a0037ad2845a3fbba9da380a8b8a576['h012f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0097d] =  I8a0037ad2845a3fbba9da380a8b8a576['h012fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0097e] =  I8a0037ad2845a3fbba9da380a8b8a576['h012fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0097f] =  I8a0037ad2845a3fbba9da380a8b8a576['h012fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00980] =  I8a0037ad2845a3fbba9da380a8b8a576['h01300] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00981] =  I8a0037ad2845a3fbba9da380a8b8a576['h01302] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00982] =  I8a0037ad2845a3fbba9da380a8b8a576['h01304] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00983] =  I8a0037ad2845a3fbba9da380a8b8a576['h01306] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00984] =  I8a0037ad2845a3fbba9da380a8b8a576['h01308] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00985] =  I8a0037ad2845a3fbba9da380a8b8a576['h0130a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00986] =  I8a0037ad2845a3fbba9da380a8b8a576['h0130c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00987] =  I8a0037ad2845a3fbba9da380a8b8a576['h0130e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00988] =  I8a0037ad2845a3fbba9da380a8b8a576['h01310] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00989] =  I8a0037ad2845a3fbba9da380a8b8a576['h01312] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0098a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01314] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0098b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01316] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0098c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01318] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0098d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0131a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0098e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0131c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0098f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0131e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00990] =  I8a0037ad2845a3fbba9da380a8b8a576['h01320] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00991] =  I8a0037ad2845a3fbba9da380a8b8a576['h01322] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00992] =  I8a0037ad2845a3fbba9da380a8b8a576['h01324] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00993] =  I8a0037ad2845a3fbba9da380a8b8a576['h01326] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00994] =  I8a0037ad2845a3fbba9da380a8b8a576['h01328] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00995] =  I8a0037ad2845a3fbba9da380a8b8a576['h0132a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00996] =  I8a0037ad2845a3fbba9da380a8b8a576['h0132c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00997] =  I8a0037ad2845a3fbba9da380a8b8a576['h0132e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00998] =  I8a0037ad2845a3fbba9da380a8b8a576['h01330] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00999] =  I8a0037ad2845a3fbba9da380a8b8a576['h01332] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0099a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01334] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0099b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01336] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0099c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01338] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0099d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0133a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0099e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0133c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0099f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0133e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01340] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01342] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01344] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01346] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01348] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0134a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0134c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0134e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01350] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01352] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h01354] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h01356] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h01358] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0135a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0135c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009af] =  I8a0037ad2845a3fbba9da380a8b8a576['h0135e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01360] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01362] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01364] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01366] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01368] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0136a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0136c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0136e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01370] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01372] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h01374] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h01376] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h01378] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0137a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009be] =  I8a0037ad2845a3fbba9da380a8b8a576['h0137c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0137e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01380] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01382] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01384] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01386] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01388] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0138a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0138c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0138e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01390] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01392] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h01394] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h01396] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h01398] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0139a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0139c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0139e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h013a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h013a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h013a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h013a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h013a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h013aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h013ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h013ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h013b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h013b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009da] =  I8a0037ad2845a3fbba9da380a8b8a576['h013b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009db] =  I8a0037ad2845a3fbba9da380a8b8a576['h013b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h013b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h013ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009de] =  I8a0037ad2845a3fbba9da380a8b8a576['h013bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009df] =  I8a0037ad2845a3fbba9da380a8b8a576['h013be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h013c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h013c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h013c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h013c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h013c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h013ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h013cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h013ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h013d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h013d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h013d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h013d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h013d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h013da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h013dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h013de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h013e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h013e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h013e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h013e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h013e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h013ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h013ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h013ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h013f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h013f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h013f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h013f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h013f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h013fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h013fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h009ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h013fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a00] =  I8a0037ad2845a3fbba9da380a8b8a576['h01400] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a01] =  I8a0037ad2845a3fbba9da380a8b8a576['h01402] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a02] =  I8a0037ad2845a3fbba9da380a8b8a576['h01404] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a03] =  I8a0037ad2845a3fbba9da380a8b8a576['h01406] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a04] =  I8a0037ad2845a3fbba9da380a8b8a576['h01408] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a05] =  I8a0037ad2845a3fbba9da380a8b8a576['h0140a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a06] =  I8a0037ad2845a3fbba9da380a8b8a576['h0140c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a07] =  I8a0037ad2845a3fbba9da380a8b8a576['h0140e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a08] =  I8a0037ad2845a3fbba9da380a8b8a576['h01410] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a09] =  I8a0037ad2845a3fbba9da380a8b8a576['h01412] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a0a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01414] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a0b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01416] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a0c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01418] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a0d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0141a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a0e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0141c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a0f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0141e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a10] =  I8a0037ad2845a3fbba9da380a8b8a576['h01420] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a11] =  I8a0037ad2845a3fbba9da380a8b8a576['h01422] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a12] =  I8a0037ad2845a3fbba9da380a8b8a576['h01424] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a13] =  I8a0037ad2845a3fbba9da380a8b8a576['h01426] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a14] =  I8a0037ad2845a3fbba9da380a8b8a576['h01428] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a15] =  I8a0037ad2845a3fbba9da380a8b8a576['h0142a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a16] =  I8a0037ad2845a3fbba9da380a8b8a576['h0142c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a17] =  I8a0037ad2845a3fbba9da380a8b8a576['h0142e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a18] =  I8a0037ad2845a3fbba9da380a8b8a576['h01430] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a19] =  I8a0037ad2845a3fbba9da380a8b8a576['h01432] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a1a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01434] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a1b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01436] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a1c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01438] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a1d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0143a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a1e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0143c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a1f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0143e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a20] =  I8a0037ad2845a3fbba9da380a8b8a576['h01440] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a21] =  I8a0037ad2845a3fbba9da380a8b8a576['h01442] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a22] =  I8a0037ad2845a3fbba9da380a8b8a576['h01444] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a23] =  I8a0037ad2845a3fbba9da380a8b8a576['h01446] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a24] =  I8a0037ad2845a3fbba9da380a8b8a576['h01448] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a25] =  I8a0037ad2845a3fbba9da380a8b8a576['h0144a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a26] =  I8a0037ad2845a3fbba9da380a8b8a576['h0144c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a27] =  I8a0037ad2845a3fbba9da380a8b8a576['h0144e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a28] =  I8a0037ad2845a3fbba9da380a8b8a576['h01450] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a29] =  I8a0037ad2845a3fbba9da380a8b8a576['h01452] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a2a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01454] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a2b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01456] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a2c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01458] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a2d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0145a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a2e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0145c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a2f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0145e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a30] =  I8a0037ad2845a3fbba9da380a8b8a576['h01460] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a31] =  I8a0037ad2845a3fbba9da380a8b8a576['h01462] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a32] =  I8a0037ad2845a3fbba9da380a8b8a576['h01464] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a33] =  I8a0037ad2845a3fbba9da380a8b8a576['h01466] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a34] =  I8a0037ad2845a3fbba9da380a8b8a576['h01468] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a35] =  I8a0037ad2845a3fbba9da380a8b8a576['h0146a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a36] =  I8a0037ad2845a3fbba9da380a8b8a576['h0146c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a37] =  I8a0037ad2845a3fbba9da380a8b8a576['h0146e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a38] =  I8a0037ad2845a3fbba9da380a8b8a576['h01470] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a39] =  I8a0037ad2845a3fbba9da380a8b8a576['h01472] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a3a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01474] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a3b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01476] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a3c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01478] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a3d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0147a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a3e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0147c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a3f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0147e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a40] =  I8a0037ad2845a3fbba9da380a8b8a576['h01480] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a41] =  I8a0037ad2845a3fbba9da380a8b8a576['h01482] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a42] =  I8a0037ad2845a3fbba9da380a8b8a576['h01484] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a43] =  I8a0037ad2845a3fbba9da380a8b8a576['h01486] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a44] =  I8a0037ad2845a3fbba9da380a8b8a576['h01488] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a45] =  I8a0037ad2845a3fbba9da380a8b8a576['h0148a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a46] =  I8a0037ad2845a3fbba9da380a8b8a576['h0148c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a47] =  I8a0037ad2845a3fbba9da380a8b8a576['h0148e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a48] =  I8a0037ad2845a3fbba9da380a8b8a576['h01490] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a49] =  I8a0037ad2845a3fbba9da380a8b8a576['h01492] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a4a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01494] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a4b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01496] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a4c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01498] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a4d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0149a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a4e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0149c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a4f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0149e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a50] =  I8a0037ad2845a3fbba9da380a8b8a576['h014a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a51] =  I8a0037ad2845a3fbba9da380a8b8a576['h014a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a52] =  I8a0037ad2845a3fbba9da380a8b8a576['h014a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a53] =  I8a0037ad2845a3fbba9da380a8b8a576['h014a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a54] =  I8a0037ad2845a3fbba9da380a8b8a576['h014a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a55] =  I8a0037ad2845a3fbba9da380a8b8a576['h014aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a56] =  I8a0037ad2845a3fbba9da380a8b8a576['h014ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a57] =  I8a0037ad2845a3fbba9da380a8b8a576['h014ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a58] =  I8a0037ad2845a3fbba9da380a8b8a576['h014b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a59] =  I8a0037ad2845a3fbba9da380a8b8a576['h014b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a5a] =  I8a0037ad2845a3fbba9da380a8b8a576['h014b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a5b] =  I8a0037ad2845a3fbba9da380a8b8a576['h014b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a5c] =  I8a0037ad2845a3fbba9da380a8b8a576['h014b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a5d] =  I8a0037ad2845a3fbba9da380a8b8a576['h014ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a5e] =  I8a0037ad2845a3fbba9da380a8b8a576['h014bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a5f] =  I8a0037ad2845a3fbba9da380a8b8a576['h014be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a60] =  I8a0037ad2845a3fbba9da380a8b8a576['h014c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a61] =  I8a0037ad2845a3fbba9da380a8b8a576['h014c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a62] =  I8a0037ad2845a3fbba9da380a8b8a576['h014c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a63] =  I8a0037ad2845a3fbba9da380a8b8a576['h014c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a64] =  I8a0037ad2845a3fbba9da380a8b8a576['h014c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a65] =  I8a0037ad2845a3fbba9da380a8b8a576['h014ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a66] =  I8a0037ad2845a3fbba9da380a8b8a576['h014cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a67] =  I8a0037ad2845a3fbba9da380a8b8a576['h014ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a68] =  I8a0037ad2845a3fbba9da380a8b8a576['h014d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a69] =  I8a0037ad2845a3fbba9da380a8b8a576['h014d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a6a] =  I8a0037ad2845a3fbba9da380a8b8a576['h014d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a6b] =  I8a0037ad2845a3fbba9da380a8b8a576['h014d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a6c] =  I8a0037ad2845a3fbba9da380a8b8a576['h014d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a6d] =  I8a0037ad2845a3fbba9da380a8b8a576['h014da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a6e] =  I8a0037ad2845a3fbba9da380a8b8a576['h014dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a6f] =  I8a0037ad2845a3fbba9da380a8b8a576['h014de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a70] =  I8a0037ad2845a3fbba9da380a8b8a576['h014e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a71] =  I8a0037ad2845a3fbba9da380a8b8a576['h014e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a72] =  I8a0037ad2845a3fbba9da380a8b8a576['h014e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a73] =  I8a0037ad2845a3fbba9da380a8b8a576['h014e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a74] =  I8a0037ad2845a3fbba9da380a8b8a576['h014e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a75] =  I8a0037ad2845a3fbba9da380a8b8a576['h014ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a76] =  I8a0037ad2845a3fbba9da380a8b8a576['h014ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a77] =  I8a0037ad2845a3fbba9da380a8b8a576['h014ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a78] =  I8a0037ad2845a3fbba9da380a8b8a576['h014f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a79] =  I8a0037ad2845a3fbba9da380a8b8a576['h014f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a7a] =  I8a0037ad2845a3fbba9da380a8b8a576['h014f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a7b] =  I8a0037ad2845a3fbba9da380a8b8a576['h014f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a7c] =  I8a0037ad2845a3fbba9da380a8b8a576['h014f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a7d] =  I8a0037ad2845a3fbba9da380a8b8a576['h014fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a7e] =  I8a0037ad2845a3fbba9da380a8b8a576['h014fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a7f] =  I8a0037ad2845a3fbba9da380a8b8a576['h014fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a80] =  I8a0037ad2845a3fbba9da380a8b8a576['h01500] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a81] =  I8a0037ad2845a3fbba9da380a8b8a576['h01502] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a82] =  I8a0037ad2845a3fbba9da380a8b8a576['h01504] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a83] =  I8a0037ad2845a3fbba9da380a8b8a576['h01506] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a84] =  I8a0037ad2845a3fbba9da380a8b8a576['h01508] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a85] =  I8a0037ad2845a3fbba9da380a8b8a576['h0150a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a86] =  I8a0037ad2845a3fbba9da380a8b8a576['h0150c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a87] =  I8a0037ad2845a3fbba9da380a8b8a576['h0150e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a88] =  I8a0037ad2845a3fbba9da380a8b8a576['h01510] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a89] =  I8a0037ad2845a3fbba9da380a8b8a576['h01512] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a8a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01514] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a8b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01516] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a8c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01518] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a8d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0151a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a8e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0151c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a8f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0151e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a90] =  I8a0037ad2845a3fbba9da380a8b8a576['h01520] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a91] =  I8a0037ad2845a3fbba9da380a8b8a576['h01522] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a92] =  I8a0037ad2845a3fbba9da380a8b8a576['h01524] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a93] =  I8a0037ad2845a3fbba9da380a8b8a576['h01526] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a94] =  I8a0037ad2845a3fbba9da380a8b8a576['h01528] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a95] =  I8a0037ad2845a3fbba9da380a8b8a576['h0152a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a96] =  I8a0037ad2845a3fbba9da380a8b8a576['h0152c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a97] =  I8a0037ad2845a3fbba9da380a8b8a576['h0152e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a98] =  I8a0037ad2845a3fbba9da380a8b8a576['h01530] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a99] =  I8a0037ad2845a3fbba9da380a8b8a576['h01532] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a9a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01534] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a9b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01536] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a9c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01538] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a9d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0153a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a9e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0153c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00a9f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0153e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00aa0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01540] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00aa1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01542] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00aa2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01544] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00aa3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01546] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00aa4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01548] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00aa5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0154a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00aa6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0154c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00aa7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0154e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00aa8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01550] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00aa9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01552] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00aaa] =  I8a0037ad2845a3fbba9da380a8b8a576['h01554] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00aab] =  I8a0037ad2845a3fbba9da380a8b8a576['h01556] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00aac] =  I8a0037ad2845a3fbba9da380a8b8a576['h01558] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00aad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0155a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00aae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0155c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00aaf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0155e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ab0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01560] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ab1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01562] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ab2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01564] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ab3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01566] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ab4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01568] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ab5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0156a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ab6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0156c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ab7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0156e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ab8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01570] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ab9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01572] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00aba] =  I8a0037ad2845a3fbba9da380a8b8a576['h01574] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00abb] =  I8a0037ad2845a3fbba9da380a8b8a576['h01576] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00abc] =  I8a0037ad2845a3fbba9da380a8b8a576['h01578] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00abd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0157a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00abe] =  I8a0037ad2845a3fbba9da380a8b8a576['h0157c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00abf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0157e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ac0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01580] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ac1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01582] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ac2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01584] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ac3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01586] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ac4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01588] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ac5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0158a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ac6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0158c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ac7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0158e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ac8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01590] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ac9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01592] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00aca] =  I8a0037ad2845a3fbba9da380a8b8a576['h01594] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00acb] =  I8a0037ad2845a3fbba9da380a8b8a576['h01596] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00acc] =  I8a0037ad2845a3fbba9da380a8b8a576['h01598] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00acd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0159a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ace] =  I8a0037ad2845a3fbba9da380a8b8a576['h0159c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00acf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0159e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ad0] =  I8a0037ad2845a3fbba9da380a8b8a576['h015a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ad1] =  I8a0037ad2845a3fbba9da380a8b8a576['h015a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ad2] =  I8a0037ad2845a3fbba9da380a8b8a576['h015a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ad3] =  I8a0037ad2845a3fbba9da380a8b8a576['h015a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ad4] =  I8a0037ad2845a3fbba9da380a8b8a576['h015a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ad5] =  I8a0037ad2845a3fbba9da380a8b8a576['h015aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ad6] =  I8a0037ad2845a3fbba9da380a8b8a576['h015ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ad7] =  I8a0037ad2845a3fbba9da380a8b8a576['h015ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ad8] =  I8a0037ad2845a3fbba9da380a8b8a576['h015b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ad9] =  I8a0037ad2845a3fbba9da380a8b8a576['h015b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ada] =  I8a0037ad2845a3fbba9da380a8b8a576['h015b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00adb] =  I8a0037ad2845a3fbba9da380a8b8a576['h015b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00adc] =  I8a0037ad2845a3fbba9da380a8b8a576['h015b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00add] =  I8a0037ad2845a3fbba9da380a8b8a576['h015ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ade] =  I8a0037ad2845a3fbba9da380a8b8a576['h015bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00adf] =  I8a0037ad2845a3fbba9da380a8b8a576['h015be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ae0] =  I8a0037ad2845a3fbba9da380a8b8a576['h015c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ae1] =  I8a0037ad2845a3fbba9da380a8b8a576['h015c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ae2] =  I8a0037ad2845a3fbba9da380a8b8a576['h015c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ae3] =  I8a0037ad2845a3fbba9da380a8b8a576['h015c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ae4] =  I8a0037ad2845a3fbba9da380a8b8a576['h015c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ae5] =  I8a0037ad2845a3fbba9da380a8b8a576['h015ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ae6] =  I8a0037ad2845a3fbba9da380a8b8a576['h015cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ae7] =  I8a0037ad2845a3fbba9da380a8b8a576['h015ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ae8] =  I8a0037ad2845a3fbba9da380a8b8a576['h015d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ae9] =  I8a0037ad2845a3fbba9da380a8b8a576['h015d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00aea] =  I8a0037ad2845a3fbba9da380a8b8a576['h015d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00aeb] =  I8a0037ad2845a3fbba9da380a8b8a576['h015d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00aec] =  I8a0037ad2845a3fbba9da380a8b8a576['h015d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00aed] =  I8a0037ad2845a3fbba9da380a8b8a576['h015da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00aee] =  I8a0037ad2845a3fbba9da380a8b8a576['h015dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00aef] =  I8a0037ad2845a3fbba9da380a8b8a576['h015de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00af0] =  I8a0037ad2845a3fbba9da380a8b8a576['h015e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00af1] =  I8a0037ad2845a3fbba9da380a8b8a576['h015e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00af2] =  I8a0037ad2845a3fbba9da380a8b8a576['h015e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00af3] =  I8a0037ad2845a3fbba9da380a8b8a576['h015e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00af4] =  I8a0037ad2845a3fbba9da380a8b8a576['h015e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00af5] =  I8a0037ad2845a3fbba9da380a8b8a576['h015ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00af6] =  I8a0037ad2845a3fbba9da380a8b8a576['h015ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00af7] =  I8a0037ad2845a3fbba9da380a8b8a576['h015ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00af8] =  I8a0037ad2845a3fbba9da380a8b8a576['h015f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00af9] =  I8a0037ad2845a3fbba9da380a8b8a576['h015f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00afa] =  I8a0037ad2845a3fbba9da380a8b8a576['h015f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00afb] =  I8a0037ad2845a3fbba9da380a8b8a576['h015f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00afc] =  I8a0037ad2845a3fbba9da380a8b8a576['h015f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00afd] =  I8a0037ad2845a3fbba9da380a8b8a576['h015fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00afe] =  I8a0037ad2845a3fbba9da380a8b8a576['h015fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00aff] =  I8a0037ad2845a3fbba9da380a8b8a576['h015fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b00] =  I8a0037ad2845a3fbba9da380a8b8a576['h01600] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b01] =  I8a0037ad2845a3fbba9da380a8b8a576['h01602] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b02] =  I8a0037ad2845a3fbba9da380a8b8a576['h01604] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b03] =  I8a0037ad2845a3fbba9da380a8b8a576['h01606] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b04] =  I8a0037ad2845a3fbba9da380a8b8a576['h01608] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b05] =  I8a0037ad2845a3fbba9da380a8b8a576['h0160a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b06] =  I8a0037ad2845a3fbba9da380a8b8a576['h0160c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b07] =  I8a0037ad2845a3fbba9da380a8b8a576['h0160e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b08] =  I8a0037ad2845a3fbba9da380a8b8a576['h01610] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b09] =  I8a0037ad2845a3fbba9da380a8b8a576['h01612] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b0a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01614] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b0b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01616] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b0c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01618] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b0d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0161a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b0e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0161c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b0f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0161e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b10] =  I8a0037ad2845a3fbba9da380a8b8a576['h01620] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b11] =  I8a0037ad2845a3fbba9da380a8b8a576['h01622] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b12] =  I8a0037ad2845a3fbba9da380a8b8a576['h01624] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b13] =  I8a0037ad2845a3fbba9da380a8b8a576['h01626] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b14] =  I8a0037ad2845a3fbba9da380a8b8a576['h01628] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b15] =  I8a0037ad2845a3fbba9da380a8b8a576['h0162a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b16] =  I8a0037ad2845a3fbba9da380a8b8a576['h0162c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b17] =  I8a0037ad2845a3fbba9da380a8b8a576['h0162e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b18] =  I8a0037ad2845a3fbba9da380a8b8a576['h01630] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b19] =  I8a0037ad2845a3fbba9da380a8b8a576['h01632] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b1a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01634] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b1b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01636] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b1c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01638] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b1d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0163a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b1e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0163c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b1f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0163e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b20] =  I8a0037ad2845a3fbba9da380a8b8a576['h01640] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b21] =  I8a0037ad2845a3fbba9da380a8b8a576['h01642] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b22] =  I8a0037ad2845a3fbba9da380a8b8a576['h01644] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b23] =  I8a0037ad2845a3fbba9da380a8b8a576['h01646] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b24] =  I8a0037ad2845a3fbba9da380a8b8a576['h01648] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b25] =  I8a0037ad2845a3fbba9da380a8b8a576['h0164a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b26] =  I8a0037ad2845a3fbba9da380a8b8a576['h0164c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b27] =  I8a0037ad2845a3fbba9da380a8b8a576['h0164e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b28] =  I8a0037ad2845a3fbba9da380a8b8a576['h01650] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b29] =  I8a0037ad2845a3fbba9da380a8b8a576['h01652] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b2a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01654] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b2b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01656] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b2c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01658] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b2d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0165a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b2e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0165c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b2f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0165e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b30] =  I8a0037ad2845a3fbba9da380a8b8a576['h01660] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b31] =  I8a0037ad2845a3fbba9da380a8b8a576['h01662] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b32] =  I8a0037ad2845a3fbba9da380a8b8a576['h01664] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b33] =  I8a0037ad2845a3fbba9da380a8b8a576['h01666] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b34] =  I8a0037ad2845a3fbba9da380a8b8a576['h01668] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b35] =  I8a0037ad2845a3fbba9da380a8b8a576['h0166a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b36] =  I8a0037ad2845a3fbba9da380a8b8a576['h0166c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b37] =  I8a0037ad2845a3fbba9da380a8b8a576['h0166e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b38] =  I8a0037ad2845a3fbba9da380a8b8a576['h01670] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b39] =  I8a0037ad2845a3fbba9da380a8b8a576['h01672] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b3a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01674] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b3b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01676] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b3c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01678] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b3d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0167a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b3e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0167c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b3f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0167e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b40] =  I8a0037ad2845a3fbba9da380a8b8a576['h01680] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b41] =  I8a0037ad2845a3fbba9da380a8b8a576['h01682] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b42] =  I8a0037ad2845a3fbba9da380a8b8a576['h01684] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b43] =  I8a0037ad2845a3fbba9da380a8b8a576['h01686] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b44] =  I8a0037ad2845a3fbba9da380a8b8a576['h01688] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b45] =  I8a0037ad2845a3fbba9da380a8b8a576['h0168a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b46] =  I8a0037ad2845a3fbba9da380a8b8a576['h0168c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b47] =  I8a0037ad2845a3fbba9da380a8b8a576['h0168e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b48] =  I8a0037ad2845a3fbba9da380a8b8a576['h01690] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b49] =  I8a0037ad2845a3fbba9da380a8b8a576['h01692] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b4a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01694] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b4b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01696] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b4c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01698] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b4d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0169a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b4e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0169c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b4f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0169e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b50] =  I8a0037ad2845a3fbba9da380a8b8a576['h016a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b51] =  I8a0037ad2845a3fbba9da380a8b8a576['h016a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b52] =  I8a0037ad2845a3fbba9da380a8b8a576['h016a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b53] =  I8a0037ad2845a3fbba9da380a8b8a576['h016a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b54] =  I8a0037ad2845a3fbba9da380a8b8a576['h016a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b55] =  I8a0037ad2845a3fbba9da380a8b8a576['h016aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b56] =  I8a0037ad2845a3fbba9da380a8b8a576['h016ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b57] =  I8a0037ad2845a3fbba9da380a8b8a576['h016ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b58] =  I8a0037ad2845a3fbba9da380a8b8a576['h016b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b59] =  I8a0037ad2845a3fbba9da380a8b8a576['h016b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b5a] =  I8a0037ad2845a3fbba9da380a8b8a576['h016b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b5b] =  I8a0037ad2845a3fbba9da380a8b8a576['h016b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b5c] =  I8a0037ad2845a3fbba9da380a8b8a576['h016b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b5d] =  I8a0037ad2845a3fbba9da380a8b8a576['h016ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b5e] =  I8a0037ad2845a3fbba9da380a8b8a576['h016bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b5f] =  I8a0037ad2845a3fbba9da380a8b8a576['h016be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b60] =  I8a0037ad2845a3fbba9da380a8b8a576['h016c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b61] =  I8a0037ad2845a3fbba9da380a8b8a576['h016c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b62] =  I8a0037ad2845a3fbba9da380a8b8a576['h016c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b63] =  I8a0037ad2845a3fbba9da380a8b8a576['h016c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b64] =  I8a0037ad2845a3fbba9da380a8b8a576['h016c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b65] =  I8a0037ad2845a3fbba9da380a8b8a576['h016ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b66] =  I8a0037ad2845a3fbba9da380a8b8a576['h016cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b67] =  I8a0037ad2845a3fbba9da380a8b8a576['h016ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b68] =  I8a0037ad2845a3fbba9da380a8b8a576['h016d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b69] =  I8a0037ad2845a3fbba9da380a8b8a576['h016d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b6a] =  I8a0037ad2845a3fbba9da380a8b8a576['h016d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b6b] =  I8a0037ad2845a3fbba9da380a8b8a576['h016d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b6c] =  I8a0037ad2845a3fbba9da380a8b8a576['h016d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b6d] =  I8a0037ad2845a3fbba9da380a8b8a576['h016da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b6e] =  I8a0037ad2845a3fbba9da380a8b8a576['h016dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b6f] =  I8a0037ad2845a3fbba9da380a8b8a576['h016de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b70] =  I8a0037ad2845a3fbba9da380a8b8a576['h016e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b71] =  I8a0037ad2845a3fbba9da380a8b8a576['h016e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b72] =  I8a0037ad2845a3fbba9da380a8b8a576['h016e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b73] =  I8a0037ad2845a3fbba9da380a8b8a576['h016e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b74] =  I8a0037ad2845a3fbba9da380a8b8a576['h016e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b75] =  I8a0037ad2845a3fbba9da380a8b8a576['h016ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b76] =  I8a0037ad2845a3fbba9da380a8b8a576['h016ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b77] =  I8a0037ad2845a3fbba9da380a8b8a576['h016ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b78] =  I8a0037ad2845a3fbba9da380a8b8a576['h016f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b79] =  I8a0037ad2845a3fbba9da380a8b8a576['h016f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b7a] =  I8a0037ad2845a3fbba9da380a8b8a576['h016f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b7b] =  I8a0037ad2845a3fbba9da380a8b8a576['h016f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b7c] =  I8a0037ad2845a3fbba9da380a8b8a576['h016f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b7d] =  I8a0037ad2845a3fbba9da380a8b8a576['h016fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b7e] =  I8a0037ad2845a3fbba9da380a8b8a576['h016fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b7f] =  I8a0037ad2845a3fbba9da380a8b8a576['h016fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b80] =  I8a0037ad2845a3fbba9da380a8b8a576['h01700] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b81] =  I8a0037ad2845a3fbba9da380a8b8a576['h01702] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b82] =  I8a0037ad2845a3fbba9da380a8b8a576['h01704] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b83] =  I8a0037ad2845a3fbba9da380a8b8a576['h01706] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b84] =  I8a0037ad2845a3fbba9da380a8b8a576['h01708] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b85] =  I8a0037ad2845a3fbba9da380a8b8a576['h0170a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b86] =  I8a0037ad2845a3fbba9da380a8b8a576['h0170c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b87] =  I8a0037ad2845a3fbba9da380a8b8a576['h0170e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b88] =  I8a0037ad2845a3fbba9da380a8b8a576['h01710] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b89] =  I8a0037ad2845a3fbba9da380a8b8a576['h01712] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b8a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01714] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b8b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01716] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b8c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01718] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b8d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0171a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b8e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0171c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b8f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0171e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b90] =  I8a0037ad2845a3fbba9da380a8b8a576['h01720] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b91] =  I8a0037ad2845a3fbba9da380a8b8a576['h01722] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b92] =  I8a0037ad2845a3fbba9da380a8b8a576['h01724] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b93] =  I8a0037ad2845a3fbba9da380a8b8a576['h01726] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b94] =  I8a0037ad2845a3fbba9da380a8b8a576['h01728] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b95] =  I8a0037ad2845a3fbba9da380a8b8a576['h0172a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b96] =  I8a0037ad2845a3fbba9da380a8b8a576['h0172c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b97] =  I8a0037ad2845a3fbba9da380a8b8a576['h0172e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b98] =  I8a0037ad2845a3fbba9da380a8b8a576['h01730] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b99] =  I8a0037ad2845a3fbba9da380a8b8a576['h01732] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b9a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01734] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b9b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01736] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b9c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01738] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b9d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0173a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b9e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0173c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00b9f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0173e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ba0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01740] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ba1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01742] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ba2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01744] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ba3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01746] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ba4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01748] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ba5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0174a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ba6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0174c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ba7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0174e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ba8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01750] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ba9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01752] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00baa] =  I8a0037ad2845a3fbba9da380a8b8a576['h01754] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bab] =  I8a0037ad2845a3fbba9da380a8b8a576['h01756] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bac] =  I8a0037ad2845a3fbba9da380a8b8a576['h01758] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0175a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0175c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00baf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0175e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bb0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01760] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bb1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01762] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bb2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01764] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bb3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01766] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bb4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01768] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bb5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0176a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bb6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0176c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bb7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0176e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bb8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01770] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bb9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01772] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bba] =  I8a0037ad2845a3fbba9da380a8b8a576['h01774] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bbb] =  I8a0037ad2845a3fbba9da380a8b8a576['h01776] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bbc] =  I8a0037ad2845a3fbba9da380a8b8a576['h01778] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bbd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0177a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bbe] =  I8a0037ad2845a3fbba9da380a8b8a576['h0177c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bbf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0177e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bc0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01780] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bc1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01782] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bc2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01784] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bc3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01786] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bc4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01788] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bc5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0178a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bc6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0178c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bc7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0178e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bc8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01790] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bc9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01792] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bca] =  I8a0037ad2845a3fbba9da380a8b8a576['h01794] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bcb] =  I8a0037ad2845a3fbba9da380a8b8a576['h01796] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bcc] =  I8a0037ad2845a3fbba9da380a8b8a576['h01798] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bcd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0179a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0179c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bcf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0179e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bd0] =  I8a0037ad2845a3fbba9da380a8b8a576['h017a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bd1] =  I8a0037ad2845a3fbba9da380a8b8a576['h017a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bd2] =  I8a0037ad2845a3fbba9da380a8b8a576['h017a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bd3] =  I8a0037ad2845a3fbba9da380a8b8a576['h017a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bd4] =  I8a0037ad2845a3fbba9da380a8b8a576['h017a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bd5] =  I8a0037ad2845a3fbba9da380a8b8a576['h017aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bd6] =  I8a0037ad2845a3fbba9da380a8b8a576['h017ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bd7] =  I8a0037ad2845a3fbba9da380a8b8a576['h017ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bd8] =  I8a0037ad2845a3fbba9da380a8b8a576['h017b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bd9] =  I8a0037ad2845a3fbba9da380a8b8a576['h017b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bda] =  I8a0037ad2845a3fbba9da380a8b8a576['h017b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bdb] =  I8a0037ad2845a3fbba9da380a8b8a576['h017b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bdc] =  I8a0037ad2845a3fbba9da380a8b8a576['h017b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bdd] =  I8a0037ad2845a3fbba9da380a8b8a576['h017ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bde] =  I8a0037ad2845a3fbba9da380a8b8a576['h017bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bdf] =  I8a0037ad2845a3fbba9da380a8b8a576['h017be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00be0] =  I8a0037ad2845a3fbba9da380a8b8a576['h017c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00be1] =  I8a0037ad2845a3fbba9da380a8b8a576['h017c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00be2] =  I8a0037ad2845a3fbba9da380a8b8a576['h017c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00be3] =  I8a0037ad2845a3fbba9da380a8b8a576['h017c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00be4] =  I8a0037ad2845a3fbba9da380a8b8a576['h017c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00be5] =  I8a0037ad2845a3fbba9da380a8b8a576['h017ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00be6] =  I8a0037ad2845a3fbba9da380a8b8a576['h017cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00be7] =  I8a0037ad2845a3fbba9da380a8b8a576['h017ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00be8] =  I8a0037ad2845a3fbba9da380a8b8a576['h017d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00be9] =  I8a0037ad2845a3fbba9da380a8b8a576['h017d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bea] =  I8a0037ad2845a3fbba9da380a8b8a576['h017d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00beb] =  I8a0037ad2845a3fbba9da380a8b8a576['h017d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bec] =  I8a0037ad2845a3fbba9da380a8b8a576['h017d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bed] =  I8a0037ad2845a3fbba9da380a8b8a576['h017da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bee] =  I8a0037ad2845a3fbba9da380a8b8a576['h017dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bef] =  I8a0037ad2845a3fbba9da380a8b8a576['h017de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bf0] =  I8a0037ad2845a3fbba9da380a8b8a576['h017e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bf1] =  I8a0037ad2845a3fbba9da380a8b8a576['h017e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bf2] =  I8a0037ad2845a3fbba9da380a8b8a576['h017e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bf3] =  I8a0037ad2845a3fbba9da380a8b8a576['h017e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bf4] =  I8a0037ad2845a3fbba9da380a8b8a576['h017e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bf5] =  I8a0037ad2845a3fbba9da380a8b8a576['h017ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bf6] =  I8a0037ad2845a3fbba9da380a8b8a576['h017ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bf7] =  I8a0037ad2845a3fbba9da380a8b8a576['h017ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bf8] =  I8a0037ad2845a3fbba9da380a8b8a576['h017f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bf9] =  I8a0037ad2845a3fbba9da380a8b8a576['h017f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bfa] =  I8a0037ad2845a3fbba9da380a8b8a576['h017f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bfb] =  I8a0037ad2845a3fbba9da380a8b8a576['h017f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bfc] =  I8a0037ad2845a3fbba9da380a8b8a576['h017f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bfd] =  I8a0037ad2845a3fbba9da380a8b8a576['h017fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bfe] =  I8a0037ad2845a3fbba9da380a8b8a576['h017fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00bff] =  I8a0037ad2845a3fbba9da380a8b8a576['h017fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c00] =  I8a0037ad2845a3fbba9da380a8b8a576['h01800] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c01] =  I8a0037ad2845a3fbba9da380a8b8a576['h01802] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c02] =  I8a0037ad2845a3fbba9da380a8b8a576['h01804] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c03] =  I8a0037ad2845a3fbba9da380a8b8a576['h01806] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c04] =  I8a0037ad2845a3fbba9da380a8b8a576['h01808] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c05] =  I8a0037ad2845a3fbba9da380a8b8a576['h0180a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c06] =  I8a0037ad2845a3fbba9da380a8b8a576['h0180c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c07] =  I8a0037ad2845a3fbba9da380a8b8a576['h0180e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c08] =  I8a0037ad2845a3fbba9da380a8b8a576['h01810] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c09] =  I8a0037ad2845a3fbba9da380a8b8a576['h01812] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c0a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01814] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c0b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01816] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c0c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01818] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c0d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0181a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c0e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0181c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c0f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0181e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c10] =  I8a0037ad2845a3fbba9da380a8b8a576['h01820] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c11] =  I8a0037ad2845a3fbba9da380a8b8a576['h01822] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c12] =  I8a0037ad2845a3fbba9da380a8b8a576['h01824] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c13] =  I8a0037ad2845a3fbba9da380a8b8a576['h01826] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c14] =  I8a0037ad2845a3fbba9da380a8b8a576['h01828] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c15] =  I8a0037ad2845a3fbba9da380a8b8a576['h0182a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c16] =  I8a0037ad2845a3fbba9da380a8b8a576['h0182c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c17] =  I8a0037ad2845a3fbba9da380a8b8a576['h0182e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c18] =  I8a0037ad2845a3fbba9da380a8b8a576['h01830] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c19] =  I8a0037ad2845a3fbba9da380a8b8a576['h01832] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c1a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01834] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c1b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01836] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c1c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01838] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c1d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0183a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c1e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0183c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c1f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0183e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c20] =  I8a0037ad2845a3fbba9da380a8b8a576['h01840] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c21] =  I8a0037ad2845a3fbba9da380a8b8a576['h01842] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c22] =  I8a0037ad2845a3fbba9da380a8b8a576['h01844] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c23] =  I8a0037ad2845a3fbba9da380a8b8a576['h01846] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c24] =  I8a0037ad2845a3fbba9da380a8b8a576['h01848] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c25] =  I8a0037ad2845a3fbba9da380a8b8a576['h0184a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c26] =  I8a0037ad2845a3fbba9da380a8b8a576['h0184c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c27] =  I8a0037ad2845a3fbba9da380a8b8a576['h0184e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c28] =  I8a0037ad2845a3fbba9da380a8b8a576['h01850] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c29] =  I8a0037ad2845a3fbba9da380a8b8a576['h01852] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c2a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01854] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c2b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01856] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c2c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01858] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c2d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0185a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c2e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0185c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c2f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0185e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c30] =  I8a0037ad2845a3fbba9da380a8b8a576['h01860] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c31] =  I8a0037ad2845a3fbba9da380a8b8a576['h01862] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c32] =  I8a0037ad2845a3fbba9da380a8b8a576['h01864] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c33] =  I8a0037ad2845a3fbba9da380a8b8a576['h01866] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c34] =  I8a0037ad2845a3fbba9da380a8b8a576['h01868] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c35] =  I8a0037ad2845a3fbba9da380a8b8a576['h0186a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c36] =  I8a0037ad2845a3fbba9da380a8b8a576['h0186c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c37] =  I8a0037ad2845a3fbba9da380a8b8a576['h0186e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c38] =  I8a0037ad2845a3fbba9da380a8b8a576['h01870] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c39] =  I8a0037ad2845a3fbba9da380a8b8a576['h01872] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c3a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01874] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c3b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01876] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c3c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01878] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c3d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0187a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c3e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0187c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c3f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0187e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c40] =  I8a0037ad2845a3fbba9da380a8b8a576['h01880] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c41] =  I8a0037ad2845a3fbba9da380a8b8a576['h01882] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c42] =  I8a0037ad2845a3fbba9da380a8b8a576['h01884] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c43] =  I8a0037ad2845a3fbba9da380a8b8a576['h01886] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c44] =  I8a0037ad2845a3fbba9da380a8b8a576['h01888] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c45] =  I8a0037ad2845a3fbba9da380a8b8a576['h0188a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c46] =  I8a0037ad2845a3fbba9da380a8b8a576['h0188c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c47] =  I8a0037ad2845a3fbba9da380a8b8a576['h0188e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c48] =  I8a0037ad2845a3fbba9da380a8b8a576['h01890] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c49] =  I8a0037ad2845a3fbba9da380a8b8a576['h01892] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c4a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01894] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c4b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01896] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c4c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01898] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c4d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0189a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c4e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0189c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c4f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0189e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c50] =  I8a0037ad2845a3fbba9da380a8b8a576['h018a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c51] =  I8a0037ad2845a3fbba9da380a8b8a576['h018a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c52] =  I8a0037ad2845a3fbba9da380a8b8a576['h018a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c53] =  I8a0037ad2845a3fbba9da380a8b8a576['h018a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c54] =  I8a0037ad2845a3fbba9da380a8b8a576['h018a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c55] =  I8a0037ad2845a3fbba9da380a8b8a576['h018aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c56] =  I8a0037ad2845a3fbba9da380a8b8a576['h018ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c57] =  I8a0037ad2845a3fbba9da380a8b8a576['h018ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c58] =  I8a0037ad2845a3fbba9da380a8b8a576['h018b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c59] =  I8a0037ad2845a3fbba9da380a8b8a576['h018b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c5a] =  I8a0037ad2845a3fbba9da380a8b8a576['h018b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c5b] =  I8a0037ad2845a3fbba9da380a8b8a576['h018b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c5c] =  I8a0037ad2845a3fbba9da380a8b8a576['h018b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c5d] =  I8a0037ad2845a3fbba9da380a8b8a576['h018ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c5e] =  I8a0037ad2845a3fbba9da380a8b8a576['h018bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c5f] =  I8a0037ad2845a3fbba9da380a8b8a576['h018be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c60] =  I8a0037ad2845a3fbba9da380a8b8a576['h018c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c61] =  I8a0037ad2845a3fbba9da380a8b8a576['h018c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c62] =  I8a0037ad2845a3fbba9da380a8b8a576['h018c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c63] =  I8a0037ad2845a3fbba9da380a8b8a576['h018c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c64] =  I8a0037ad2845a3fbba9da380a8b8a576['h018c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c65] =  I8a0037ad2845a3fbba9da380a8b8a576['h018ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c66] =  I8a0037ad2845a3fbba9da380a8b8a576['h018cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c67] =  I8a0037ad2845a3fbba9da380a8b8a576['h018ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c68] =  I8a0037ad2845a3fbba9da380a8b8a576['h018d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c69] =  I8a0037ad2845a3fbba9da380a8b8a576['h018d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c6a] =  I8a0037ad2845a3fbba9da380a8b8a576['h018d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c6b] =  I8a0037ad2845a3fbba9da380a8b8a576['h018d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c6c] =  I8a0037ad2845a3fbba9da380a8b8a576['h018d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c6d] =  I8a0037ad2845a3fbba9da380a8b8a576['h018da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c6e] =  I8a0037ad2845a3fbba9da380a8b8a576['h018dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c6f] =  I8a0037ad2845a3fbba9da380a8b8a576['h018de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c70] =  I8a0037ad2845a3fbba9da380a8b8a576['h018e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c71] =  I8a0037ad2845a3fbba9da380a8b8a576['h018e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c72] =  I8a0037ad2845a3fbba9da380a8b8a576['h018e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c73] =  I8a0037ad2845a3fbba9da380a8b8a576['h018e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c74] =  I8a0037ad2845a3fbba9da380a8b8a576['h018e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c75] =  I8a0037ad2845a3fbba9da380a8b8a576['h018ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c76] =  I8a0037ad2845a3fbba9da380a8b8a576['h018ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c77] =  I8a0037ad2845a3fbba9da380a8b8a576['h018ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c78] =  I8a0037ad2845a3fbba9da380a8b8a576['h018f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c79] =  I8a0037ad2845a3fbba9da380a8b8a576['h018f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c7a] =  I8a0037ad2845a3fbba9da380a8b8a576['h018f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c7b] =  I8a0037ad2845a3fbba9da380a8b8a576['h018f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c7c] =  I8a0037ad2845a3fbba9da380a8b8a576['h018f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c7d] =  I8a0037ad2845a3fbba9da380a8b8a576['h018fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c7e] =  I8a0037ad2845a3fbba9da380a8b8a576['h018fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c7f] =  I8a0037ad2845a3fbba9da380a8b8a576['h018fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c80] =  I8a0037ad2845a3fbba9da380a8b8a576['h01900] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c81] =  I8a0037ad2845a3fbba9da380a8b8a576['h01902] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c82] =  I8a0037ad2845a3fbba9da380a8b8a576['h01904] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c83] =  I8a0037ad2845a3fbba9da380a8b8a576['h01906] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c84] =  I8a0037ad2845a3fbba9da380a8b8a576['h01908] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c85] =  I8a0037ad2845a3fbba9da380a8b8a576['h0190a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c86] =  I8a0037ad2845a3fbba9da380a8b8a576['h0190c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c87] =  I8a0037ad2845a3fbba9da380a8b8a576['h0190e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c88] =  I8a0037ad2845a3fbba9da380a8b8a576['h01910] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c89] =  I8a0037ad2845a3fbba9da380a8b8a576['h01912] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c8a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01914] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c8b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01916] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c8c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01918] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c8d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0191a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c8e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0191c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c8f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0191e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c90] =  I8a0037ad2845a3fbba9da380a8b8a576['h01920] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c91] =  I8a0037ad2845a3fbba9da380a8b8a576['h01922] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c92] =  I8a0037ad2845a3fbba9da380a8b8a576['h01924] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c93] =  I8a0037ad2845a3fbba9da380a8b8a576['h01926] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c94] =  I8a0037ad2845a3fbba9da380a8b8a576['h01928] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c95] =  I8a0037ad2845a3fbba9da380a8b8a576['h0192a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c96] =  I8a0037ad2845a3fbba9da380a8b8a576['h0192c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c97] =  I8a0037ad2845a3fbba9da380a8b8a576['h0192e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c98] =  I8a0037ad2845a3fbba9da380a8b8a576['h01930] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c99] =  I8a0037ad2845a3fbba9da380a8b8a576['h01932] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c9a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01934] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c9b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01936] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c9c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01938] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c9d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0193a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c9e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0193c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00c9f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0193e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ca0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01940] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ca1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01942] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ca2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01944] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ca3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01946] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ca4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01948] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ca5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0194a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ca6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0194c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ca7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0194e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ca8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01950] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ca9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01952] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00caa] =  I8a0037ad2845a3fbba9da380a8b8a576['h01954] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cab] =  I8a0037ad2845a3fbba9da380a8b8a576['h01956] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cac] =  I8a0037ad2845a3fbba9da380a8b8a576['h01958] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0195a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0195c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00caf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0195e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cb0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01960] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cb1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01962] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cb2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01964] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cb3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01966] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cb4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01968] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cb5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0196a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cb6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0196c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cb7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0196e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cb8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01970] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cb9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01972] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cba] =  I8a0037ad2845a3fbba9da380a8b8a576['h01974] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cbb] =  I8a0037ad2845a3fbba9da380a8b8a576['h01976] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cbc] =  I8a0037ad2845a3fbba9da380a8b8a576['h01978] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cbd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0197a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cbe] =  I8a0037ad2845a3fbba9da380a8b8a576['h0197c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cbf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0197e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cc0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01980] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cc1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01982] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cc2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01984] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cc3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01986] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cc4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01988] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cc5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0198a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cc6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0198c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cc7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0198e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cc8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01990] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cc9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01992] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cca] =  I8a0037ad2845a3fbba9da380a8b8a576['h01994] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ccb] =  I8a0037ad2845a3fbba9da380a8b8a576['h01996] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ccc] =  I8a0037ad2845a3fbba9da380a8b8a576['h01998] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ccd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0199a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0199c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ccf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0199e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cd0] =  I8a0037ad2845a3fbba9da380a8b8a576['h019a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cd1] =  I8a0037ad2845a3fbba9da380a8b8a576['h019a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cd2] =  I8a0037ad2845a3fbba9da380a8b8a576['h019a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cd3] =  I8a0037ad2845a3fbba9da380a8b8a576['h019a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cd4] =  I8a0037ad2845a3fbba9da380a8b8a576['h019a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cd5] =  I8a0037ad2845a3fbba9da380a8b8a576['h019aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cd6] =  I8a0037ad2845a3fbba9da380a8b8a576['h019ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cd7] =  I8a0037ad2845a3fbba9da380a8b8a576['h019ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cd8] =  I8a0037ad2845a3fbba9da380a8b8a576['h019b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cd9] =  I8a0037ad2845a3fbba9da380a8b8a576['h019b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cda] =  I8a0037ad2845a3fbba9da380a8b8a576['h019b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cdb] =  I8a0037ad2845a3fbba9da380a8b8a576['h019b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cdc] =  I8a0037ad2845a3fbba9da380a8b8a576['h019b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cdd] =  I8a0037ad2845a3fbba9da380a8b8a576['h019ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cde] =  I8a0037ad2845a3fbba9da380a8b8a576['h019bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cdf] =  I8a0037ad2845a3fbba9da380a8b8a576['h019be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ce0] =  I8a0037ad2845a3fbba9da380a8b8a576['h019c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ce1] =  I8a0037ad2845a3fbba9da380a8b8a576['h019c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ce2] =  I8a0037ad2845a3fbba9da380a8b8a576['h019c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ce3] =  I8a0037ad2845a3fbba9da380a8b8a576['h019c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ce4] =  I8a0037ad2845a3fbba9da380a8b8a576['h019c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ce5] =  I8a0037ad2845a3fbba9da380a8b8a576['h019ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ce6] =  I8a0037ad2845a3fbba9da380a8b8a576['h019cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ce7] =  I8a0037ad2845a3fbba9da380a8b8a576['h019ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ce8] =  I8a0037ad2845a3fbba9da380a8b8a576['h019d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ce9] =  I8a0037ad2845a3fbba9da380a8b8a576['h019d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cea] =  I8a0037ad2845a3fbba9da380a8b8a576['h019d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ceb] =  I8a0037ad2845a3fbba9da380a8b8a576['h019d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cec] =  I8a0037ad2845a3fbba9da380a8b8a576['h019d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ced] =  I8a0037ad2845a3fbba9da380a8b8a576['h019da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cee] =  I8a0037ad2845a3fbba9da380a8b8a576['h019dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cef] =  I8a0037ad2845a3fbba9da380a8b8a576['h019de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cf0] =  I8a0037ad2845a3fbba9da380a8b8a576['h019e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cf1] =  I8a0037ad2845a3fbba9da380a8b8a576['h019e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cf2] =  I8a0037ad2845a3fbba9da380a8b8a576['h019e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cf3] =  I8a0037ad2845a3fbba9da380a8b8a576['h019e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cf4] =  I8a0037ad2845a3fbba9da380a8b8a576['h019e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cf5] =  I8a0037ad2845a3fbba9da380a8b8a576['h019ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cf6] =  I8a0037ad2845a3fbba9da380a8b8a576['h019ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cf7] =  I8a0037ad2845a3fbba9da380a8b8a576['h019ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cf8] =  I8a0037ad2845a3fbba9da380a8b8a576['h019f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cf9] =  I8a0037ad2845a3fbba9da380a8b8a576['h019f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cfa] =  I8a0037ad2845a3fbba9da380a8b8a576['h019f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cfb] =  I8a0037ad2845a3fbba9da380a8b8a576['h019f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cfc] =  I8a0037ad2845a3fbba9da380a8b8a576['h019f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cfd] =  I8a0037ad2845a3fbba9da380a8b8a576['h019fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cfe] =  I8a0037ad2845a3fbba9da380a8b8a576['h019fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00cff] =  I8a0037ad2845a3fbba9da380a8b8a576['h019fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d00] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d01] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d02] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d03] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d04] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d05] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d06] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d07] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d08] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d09] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d0a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d0b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d0c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d0d] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d0e] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d0f] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d10] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d11] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d12] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d13] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d14] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d15] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d16] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d17] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d18] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d19] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d1a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d1b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d1c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d1d] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d1e] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d1f] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d20] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d21] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d22] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d23] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d24] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d25] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d26] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d27] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d28] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d29] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d2a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d2b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d2c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d2d] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d2e] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d2f] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d30] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d31] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d32] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d33] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d34] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d35] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d36] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d37] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d38] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d39] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d3a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d3b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d3c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d3d] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d3e] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d3f] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d40] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d41] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d42] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d43] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d44] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d45] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d46] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d47] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d48] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d49] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d4a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d4b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d4c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d4d] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d4e] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d4f] =  I8a0037ad2845a3fbba9da380a8b8a576['h01a9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d50] =  I8a0037ad2845a3fbba9da380a8b8a576['h01aa0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d51] =  I8a0037ad2845a3fbba9da380a8b8a576['h01aa2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d52] =  I8a0037ad2845a3fbba9da380a8b8a576['h01aa4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d53] =  I8a0037ad2845a3fbba9da380a8b8a576['h01aa6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d54] =  I8a0037ad2845a3fbba9da380a8b8a576['h01aa8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d55] =  I8a0037ad2845a3fbba9da380a8b8a576['h01aaa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d56] =  I8a0037ad2845a3fbba9da380a8b8a576['h01aac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d57] =  I8a0037ad2845a3fbba9da380a8b8a576['h01aae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d58] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ab0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d59] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ab2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d5a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ab4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d5b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ab6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d5c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ab8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d5d] =  I8a0037ad2845a3fbba9da380a8b8a576['h01aba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d5e] =  I8a0037ad2845a3fbba9da380a8b8a576['h01abc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d5f] =  I8a0037ad2845a3fbba9da380a8b8a576['h01abe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d60] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ac0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d61] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ac2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d62] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ac4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d63] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ac6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d64] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ac8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d65] =  I8a0037ad2845a3fbba9da380a8b8a576['h01aca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d66] =  I8a0037ad2845a3fbba9da380a8b8a576['h01acc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d67] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ace] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d68] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ad0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d69] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ad2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d6a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ad4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d6b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ad6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d6c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ad8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d6d] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ada] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d6e] =  I8a0037ad2845a3fbba9da380a8b8a576['h01adc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d6f] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ade] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d70] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ae0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d71] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ae2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d72] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ae4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d73] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ae6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d74] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ae8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d75] =  I8a0037ad2845a3fbba9da380a8b8a576['h01aea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d76] =  I8a0037ad2845a3fbba9da380a8b8a576['h01aec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d77] =  I8a0037ad2845a3fbba9da380a8b8a576['h01aee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d78] =  I8a0037ad2845a3fbba9da380a8b8a576['h01af0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d79] =  I8a0037ad2845a3fbba9da380a8b8a576['h01af2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d7a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01af4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d7b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01af6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d7c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01af8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d7d] =  I8a0037ad2845a3fbba9da380a8b8a576['h01afa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d7e] =  I8a0037ad2845a3fbba9da380a8b8a576['h01afc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d7f] =  I8a0037ad2845a3fbba9da380a8b8a576['h01afe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d80] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d81] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d82] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d83] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d84] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d85] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d86] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d87] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d88] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d89] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d8a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d8b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d8c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d8d] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d8e] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d8f] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d90] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d91] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d92] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d93] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d94] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d95] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d96] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d97] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d98] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d99] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d9a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d9b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d9c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d9d] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d9e] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00d9f] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00da0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00da1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00da2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00da3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00da4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00da5] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00da6] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00da7] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00da8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00da9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00daa] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dab] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dac] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dad] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dae] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00daf] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00db0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00db1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00db2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00db3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00db4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00db5] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00db6] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00db7] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00db8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00db9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dba] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dbb] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dbc] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dbd] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dbe] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dbf] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dc0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dc1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dc2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dc3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dc4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dc5] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dc6] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dc7] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dc8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dc9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dca] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dcb] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dcc] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dcd] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dce] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dcf] =  I8a0037ad2845a3fbba9da380a8b8a576['h01b9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dd0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ba0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dd1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ba2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dd2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ba4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dd3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ba6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dd4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ba8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dd5] =  I8a0037ad2845a3fbba9da380a8b8a576['h01baa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dd6] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dd7] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dd8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dd9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dda] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ddb] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ddc] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ddd] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dde] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ddf] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00de0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00de1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00de2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00de3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00de4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00de5] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00de6] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bcc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00de7] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00de8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00de9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dea] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00deb] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dec] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ded] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dee] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bdc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00def] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00df0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01be0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00df1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01be2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00df2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01be4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00df3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01be6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00df4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01be8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00df5] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00df6] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00df7] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00df8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bf0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00df9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bf2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dfa] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bf4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dfb] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bf6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dfc] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bf8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dfd] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bfa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dfe] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bfc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00dff] =  I8a0037ad2845a3fbba9da380a8b8a576['h01bfe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e00] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e01] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e02] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e03] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e04] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e05] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e06] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e07] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e08] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e09] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e0a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e0b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e0c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e0d] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e0e] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e0f] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e10] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e11] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e12] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e13] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e14] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e15] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e16] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e17] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e18] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e19] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e1a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e1b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e1c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e1d] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e1e] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e1f] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e20] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e21] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e22] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e23] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e24] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e25] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e26] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e27] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e28] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e29] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e2a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e2b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e2c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e2d] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e2e] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e2f] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e30] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e31] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e32] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e33] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e34] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e35] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e36] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e37] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e38] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e39] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e3a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e3b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e3c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e3d] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e3e] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e3f] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e40] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e41] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e42] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e43] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e44] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e45] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e46] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e47] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e48] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e49] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e4a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e4b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e4c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e4d] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e4e] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e4f] =  I8a0037ad2845a3fbba9da380a8b8a576['h01c9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e50] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ca0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e51] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ca2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e52] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ca4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e53] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ca6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e54] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ca8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e55] =  I8a0037ad2845a3fbba9da380a8b8a576['h01caa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e56] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e57] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e58] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e59] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e5a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e5b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e5c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e5d] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e5e] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e5f] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e60] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e61] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e62] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e63] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e64] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e65] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e66] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ccc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e67] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e68] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e69] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e6a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e6b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e6c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e6d] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e6e] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cdc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e6f] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e70] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ce0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e71] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ce2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e72] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ce4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e73] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ce6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e74] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ce8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e75] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e76] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e77] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e78] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cf0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e79] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cf2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e7a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cf4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e7b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cf6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e7c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cf8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e7d] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cfa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e7e] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cfc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e7f] =  I8a0037ad2845a3fbba9da380a8b8a576['h01cfe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e80] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e81] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e82] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e83] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e84] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e85] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e86] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e87] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e88] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e89] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e8a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e8b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e8c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e8d] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e8e] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e8f] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e90] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e91] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e92] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e93] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e94] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e95] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e96] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e97] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e98] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e99] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e9a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e9b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e9c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e9d] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e9e] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00e9f] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ea0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ea1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ea2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ea3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ea4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ea5] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ea6] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ea7] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ea8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ea9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00eaa] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00eab] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00eac] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ead] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00eae] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00eaf] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00eb0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00eb1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00eb2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00eb3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00eb4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00eb5] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00eb6] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00eb7] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00eb8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00eb9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00eba] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ebb] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ebc] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ebd] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ebe] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ebf] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ec0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ec1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ec2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ec3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ec4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ec5] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ec6] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ec7] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ec8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ec9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00eca] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ecb] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ecc] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ecd] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ece] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ecf] =  I8a0037ad2845a3fbba9da380a8b8a576['h01d9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ed0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01da0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ed1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01da2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ed2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01da4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ed3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01da6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ed4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01da8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ed5] =  I8a0037ad2845a3fbba9da380a8b8a576['h01daa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ed6] =  I8a0037ad2845a3fbba9da380a8b8a576['h01dac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ed7] =  I8a0037ad2845a3fbba9da380a8b8a576['h01dae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ed8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01db0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ed9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01db2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00eda] =  I8a0037ad2845a3fbba9da380a8b8a576['h01db4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00edb] =  I8a0037ad2845a3fbba9da380a8b8a576['h01db6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00edc] =  I8a0037ad2845a3fbba9da380a8b8a576['h01db8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00edd] =  I8a0037ad2845a3fbba9da380a8b8a576['h01dba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ede] =  I8a0037ad2845a3fbba9da380a8b8a576['h01dbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00edf] =  I8a0037ad2845a3fbba9da380a8b8a576['h01dbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ee0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01dc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ee1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01dc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ee2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01dc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ee3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01dc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ee4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01dc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ee5] =  I8a0037ad2845a3fbba9da380a8b8a576['h01dca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ee6] =  I8a0037ad2845a3fbba9da380a8b8a576['h01dcc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ee7] =  I8a0037ad2845a3fbba9da380a8b8a576['h01dce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ee8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01dd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ee9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01dd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00eea] =  I8a0037ad2845a3fbba9da380a8b8a576['h01dd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00eeb] =  I8a0037ad2845a3fbba9da380a8b8a576['h01dd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00eec] =  I8a0037ad2845a3fbba9da380a8b8a576['h01dd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00eed] =  I8a0037ad2845a3fbba9da380a8b8a576['h01dda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00eee] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ddc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00eef] =  I8a0037ad2845a3fbba9da380a8b8a576['h01dde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ef0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01de0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ef1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01de2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ef2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01de4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ef3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01de6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ef4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01de8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ef5] =  I8a0037ad2845a3fbba9da380a8b8a576['h01dea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ef6] =  I8a0037ad2845a3fbba9da380a8b8a576['h01dec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ef7] =  I8a0037ad2845a3fbba9da380a8b8a576['h01dee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ef8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01df0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ef9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01df2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00efa] =  I8a0037ad2845a3fbba9da380a8b8a576['h01df4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00efb] =  I8a0037ad2845a3fbba9da380a8b8a576['h01df6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00efc] =  I8a0037ad2845a3fbba9da380a8b8a576['h01df8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00efd] =  I8a0037ad2845a3fbba9da380a8b8a576['h01dfa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00efe] =  I8a0037ad2845a3fbba9da380a8b8a576['h01dfc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00eff] =  I8a0037ad2845a3fbba9da380a8b8a576['h01dfe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f00] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f01] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f02] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f03] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f04] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f05] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f06] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f07] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f08] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f09] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f0a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f0b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f0c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f0d] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f0e] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f0f] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f10] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f11] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f12] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f13] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f14] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f15] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f16] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f17] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f18] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f19] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f1a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f1b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f1c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f1d] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f1e] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f1f] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f20] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f21] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f22] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f23] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f24] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f25] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f26] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f27] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f28] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f29] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f2a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f2b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f2c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f2d] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f2e] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f2f] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f30] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f31] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f32] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f33] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f34] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f35] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f36] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f37] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f38] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f39] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f3a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f3b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f3c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f3d] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f3e] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f3f] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f40] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f41] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f42] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f43] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f44] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f45] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f46] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f47] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f48] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f49] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f4a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f4b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f4c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f4d] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f4e] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f4f] =  I8a0037ad2845a3fbba9da380a8b8a576['h01e9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f50] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ea0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f51] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ea2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f52] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ea4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f53] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ea6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f54] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ea8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f55] =  I8a0037ad2845a3fbba9da380a8b8a576['h01eaa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f56] =  I8a0037ad2845a3fbba9da380a8b8a576['h01eac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f57] =  I8a0037ad2845a3fbba9da380a8b8a576['h01eae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f58] =  I8a0037ad2845a3fbba9da380a8b8a576['h01eb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f59] =  I8a0037ad2845a3fbba9da380a8b8a576['h01eb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f5a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01eb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f5b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01eb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f5c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01eb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f5d] =  I8a0037ad2845a3fbba9da380a8b8a576['h01eba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f5e] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ebc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f5f] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ebe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f60] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ec0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f61] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ec2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f62] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ec4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f63] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ec6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f64] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ec8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f65] =  I8a0037ad2845a3fbba9da380a8b8a576['h01eca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f66] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ecc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f67] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ece] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f68] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ed0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f69] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ed2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f6a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ed4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f6b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ed6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f6c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ed8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f6d] =  I8a0037ad2845a3fbba9da380a8b8a576['h01eda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f6e] =  I8a0037ad2845a3fbba9da380a8b8a576['h01edc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f6f] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ede] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f70] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ee0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f71] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ee2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f72] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ee4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f73] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ee6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f74] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ee8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f75] =  I8a0037ad2845a3fbba9da380a8b8a576['h01eea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f76] =  I8a0037ad2845a3fbba9da380a8b8a576['h01eec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f77] =  I8a0037ad2845a3fbba9da380a8b8a576['h01eee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f78] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ef0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f79] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ef2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f7a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ef4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f7b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ef6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f7c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ef8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f7d] =  I8a0037ad2845a3fbba9da380a8b8a576['h01efa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f7e] =  I8a0037ad2845a3fbba9da380a8b8a576['h01efc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f7f] =  I8a0037ad2845a3fbba9da380a8b8a576['h01efe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f80] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f81] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f82] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f83] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f84] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f85] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f86] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f87] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f88] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f89] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f8a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f8b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f8c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f8d] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f8e] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f8f] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f90] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f91] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f92] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f93] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f94] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f95] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f96] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f97] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f98] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f99] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f9a] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f9b] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f9c] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f9d] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f9e] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00f9f] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fa0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fa1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fa2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fa3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fa4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fa5] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fa6] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fa7] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fa8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fa9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00faa] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fab] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fac] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fad] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fae] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00faf] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fb0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fb1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fb2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fb3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fb4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fb5] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fb6] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fb7] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fb8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fb9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fba] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fbb] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fbc] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fbd] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fbe] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fbf] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fc0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fc1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fc2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fc3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fc4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fc5] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fc6] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fc7] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fc8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fc9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fca] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fcb] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fcc] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fcd] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fce] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fcf] =  I8a0037ad2845a3fbba9da380a8b8a576['h01f9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fd0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fa0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fd1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fa2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fd2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fa4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fd3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fa6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fd4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fa8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fd5] =  I8a0037ad2845a3fbba9da380a8b8a576['h01faa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fd6] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fd7] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fd8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fd9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fda] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fdb] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fdc] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fdd] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fde] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fdf] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fe0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fe1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fe2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fe3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fe4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fe5] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fe6] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fcc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fe7] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fe8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fe9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fea] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00feb] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fec] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fed] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fee] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fdc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fef] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ff0] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fe0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ff1] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fe2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ff2] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fe4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ff3] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fe6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ff4] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fe8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ff5] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ff6] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ff7] =  I8a0037ad2845a3fbba9da380a8b8a576['h01fee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ff8] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ff0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ff9] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ff2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ffa] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ff4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ffb] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ff6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ffc] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ff8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ffd] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ffa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00ffe] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ffc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h00fff] =  I8a0037ad2845a3fbba9da380a8b8a576['h01ffe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01000] =  I8a0037ad2845a3fbba9da380a8b8a576['h02000] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01001] =  I8a0037ad2845a3fbba9da380a8b8a576['h02002] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01002] =  I8a0037ad2845a3fbba9da380a8b8a576['h02004] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01003] =  I8a0037ad2845a3fbba9da380a8b8a576['h02006] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01004] =  I8a0037ad2845a3fbba9da380a8b8a576['h02008] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01005] =  I8a0037ad2845a3fbba9da380a8b8a576['h0200a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01006] =  I8a0037ad2845a3fbba9da380a8b8a576['h0200c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01007] =  I8a0037ad2845a3fbba9da380a8b8a576['h0200e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01008] =  I8a0037ad2845a3fbba9da380a8b8a576['h02010] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01009] =  I8a0037ad2845a3fbba9da380a8b8a576['h02012] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0100a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02014] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0100b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02016] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0100c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02018] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0100d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0201a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0100e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0201c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0100f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0201e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01010] =  I8a0037ad2845a3fbba9da380a8b8a576['h02020] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01011] =  I8a0037ad2845a3fbba9da380a8b8a576['h02022] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01012] =  I8a0037ad2845a3fbba9da380a8b8a576['h02024] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01013] =  I8a0037ad2845a3fbba9da380a8b8a576['h02026] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01014] =  I8a0037ad2845a3fbba9da380a8b8a576['h02028] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01015] =  I8a0037ad2845a3fbba9da380a8b8a576['h0202a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01016] =  I8a0037ad2845a3fbba9da380a8b8a576['h0202c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01017] =  I8a0037ad2845a3fbba9da380a8b8a576['h0202e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01018] =  I8a0037ad2845a3fbba9da380a8b8a576['h02030] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01019] =  I8a0037ad2845a3fbba9da380a8b8a576['h02032] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0101a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02034] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0101b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02036] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0101c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02038] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0101d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0203a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0101e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0203c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0101f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0203e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01020] =  I8a0037ad2845a3fbba9da380a8b8a576['h02040] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01021] =  I8a0037ad2845a3fbba9da380a8b8a576['h02042] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01022] =  I8a0037ad2845a3fbba9da380a8b8a576['h02044] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01023] =  I8a0037ad2845a3fbba9da380a8b8a576['h02046] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01024] =  I8a0037ad2845a3fbba9da380a8b8a576['h02048] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01025] =  I8a0037ad2845a3fbba9da380a8b8a576['h0204a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01026] =  I8a0037ad2845a3fbba9da380a8b8a576['h0204c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01027] =  I8a0037ad2845a3fbba9da380a8b8a576['h0204e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01028] =  I8a0037ad2845a3fbba9da380a8b8a576['h02050] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01029] =  I8a0037ad2845a3fbba9da380a8b8a576['h02052] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0102a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02054] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0102b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02056] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0102c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02058] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0102d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0205a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0102e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0205c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0102f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0205e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01030] =  I8a0037ad2845a3fbba9da380a8b8a576['h02060] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01031] =  I8a0037ad2845a3fbba9da380a8b8a576['h02062] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01032] =  I8a0037ad2845a3fbba9da380a8b8a576['h02064] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01033] =  I8a0037ad2845a3fbba9da380a8b8a576['h02066] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01034] =  I8a0037ad2845a3fbba9da380a8b8a576['h02068] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01035] =  I8a0037ad2845a3fbba9da380a8b8a576['h0206a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01036] =  I8a0037ad2845a3fbba9da380a8b8a576['h0206c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01037] =  I8a0037ad2845a3fbba9da380a8b8a576['h0206e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01038] =  I8a0037ad2845a3fbba9da380a8b8a576['h02070] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01039] =  I8a0037ad2845a3fbba9da380a8b8a576['h02072] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0103a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02074] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0103b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02076] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0103c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02078] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0103d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0207a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0103e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0207c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0103f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0207e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01040] =  I8a0037ad2845a3fbba9da380a8b8a576['h02080] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01041] =  I8a0037ad2845a3fbba9da380a8b8a576['h02082] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01042] =  I8a0037ad2845a3fbba9da380a8b8a576['h02084] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01043] =  I8a0037ad2845a3fbba9da380a8b8a576['h02086] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01044] =  I8a0037ad2845a3fbba9da380a8b8a576['h02088] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01045] =  I8a0037ad2845a3fbba9da380a8b8a576['h0208a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01046] =  I8a0037ad2845a3fbba9da380a8b8a576['h0208c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01047] =  I8a0037ad2845a3fbba9da380a8b8a576['h0208e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01048] =  I8a0037ad2845a3fbba9da380a8b8a576['h02090] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01049] =  I8a0037ad2845a3fbba9da380a8b8a576['h02092] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0104a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02094] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0104b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02096] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0104c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02098] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0104d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0209a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0104e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0209c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0104f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0209e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01050] =  I8a0037ad2845a3fbba9da380a8b8a576['h020a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01051] =  I8a0037ad2845a3fbba9da380a8b8a576['h020a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01052] =  I8a0037ad2845a3fbba9da380a8b8a576['h020a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01053] =  I8a0037ad2845a3fbba9da380a8b8a576['h020a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01054] =  I8a0037ad2845a3fbba9da380a8b8a576['h020a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01055] =  I8a0037ad2845a3fbba9da380a8b8a576['h020aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01056] =  I8a0037ad2845a3fbba9da380a8b8a576['h020ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01057] =  I8a0037ad2845a3fbba9da380a8b8a576['h020ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01058] =  I8a0037ad2845a3fbba9da380a8b8a576['h020b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01059] =  I8a0037ad2845a3fbba9da380a8b8a576['h020b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0105a] =  I8a0037ad2845a3fbba9da380a8b8a576['h020b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0105b] =  I8a0037ad2845a3fbba9da380a8b8a576['h020b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0105c] =  I8a0037ad2845a3fbba9da380a8b8a576['h020b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0105d] =  I8a0037ad2845a3fbba9da380a8b8a576['h020ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0105e] =  I8a0037ad2845a3fbba9da380a8b8a576['h020bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0105f] =  I8a0037ad2845a3fbba9da380a8b8a576['h020be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01060] =  I8a0037ad2845a3fbba9da380a8b8a576['h020c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01061] =  I8a0037ad2845a3fbba9da380a8b8a576['h020c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01062] =  I8a0037ad2845a3fbba9da380a8b8a576['h020c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01063] =  I8a0037ad2845a3fbba9da380a8b8a576['h020c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01064] =  I8a0037ad2845a3fbba9da380a8b8a576['h020c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01065] =  I8a0037ad2845a3fbba9da380a8b8a576['h020ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01066] =  I8a0037ad2845a3fbba9da380a8b8a576['h020cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01067] =  I8a0037ad2845a3fbba9da380a8b8a576['h020ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01068] =  I8a0037ad2845a3fbba9da380a8b8a576['h020d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01069] =  I8a0037ad2845a3fbba9da380a8b8a576['h020d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0106a] =  I8a0037ad2845a3fbba9da380a8b8a576['h020d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0106b] =  I8a0037ad2845a3fbba9da380a8b8a576['h020d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0106c] =  I8a0037ad2845a3fbba9da380a8b8a576['h020d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0106d] =  I8a0037ad2845a3fbba9da380a8b8a576['h020da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0106e] =  I8a0037ad2845a3fbba9da380a8b8a576['h020dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0106f] =  I8a0037ad2845a3fbba9da380a8b8a576['h020de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01070] =  I8a0037ad2845a3fbba9da380a8b8a576['h020e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01071] =  I8a0037ad2845a3fbba9da380a8b8a576['h020e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01072] =  I8a0037ad2845a3fbba9da380a8b8a576['h020e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01073] =  I8a0037ad2845a3fbba9da380a8b8a576['h020e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01074] =  I8a0037ad2845a3fbba9da380a8b8a576['h020e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01075] =  I8a0037ad2845a3fbba9da380a8b8a576['h020ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01076] =  I8a0037ad2845a3fbba9da380a8b8a576['h020ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01077] =  I8a0037ad2845a3fbba9da380a8b8a576['h020ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01078] =  I8a0037ad2845a3fbba9da380a8b8a576['h020f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01079] =  I8a0037ad2845a3fbba9da380a8b8a576['h020f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0107a] =  I8a0037ad2845a3fbba9da380a8b8a576['h020f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0107b] =  I8a0037ad2845a3fbba9da380a8b8a576['h020f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0107c] =  I8a0037ad2845a3fbba9da380a8b8a576['h020f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0107d] =  I8a0037ad2845a3fbba9da380a8b8a576['h020fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0107e] =  I8a0037ad2845a3fbba9da380a8b8a576['h020fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0107f] =  I8a0037ad2845a3fbba9da380a8b8a576['h020fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01080] =  I8a0037ad2845a3fbba9da380a8b8a576['h02100] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01081] =  I8a0037ad2845a3fbba9da380a8b8a576['h02102] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01082] =  I8a0037ad2845a3fbba9da380a8b8a576['h02104] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01083] =  I8a0037ad2845a3fbba9da380a8b8a576['h02106] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01084] =  I8a0037ad2845a3fbba9da380a8b8a576['h02108] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01085] =  I8a0037ad2845a3fbba9da380a8b8a576['h0210a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01086] =  I8a0037ad2845a3fbba9da380a8b8a576['h0210c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01087] =  I8a0037ad2845a3fbba9da380a8b8a576['h0210e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01088] =  I8a0037ad2845a3fbba9da380a8b8a576['h02110] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01089] =  I8a0037ad2845a3fbba9da380a8b8a576['h02112] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0108a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02114] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0108b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02116] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0108c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02118] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0108d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0211a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0108e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0211c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0108f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0211e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01090] =  I8a0037ad2845a3fbba9da380a8b8a576['h02120] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01091] =  I8a0037ad2845a3fbba9da380a8b8a576['h02122] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01092] =  I8a0037ad2845a3fbba9da380a8b8a576['h02124] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01093] =  I8a0037ad2845a3fbba9da380a8b8a576['h02126] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01094] =  I8a0037ad2845a3fbba9da380a8b8a576['h02128] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01095] =  I8a0037ad2845a3fbba9da380a8b8a576['h0212a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01096] =  I8a0037ad2845a3fbba9da380a8b8a576['h0212c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01097] =  I8a0037ad2845a3fbba9da380a8b8a576['h0212e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01098] =  I8a0037ad2845a3fbba9da380a8b8a576['h02130] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01099] =  I8a0037ad2845a3fbba9da380a8b8a576['h02132] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0109a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02134] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0109b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02136] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0109c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02138] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0109d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0213a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0109e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0213c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0109f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0213e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02140] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02142] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02144] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02146] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02148] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0214a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0214c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0214e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02150] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02152] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h02154] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h02156] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h02158] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0215a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0215c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010af] =  I8a0037ad2845a3fbba9da380a8b8a576['h0215e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02160] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02162] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02164] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02166] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02168] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0216a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0216c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0216e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02170] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02172] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h02174] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h02176] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h02178] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0217a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010be] =  I8a0037ad2845a3fbba9da380a8b8a576['h0217c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0217e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02180] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02182] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02184] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02186] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02188] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0218a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0218c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0218e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02190] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02192] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h02194] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h02196] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h02198] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0219a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0219c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0219e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h021a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h021a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h021a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h021a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h021a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h021aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h021ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h021ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h021b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h021b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010da] =  I8a0037ad2845a3fbba9da380a8b8a576['h021b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010db] =  I8a0037ad2845a3fbba9da380a8b8a576['h021b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h021b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h021ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010de] =  I8a0037ad2845a3fbba9da380a8b8a576['h021bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010df] =  I8a0037ad2845a3fbba9da380a8b8a576['h021be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h021c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h021c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h021c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h021c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h021c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h021ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h021cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h021ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h021d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h021d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h021d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h021d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h021d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h021da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h021dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h021de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h021e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h021e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h021e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h021e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h021e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h021ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h021ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h021ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h021f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h021f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h021f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h021f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h021f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h021fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h021fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h010ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h021fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01100] =  I8a0037ad2845a3fbba9da380a8b8a576['h02200] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01101] =  I8a0037ad2845a3fbba9da380a8b8a576['h02202] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01102] =  I8a0037ad2845a3fbba9da380a8b8a576['h02204] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01103] =  I8a0037ad2845a3fbba9da380a8b8a576['h02206] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01104] =  I8a0037ad2845a3fbba9da380a8b8a576['h02208] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01105] =  I8a0037ad2845a3fbba9da380a8b8a576['h0220a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01106] =  I8a0037ad2845a3fbba9da380a8b8a576['h0220c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01107] =  I8a0037ad2845a3fbba9da380a8b8a576['h0220e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01108] =  I8a0037ad2845a3fbba9da380a8b8a576['h02210] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01109] =  I8a0037ad2845a3fbba9da380a8b8a576['h02212] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0110a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02214] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0110b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02216] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0110c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02218] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0110d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0221a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0110e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0221c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0110f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0221e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01110] =  I8a0037ad2845a3fbba9da380a8b8a576['h02220] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01111] =  I8a0037ad2845a3fbba9da380a8b8a576['h02222] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01112] =  I8a0037ad2845a3fbba9da380a8b8a576['h02224] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01113] =  I8a0037ad2845a3fbba9da380a8b8a576['h02226] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01114] =  I8a0037ad2845a3fbba9da380a8b8a576['h02228] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01115] =  I8a0037ad2845a3fbba9da380a8b8a576['h0222a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01116] =  I8a0037ad2845a3fbba9da380a8b8a576['h0222c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01117] =  I8a0037ad2845a3fbba9da380a8b8a576['h0222e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01118] =  I8a0037ad2845a3fbba9da380a8b8a576['h02230] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01119] =  I8a0037ad2845a3fbba9da380a8b8a576['h02232] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0111a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02234] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0111b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02236] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0111c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02238] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0111d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0223a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0111e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0223c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0111f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0223e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01120] =  I8a0037ad2845a3fbba9da380a8b8a576['h02240] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01121] =  I8a0037ad2845a3fbba9da380a8b8a576['h02242] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01122] =  I8a0037ad2845a3fbba9da380a8b8a576['h02244] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01123] =  I8a0037ad2845a3fbba9da380a8b8a576['h02246] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01124] =  I8a0037ad2845a3fbba9da380a8b8a576['h02248] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01125] =  I8a0037ad2845a3fbba9da380a8b8a576['h0224a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01126] =  I8a0037ad2845a3fbba9da380a8b8a576['h0224c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01127] =  I8a0037ad2845a3fbba9da380a8b8a576['h0224e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01128] =  I8a0037ad2845a3fbba9da380a8b8a576['h02250] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01129] =  I8a0037ad2845a3fbba9da380a8b8a576['h02252] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0112a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02254] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0112b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02256] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0112c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02258] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0112d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0225a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0112e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0225c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0112f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0225e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01130] =  I8a0037ad2845a3fbba9da380a8b8a576['h02260] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01131] =  I8a0037ad2845a3fbba9da380a8b8a576['h02262] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01132] =  I8a0037ad2845a3fbba9da380a8b8a576['h02264] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01133] =  I8a0037ad2845a3fbba9da380a8b8a576['h02266] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01134] =  I8a0037ad2845a3fbba9da380a8b8a576['h02268] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01135] =  I8a0037ad2845a3fbba9da380a8b8a576['h0226a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01136] =  I8a0037ad2845a3fbba9da380a8b8a576['h0226c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01137] =  I8a0037ad2845a3fbba9da380a8b8a576['h0226e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01138] =  I8a0037ad2845a3fbba9da380a8b8a576['h02270] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01139] =  I8a0037ad2845a3fbba9da380a8b8a576['h02272] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0113a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02274] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0113b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02276] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0113c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02278] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0113d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0227a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0113e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0227c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0113f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0227e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01140] =  I8a0037ad2845a3fbba9da380a8b8a576['h02280] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01141] =  I8a0037ad2845a3fbba9da380a8b8a576['h02282] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01142] =  I8a0037ad2845a3fbba9da380a8b8a576['h02284] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01143] =  I8a0037ad2845a3fbba9da380a8b8a576['h02286] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01144] =  I8a0037ad2845a3fbba9da380a8b8a576['h02288] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01145] =  I8a0037ad2845a3fbba9da380a8b8a576['h0228a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01146] =  I8a0037ad2845a3fbba9da380a8b8a576['h0228c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01147] =  I8a0037ad2845a3fbba9da380a8b8a576['h0228e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01148] =  I8a0037ad2845a3fbba9da380a8b8a576['h02290] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01149] =  I8a0037ad2845a3fbba9da380a8b8a576['h02292] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0114a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02294] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0114b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02296] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0114c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02298] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0114d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0229a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0114e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0229c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0114f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0229e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01150] =  I8a0037ad2845a3fbba9da380a8b8a576['h022a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01151] =  I8a0037ad2845a3fbba9da380a8b8a576['h022a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01152] =  I8a0037ad2845a3fbba9da380a8b8a576['h022a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01153] =  I8a0037ad2845a3fbba9da380a8b8a576['h022a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01154] =  I8a0037ad2845a3fbba9da380a8b8a576['h022a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01155] =  I8a0037ad2845a3fbba9da380a8b8a576['h022aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01156] =  I8a0037ad2845a3fbba9da380a8b8a576['h022ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01157] =  I8a0037ad2845a3fbba9da380a8b8a576['h022ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01158] =  I8a0037ad2845a3fbba9da380a8b8a576['h022b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01159] =  I8a0037ad2845a3fbba9da380a8b8a576['h022b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0115a] =  I8a0037ad2845a3fbba9da380a8b8a576['h022b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0115b] =  I8a0037ad2845a3fbba9da380a8b8a576['h022b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0115c] =  I8a0037ad2845a3fbba9da380a8b8a576['h022b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0115d] =  I8a0037ad2845a3fbba9da380a8b8a576['h022ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0115e] =  I8a0037ad2845a3fbba9da380a8b8a576['h022bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0115f] =  I8a0037ad2845a3fbba9da380a8b8a576['h022be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01160] =  I8a0037ad2845a3fbba9da380a8b8a576['h022c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01161] =  I8a0037ad2845a3fbba9da380a8b8a576['h022c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01162] =  I8a0037ad2845a3fbba9da380a8b8a576['h022c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01163] =  I8a0037ad2845a3fbba9da380a8b8a576['h022c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01164] =  I8a0037ad2845a3fbba9da380a8b8a576['h022c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01165] =  I8a0037ad2845a3fbba9da380a8b8a576['h022ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01166] =  I8a0037ad2845a3fbba9da380a8b8a576['h022cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01167] =  I8a0037ad2845a3fbba9da380a8b8a576['h022ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01168] =  I8a0037ad2845a3fbba9da380a8b8a576['h022d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01169] =  I8a0037ad2845a3fbba9da380a8b8a576['h022d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0116a] =  I8a0037ad2845a3fbba9da380a8b8a576['h022d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0116b] =  I8a0037ad2845a3fbba9da380a8b8a576['h022d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0116c] =  I8a0037ad2845a3fbba9da380a8b8a576['h022d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0116d] =  I8a0037ad2845a3fbba9da380a8b8a576['h022da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0116e] =  I8a0037ad2845a3fbba9da380a8b8a576['h022dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0116f] =  I8a0037ad2845a3fbba9da380a8b8a576['h022de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01170] =  I8a0037ad2845a3fbba9da380a8b8a576['h022e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01171] =  I8a0037ad2845a3fbba9da380a8b8a576['h022e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01172] =  I8a0037ad2845a3fbba9da380a8b8a576['h022e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01173] =  I8a0037ad2845a3fbba9da380a8b8a576['h022e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01174] =  I8a0037ad2845a3fbba9da380a8b8a576['h022e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01175] =  I8a0037ad2845a3fbba9da380a8b8a576['h022ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01176] =  I8a0037ad2845a3fbba9da380a8b8a576['h022ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01177] =  I8a0037ad2845a3fbba9da380a8b8a576['h022ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01178] =  I8a0037ad2845a3fbba9da380a8b8a576['h022f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01179] =  I8a0037ad2845a3fbba9da380a8b8a576['h022f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0117a] =  I8a0037ad2845a3fbba9da380a8b8a576['h022f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0117b] =  I8a0037ad2845a3fbba9da380a8b8a576['h022f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0117c] =  I8a0037ad2845a3fbba9da380a8b8a576['h022f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0117d] =  I8a0037ad2845a3fbba9da380a8b8a576['h022fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0117e] =  I8a0037ad2845a3fbba9da380a8b8a576['h022fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0117f] =  I8a0037ad2845a3fbba9da380a8b8a576['h022fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01180] =  I8a0037ad2845a3fbba9da380a8b8a576['h02300] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01181] =  I8a0037ad2845a3fbba9da380a8b8a576['h02302] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01182] =  I8a0037ad2845a3fbba9da380a8b8a576['h02304] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01183] =  I8a0037ad2845a3fbba9da380a8b8a576['h02306] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01184] =  I8a0037ad2845a3fbba9da380a8b8a576['h02308] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01185] =  I8a0037ad2845a3fbba9da380a8b8a576['h0230a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01186] =  I8a0037ad2845a3fbba9da380a8b8a576['h0230c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01187] =  I8a0037ad2845a3fbba9da380a8b8a576['h0230e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01188] =  I8a0037ad2845a3fbba9da380a8b8a576['h02310] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01189] =  I8a0037ad2845a3fbba9da380a8b8a576['h02312] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0118a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02314] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0118b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02316] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0118c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02318] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0118d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0231a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0118e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0231c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0118f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0231e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01190] =  I8a0037ad2845a3fbba9da380a8b8a576['h02320] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01191] =  I8a0037ad2845a3fbba9da380a8b8a576['h02322] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01192] =  I8a0037ad2845a3fbba9da380a8b8a576['h02324] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01193] =  I8a0037ad2845a3fbba9da380a8b8a576['h02326] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01194] =  I8a0037ad2845a3fbba9da380a8b8a576['h02328] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01195] =  I8a0037ad2845a3fbba9da380a8b8a576['h0232a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01196] =  I8a0037ad2845a3fbba9da380a8b8a576['h0232c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01197] =  I8a0037ad2845a3fbba9da380a8b8a576['h0232e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01198] =  I8a0037ad2845a3fbba9da380a8b8a576['h02330] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01199] =  I8a0037ad2845a3fbba9da380a8b8a576['h02332] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0119a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02334] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0119b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02336] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0119c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02338] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0119d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0233a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0119e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0233c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0119f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0233e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02340] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02342] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02344] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02346] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02348] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0234a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0234c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0234e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02350] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02352] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h02354] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h02356] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h02358] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0235a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0235c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011af] =  I8a0037ad2845a3fbba9da380a8b8a576['h0235e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02360] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02362] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02364] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02366] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02368] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0236a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0236c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0236e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02370] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02372] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h02374] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h02376] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h02378] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0237a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011be] =  I8a0037ad2845a3fbba9da380a8b8a576['h0237c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0237e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02380] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02382] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02384] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02386] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02388] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0238a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0238c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0238e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02390] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02392] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h02394] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h02396] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h02398] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0239a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0239c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0239e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h023a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h023a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h023a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h023a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h023a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h023aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h023ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h023ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h023b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h023b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011da] =  I8a0037ad2845a3fbba9da380a8b8a576['h023b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011db] =  I8a0037ad2845a3fbba9da380a8b8a576['h023b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h023b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h023ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011de] =  I8a0037ad2845a3fbba9da380a8b8a576['h023bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011df] =  I8a0037ad2845a3fbba9da380a8b8a576['h023be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h023c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h023c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h023c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h023c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h023c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h023ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h023cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h023ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h023d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h023d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h023d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h023d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h023d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h023da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h023dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h023de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h023e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h023e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h023e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h023e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h023e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h023ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h023ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h023ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h023f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h023f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h023f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h023f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h023f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h023fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h023fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h011ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h023fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01200] =  I8a0037ad2845a3fbba9da380a8b8a576['h02400] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01201] =  I8a0037ad2845a3fbba9da380a8b8a576['h02402] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01202] =  I8a0037ad2845a3fbba9da380a8b8a576['h02404] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01203] =  I8a0037ad2845a3fbba9da380a8b8a576['h02406] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01204] =  I8a0037ad2845a3fbba9da380a8b8a576['h02408] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01205] =  I8a0037ad2845a3fbba9da380a8b8a576['h0240a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01206] =  I8a0037ad2845a3fbba9da380a8b8a576['h0240c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01207] =  I8a0037ad2845a3fbba9da380a8b8a576['h0240e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01208] =  I8a0037ad2845a3fbba9da380a8b8a576['h02410] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01209] =  I8a0037ad2845a3fbba9da380a8b8a576['h02412] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0120a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02414] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0120b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02416] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0120c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02418] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0120d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0241a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0120e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0241c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0120f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0241e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01210] =  I8a0037ad2845a3fbba9da380a8b8a576['h02420] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01211] =  I8a0037ad2845a3fbba9da380a8b8a576['h02422] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01212] =  I8a0037ad2845a3fbba9da380a8b8a576['h02424] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01213] =  I8a0037ad2845a3fbba9da380a8b8a576['h02426] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01214] =  I8a0037ad2845a3fbba9da380a8b8a576['h02428] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01215] =  I8a0037ad2845a3fbba9da380a8b8a576['h0242a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01216] =  I8a0037ad2845a3fbba9da380a8b8a576['h0242c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01217] =  I8a0037ad2845a3fbba9da380a8b8a576['h0242e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01218] =  I8a0037ad2845a3fbba9da380a8b8a576['h02430] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01219] =  I8a0037ad2845a3fbba9da380a8b8a576['h02432] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0121a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02434] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0121b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02436] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0121c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02438] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0121d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0243a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0121e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0243c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0121f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0243e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01220] =  I8a0037ad2845a3fbba9da380a8b8a576['h02440] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01221] =  I8a0037ad2845a3fbba9da380a8b8a576['h02442] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01222] =  I8a0037ad2845a3fbba9da380a8b8a576['h02444] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01223] =  I8a0037ad2845a3fbba9da380a8b8a576['h02446] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01224] =  I8a0037ad2845a3fbba9da380a8b8a576['h02448] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01225] =  I8a0037ad2845a3fbba9da380a8b8a576['h0244a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01226] =  I8a0037ad2845a3fbba9da380a8b8a576['h0244c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01227] =  I8a0037ad2845a3fbba9da380a8b8a576['h0244e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01228] =  I8a0037ad2845a3fbba9da380a8b8a576['h02450] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01229] =  I8a0037ad2845a3fbba9da380a8b8a576['h02452] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0122a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02454] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0122b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02456] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0122c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02458] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0122d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0245a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0122e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0245c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0122f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0245e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01230] =  I8a0037ad2845a3fbba9da380a8b8a576['h02460] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01231] =  I8a0037ad2845a3fbba9da380a8b8a576['h02462] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01232] =  I8a0037ad2845a3fbba9da380a8b8a576['h02464] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01233] =  I8a0037ad2845a3fbba9da380a8b8a576['h02466] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01234] =  I8a0037ad2845a3fbba9da380a8b8a576['h02468] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01235] =  I8a0037ad2845a3fbba9da380a8b8a576['h0246a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01236] =  I8a0037ad2845a3fbba9da380a8b8a576['h0246c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01237] =  I8a0037ad2845a3fbba9da380a8b8a576['h0246e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01238] =  I8a0037ad2845a3fbba9da380a8b8a576['h02470] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01239] =  I8a0037ad2845a3fbba9da380a8b8a576['h02472] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0123a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02474] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0123b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02476] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0123c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02478] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0123d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0247a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0123e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0247c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0123f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0247e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01240] =  I8a0037ad2845a3fbba9da380a8b8a576['h02480] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01241] =  I8a0037ad2845a3fbba9da380a8b8a576['h02482] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01242] =  I8a0037ad2845a3fbba9da380a8b8a576['h02484] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01243] =  I8a0037ad2845a3fbba9da380a8b8a576['h02486] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01244] =  I8a0037ad2845a3fbba9da380a8b8a576['h02488] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01245] =  I8a0037ad2845a3fbba9da380a8b8a576['h0248a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01246] =  I8a0037ad2845a3fbba9da380a8b8a576['h0248c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01247] =  I8a0037ad2845a3fbba9da380a8b8a576['h0248e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01248] =  I8a0037ad2845a3fbba9da380a8b8a576['h02490] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01249] =  I8a0037ad2845a3fbba9da380a8b8a576['h02492] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0124a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02494] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0124b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02496] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0124c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02498] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0124d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0249a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0124e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0249c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0124f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0249e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01250] =  I8a0037ad2845a3fbba9da380a8b8a576['h024a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01251] =  I8a0037ad2845a3fbba9da380a8b8a576['h024a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01252] =  I8a0037ad2845a3fbba9da380a8b8a576['h024a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01253] =  I8a0037ad2845a3fbba9da380a8b8a576['h024a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01254] =  I8a0037ad2845a3fbba9da380a8b8a576['h024a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01255] =  I8a0037ad2845a3fbba9da380a8b8a576['h024aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01256] =  I8a0037ad2845a3fbba9da380a8b8a576['h024ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01257] =  I8a0037ad2845a3fbba9da380a8b8a576['h024ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01258] =  I8a0037ad2845a3fbba9da380a8b8a576['h024b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01259] =  I8a0037ad2845a3fbba9da380a8b8a576['h024b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0125a] =  I8a0037ad2845a3fbba9da380a8b8a576['h024b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0125b] =  I8a0037ad2845a3fbba9da380a8b8a576['h024b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0125c] =  I8a0037ad2845a3fbba9da380a8b8a576['h024b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0125d] =  I8a0037ad2845a3fbba9da380a8b8a576['h024ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0125e] =  I8a0037ad2845a3fbba9da380a8b8a576['h024bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0125f] =  I8a0037ad2845a3fbba9da380a8b8a576['h024be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01260] =  I8a0037ad2845a3fbba9da380a8b8a576['h024c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01261] =  I8a0037ad2845a3fbba9da380a8b8a576['h024c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01262] =  I8a0037ad2845a3fbba9da380a8b8a576['h024c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01263] =  I8a0037ad2845a3fbba9da380a8b8a576['h024c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01264] =  I8a0037ad2845a3fbba9da380a8b8a576['h024c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01265] =  I8a0037ad2845a3fbba9da380a8b8a576['h024ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01266] =  I8a0037ad2845a3fbba9da380a8b8a576['h024cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01267] =  I8a0037ad2845a3fbba9da380a8b8a576['h024ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01268] =  I8a0037ad2845a3fbba9da380a8b8a576['h024d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01269] =  I8a0037ad2845a3fbba9da380a8b8a576['h024d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0126a] =  I8a0037ad2845a3fbba9da380a8b8a576['h024d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0126b] =  I8a0037ad2845a3fbba9da380a8b8a576['h024d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0126c] =  I8a0037ad2845a3fbba9da380a8b8a576['h024d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0126d] =  I8a0037ad2845a3fbba9da380a8b8a576['h024da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0126e] =  I8a0037ad2845a3fbba9da380a8b8a576['h024dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0126f] =  I8a0037ad2845a3fbba9da380a8b8a576['h024de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01270] =  I8a0037ad2845a3fbba9da380a8b8a576['h024e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01271] =  I8a0037ad2845a3fbba9da380a8b8a576['h024e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01272] =  I8a0037ad2845a3fbba9da380a8b8a576['h024e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01273] =  I8a0037ad2845a3fbba9da380a8b8a576['h024e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01274] =  I8a0037ad2845a3fbba9da380a8b8a576['h024e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01275] =  I8a0037ad2845a3fbba9da380a8b8a576['h024ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01276] =  I8a0037ad2845a3fbba9da380a8b8a576['h024ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01277] =  I8a0037ad2845a3fbba9da380a8b8a576['h024ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01278] =  I8a0037ad2845a3fbba9da380a8b8a576['h024f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01279] =  I8a0037ad2845a3fbba9da380a8b8a576['h024f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0127a] =  I8a0037ad2845a3fbba9da380a8b8a576['h024f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0127b] =  I8a0037ad2845a3fbba9da380a8b8a576['h024f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0127c] =  I8a0037ad2845a3fbba9da380a8b8a576['h024f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0127d] =  I8a0037ad2845a3fbba9da380a8b8a576['h024fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0127e] =  I8a0037ad2845a3fbba9da380a8b8a576['h024fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0127f] =  I8a0037ad2845a3fbba9da380a8b8a576['h024fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01280] =  I8a0037ad2845a3fbba9da380a8b8a576['h02500] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01281] =  I8a0037ad2845a3fbba9da380a8b8a576['h02502] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01282] =  I8a0037ad2845a3fbba9da380a8b8a576['h02504] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01283] =  I8a0037ad2845a3fbba9da380a8b8a576['h02506] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01284] =  I8a0037ad2845a3fbba9da380a8b8a576['h02508] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01285] =  I8a0037ad2845a3fbba9da380a8b8a576['h0250a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01286] =  I8a0037ad2845a3fbba9da380a8b8a576['h0250c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01287] =  I8a0037ad2845a3fbba9da380a8b8a576['h0250e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01288] =  I8a0037ad2845a3fbba9da380a8b8a576['h02510] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01289] =  I8a0037ad2845a3fbba9da380a8b8a576['h02512] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0128a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02514] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0128b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02516] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0128c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02518] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0128d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0251a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0128e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0251c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0128f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0251e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01290] =  I8a0037ad2845a3fbba9da380a8b8a576['h02520] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01291] =  I8a0037ad2845a3fbba9da380a8b8a576['h02522] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01292] =  I8a0037ad2845a3fbba9da380a8b8a576['h02524] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01293] =  I8a0037ad2845a3fbba9da380a8b8a576['h02526] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01294] =  I8a0037ad2845a3fbba9da380a8b8a576['h02528] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01295] =  I8a0037ad2845a3fbba9da380a8b8a576['h0252a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01296] =  I8a0037ad2845a3fbba9da380a8b8a576['h0252c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01297] =  I8a0037ad2845a3fbba9da380a8b8a576['h0252e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01298] =  I8a0037ad2845a3fbba9da380a8b8a576['h02530] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01299] =  I8a0037ad2845a3fbba9da380a8b8a576['h02532] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0129a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02534] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0129b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02536] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0129c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02538] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0129d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0253a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0129e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0253c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0129f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0253e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02540] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02542] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02544] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02546] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02548] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0254a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0254c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0254e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02550] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02552] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h02554] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h02556] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h02558] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0255a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0255c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012af] =  I8a0037ad2845a3fbba9da380a8b8a576['h0255e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02560] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02562] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02564] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02566] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02568] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0256a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0256c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0256e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02570] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02572] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h02574] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h02576] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h02578] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0257a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012be] =  I8a0037ad2845a3fbba9da380a8b8a576['h0257c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0257e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02580] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02582] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02584] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02586] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02588] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0258a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0258c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0258e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02590] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02592] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h02594] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h02596] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h02598] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0259a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0259c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0259e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h025a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h025a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h025a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h025a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h025a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h025aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h025ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h025ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h025b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h025b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012da] =  I8a0037ad2845a3fbba9da380a8b8a576['h025b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012db] =  I8a0037ad2845a3fbba9da380a8b8a576['h025b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h025b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h025ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012de] =  I8a0037ad2845a3fbba9da380a8b8a576['h025bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012df] =  I8a0037ad2845a3fbba9da380a8b8a576['h025be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h025c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h025c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h025c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h025c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h025c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h025ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h025cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h025ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h025d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h025d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h025d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h025d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h025d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h025da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h025dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h025de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h025e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h025e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h025e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h025e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h025e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h025ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h025ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h025ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h025f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h025f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h025f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h025f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h025f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h025fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h025fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h012ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h025fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01300] =  I8a0037ad2845a3fbba9da380a8b8a576['h02600] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01301] =  I8a0037ad2845a3fbba9da380a8b8a576['h02602] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01302] =  I8a0037ad2845a3fbba9da380a8b8a576['h02604] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01303] =  I8a0037ad2845a3fbba9da380a8b8a576['h02606] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01304] =  I8a0037ad2845a3fbba9da380a8b8a576['h02608] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01305] =  I8a0037ad2845a3fbba9da380a8b8a576['h0260a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01306] =  I8a0037ad2845a3fbba9da380a8b8a576['h0260c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01307] =  I8a0037ad2845a3fbba9da380a8b8a576['h0260e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01308] =  I8a0037ad2845a3fbba9da380a8b8a576['h02610] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01309] =  I8a0037ad2845a3fbba9da380a8b8a576['h02612] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0130a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02614] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0130b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02616] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0130c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02618] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0130d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0261a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0130e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0261c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0130f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0261e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01310] =  I8a0037ad2845a3fbba9da380a8b8a576['h02620] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01311] =  I8a0037ad2845a3fbba9da380a8b8a576['h02622] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01312] =  I8a0037ad2845a3fbba9da380a8b8a576['h02624] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01313] =  I8a0037ad2845a3fbba9da380a8b8a576['h02626] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01314] =  I8a0037ad2845a3fbba9da380a8b8a576['h02628] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01315] =  I8a0037ad2845a3fbba9da380a8b8a576['h0262a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01316] =  I8a0037ad2845a3fbba9da380a8b8a576['h0262c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01317] =  I8a0037ad2845a3fbba9da380a8b8a576['h0262e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01318] =  I8a0037ad2845a3fbba9da380a8b8a576['h02630] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01319] =  I8a0037ad2845a3fbba9da380a8b8a576['h02632] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0131a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02634] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0131b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02636] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0131c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02638] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0131d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0263a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0131e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0263c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0131f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0263e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01320] =  I8a0037ad2845a3fbba9da380a8b8a576['h02640] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01321] =  I8a0037ad2845a3fbba9da380a8b8a576['h02642] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01322] =  I8a0037ad2845a3fbba9da380a8b8a576['h02644] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01323] =  I8a0037ad2845a3fbba9da380a8b8a576['h02646] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01324] =  I8a0037ad2845a3fbba9da380a8b8a576['h02648] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01325] =  I8a0037ad2845a3fbba9da380a8b8a576['h0264a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01326] =  I8a0037ad2845a3fbba9da380a8b8a576['h0264c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01327] =  I8a0037ad2845a3fbba9da380a8b8a576['h0264e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01328] =  I8a0037ad2845a3fbba9da380a8b8a576['h02650] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01329] =  I8a0037ad2845a3fbba9da380a8b8a576['h02652] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0132a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02654] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0132b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02656] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0132c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02658] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0132d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0265a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0132e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0265c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0132f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0265e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01330] =  I8a0037ad2845a3fbba9da380a8b8a576['h02660] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01331] =  I8a0037ad2845a3fbba9da380a8b8a576['h02662] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01332] =  I8a0037ad2845a3fbba9da380a8b8a576['h02664] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01333] =  I8a0037ad2845a3fbba9da380a8b8a576['h02666] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01334] =  I8a0037ad2845a3fbba9da380a8b8a576['h02668] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01335] =  I8a0037ad2845a3fbba9da380a8b8a576['h0266a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01336] =  I8a0037ad2845a3fbba9da380a8b8a576['h0266c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01337] =  I8a0037ad2845a3fbba9da380a8b8a576['h0266e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01338] =  I8a0037ad2845a3fbba9da380a8b8a576['h02670] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01339] =  I8a0037ad2845a3fbba9da380a8b8a576['h02672] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0133a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02674] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0133b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02676] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0133c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02678] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0133d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0267a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0133e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0267c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0133f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0267e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01340] =  I8a0037ad2845a3fbba9da380a8b8a576['h02680] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01341] =  I8a0037ad2845a3fbba9da380a8b8a576['h02682] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01342] =  I8a0037ad2845a3fbba9da380a8b8a576['h02684] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01343] =  I8a0037ad2845a3fbba9da380a8b8a576['h02686] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01344] =  I8a0037ad2845a3fbba9da380a8b8a576['h02688] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01345] =  I8a0037ad2845a3fbba9da380a8b8a576['h0268a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01346] =  I8a0037ad2845a3fbba9da380a8b8a576['h0268c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01347] =  I8a0037ad2845a3fbba9da380a8b8a576['h0268e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01348] =  I8a0037ad2845a3fbba9da380a8b8a576['h02690] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01349] =  I8a0037ad2845a3fbba9da380a8b8a576['h02692] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0134a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02694] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0134b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02696] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0134c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02698] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0134d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0269a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0134e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0269c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0134f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0269e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01350] =  I8a0037ad2845a3fbba9da380a8b8a576['h026a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01351] =  I8a0037ad2845a3fbba9da380a8b8a576['h026a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01352] =  I8a0037ad2845a3fbba9da380a8b8a576['h026a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01353] =  I8a0037ad2845a3fbba9da380a8b8a576['h026a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01354] =  I8a0037ad2845a3fbba9da380a8b8a576['h026a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01355] =  I8a0037ad2845a3fbba9da380a8b8a576['h026aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01356] =  I8a0037ad2845a3fbba9da380a8b8a576['h026ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01357] =  I8a0037ad2845a3fbba9da380a8b8a576['h026ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01358] =  I8a0037ad2845a3fbba9da380a8b8a576['h026b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01359] =  I8a0037ad2845a3fbba9da380a8b8a576['h026b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0135a] =  I8a0037ad2845a3fbba9da380a8b8a576['h026b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0135b] =  I8a0037ad2845a3fbba9da380a8b8a576['h026b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0135c] =  I8a0037ad2845a3fbba9da380a8b8a576['h026b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0135d] =  I8a0037ad2845a3fbba9da380a8b8a576['h026ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0135e] =  I8a0037ad2845a3fbba9da380a8b8a576['h026bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0135f] =  I8a0037ad2845a3fbba9da380a8b8a576['h026be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01360] =  I8a0037ad2845a3fbba9da380a8b8a576['h026c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01361] =  I8a0037ad2845a3fbba9da380a8b8a576['h026c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01362] =  I8a0037ad2845a3fbba9da380a8b8a576['h026c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01363] =  I8a0037ad2845a3fbba9da380a8b8a576['h026c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01364] =  I8a0037ad2845a3fbba9da380a8b8a576['h026c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01365] =  I8a0037ad2845a3fbba9da380a8b8a576['h026ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01366] =  I8a0037ad2845a3fbba9da380a8b8a576['h026cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01367] =  I8a0037ad2845a3fbba9da380a8b8a576['h026ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01368] =  I8a0037ad2845a3fbba9da380a8b8a576['h026d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01369] =  I8a0037ad2845a3fbba9da380a8b8a576['h026d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0136a] =  I8a0037ad2845a3fbba9da380a8b8a576['h026d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0136b] =  I8a0037ad2845a3fbba9da380a8b8a576['h026d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0136c] =  I8a0037ad2845a3fbba9da380a8b8a576['h026d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0136d] =  I8a0037ad2845a3fbba9da380a8b8a576['h026da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0136e] =  I8a0037ad2845a3fbba9da380a8b8a576['h026dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0136f] =  I8a0037ad2845a3fbba9da380a8b8a576['h026de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01370] =  I8a0037ad2845a3fbba9da380a8b8a576['h026e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01371] =  I8a0037ad2845a3fbba9da380a8b8a576['h026e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01372] =  I8a0037ad2845a3fbba9da380a8b8a576['h026e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01373] =  I8a0037ad2845a3fbba9da380a8b8a576['h026e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01374] =  I8a0037ad2845a3fbba9da380a8b8a576['h026e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01375] =  I8a0037ad2845a3fbba9da380a8b8a576['h026ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01376] =  I8a0037ad2845a3fbba9da380a8b8a576['h026ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01377] =  I8a0037ad2845a3fbba9da380a8b8a576['h026ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01378] =  I8a0037ad2845a3fbba9da380a8b8a576['h026f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01379] =  I8a0037ad2845a3fbba9da380a8b8a576['h026f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0137a] =  I8a0037ad2845a3fbba9da380a8b8a576['h026f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0137b] =  I8a0037ad2845a3fbba9da380a8b8a576['h026f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0137c] =  I8a0037ad2845a3fbba9da380a8b8a576['h026f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0137d] =  I8a0037ad2845a3fbba9da380a8b8a576['h026fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0137e] =  I8a0037ad2845a3fbba9da380a8b8a576['h026fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0137f] =  I8a0037ad2845a3fbba9da380a8b8a576['h026fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01380] =  I8a0037ad2845a3fbba9da380a8b8a576['h02700] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01381] =  I8a0037ad2845a3fbba9da380a8b8a576['h02702] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01382] =  I8a0037ad2845a3fbba9da380a8b8a576['h02704] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01383] =  I8a0037ad2845a3fbba9da380a8b8a576['h02706] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01384] =  I8a0037ad2845a3fbba9da380a8b8a576['h02708] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01385] =  I8a0037ad2845a3fbba9da380a8b8a576['h0270a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01386] =  I8a0037ad2845a3fbba9da380a8b8a576['h0270c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01387] =  I8a0037ad2845a3fbba9da380a8b8a576['h0270e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01388] =  I8a0037ad2845a3fbba9da380a8b8a576['h02710] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01389] =  I8a0037ad2845a3fbba9da380a8b8a576['h02712] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0138a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02714] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0138b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02716] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0138c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02718] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0138d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0271a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0138e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0271c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0138f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0271e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01390] =  I8a0037ad2845a3fbba9da380a8b8a576['h02720] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01391] =  I8a0037ad2845a3fbba9da380a8b8a576['h02722] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01392] =  I8a0037ad2845a3fbba9da380a8b8a576['h02724] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01393] =  I8a0037ad2845a3fbba9da380a8b8a576['h02726] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01394] =  I8a0037ad2845a3fbba9da380a8b8a576['h02728] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01395] =  I8a0037ad2845a3fbba9da380a8b8a576['h0272a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01396] =  I8a0037ad2845a3fbba9da380a8b8a576['h0272c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01397] =  I8a0037ad2845a3fbba9da380a8b8a576['h0272e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01398] =  I8a0037ad2845a3fbba9da380a8b8a576['h02730] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01399] =  I8a0037ad2845a3fbba9da380a8b8a576['h02732] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0139a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02734] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0139b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02736] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0139c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02738] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0139d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0273a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0139e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0273c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0139f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0273e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02740] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02742] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02744] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02746] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02748] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0274a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0274c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0274e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02750] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02752] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h02754] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h02756] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h02758] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0275a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0275c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013af] =  I8a0037ad2845a3fbba9da380a8b8a576['h0275e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02760] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02762] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02764] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02766] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02768] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0276a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0276c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0276e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02770] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02772] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h02774] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h02776] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h02778] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0277a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013be] =  I8a0037ad2845a3fbba9da380a8b8a576['h0277c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0277e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02780] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02782] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02784] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02786] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02788] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0278a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0278c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0278e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02790] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02792] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h02794] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h02796] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h02798] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0279a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0279c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0279e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h027a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h027a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h027a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h027a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h027a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h027aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h027ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h027ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h027b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h027b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013da] =  I8a0037ad2845a3fbba9da380a8b8a576['h027b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013db] =  I8a0037ad2845a3fbba9da380a8b8a576['h027b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h027b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h027ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013de] =  I8a0037ad2845a3fbba9da380a8b8a576['h027bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013df] =  I8a0037ad2845a3fbba9da380a8b8a576['h027be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h027c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h027c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h027c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h027c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h027c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h027ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h027cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h027ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h027d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h027d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h027d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h027d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h027d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h027da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h027dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h027de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h027e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h027e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h027e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h027e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h027e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h027ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h027ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h027ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h027f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h027f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h027f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h027f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h027f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h027fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h027fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h013ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h027fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01400] =  I8a0037ad2845a3fbba9da380a8b8a576['h02800] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01401] =  I8a0037ad2845a3fbba9da380a8b8a576['h02802] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01402] =  I8a0037ad2845a3fbba9da380a8b8a576['h02804] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01403] =  I8a0037ad2845a3fbba9da380a8b8a576['h02806] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01404] =  I8a0037ad2845a3fbba9da380a8b8a576['h02808] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01405] =  I8a0037ad2845a3fbba9da380a8b8a576['h0280a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01406] =  I8a0037ad2845a3fbba9da380a8b8a576['h0280c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01407] =  I8a0037ad2845a3fbba9da380a8b8a576['h0280e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01408] =  I8a0037ad2845a3fbba9da380a8b8a576['h02810] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01409] =  I8a0037ad2845a3fbba9da380a8b8a576['h02812] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0140a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02814] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0140b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02816] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0140c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02818] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0140d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0281a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0140e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0281c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0140f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0281e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01410] =  I8a0037ad2845a3fbba9da380a8b8a576['h02820] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01411] =  I8a0037ad2845a3fbba9da380a8b8a576['h02822] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01412] =  I8a0037ad2845a3fbba9da380a8b8a576['h02824] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01413] =  I8a0037ad2845a3fbba9da380a8b8a576['h02826] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01414] =  I8a0037ad2845a3fbba9da380a8b8a576['h02828] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01415] =  I8a0037ad2845a3fbba9da380a8b8a576['h0282a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01416] =  I8a0037ad2845a3fbba9da380a8b8a576['h0282c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01417] =  I8a0037ad2845a3fbba9da380a8b8a576['h0282e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01418] =  I8a0037ad2845a3fbba9da380a8b8a576['h02830] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01419] =  I8a0037ad2845a3fbba9da380a8b8a576['h02832] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0141a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02834] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0141b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02836] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0141c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02838] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0141d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0283a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0141e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0283c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0141f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0283e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01420] =  I8a0037ad2845a3fbba9da380a8b8a576['h02840] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01421] =  I8a0037ad2845a3fbba9da380a8b8a576['h02842] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01422] =  I8a0037ad2845a3fbba9da380a8b8a576['h02844] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01423] =  I8a0037ad2845a3fbba9da380a8b8a576['h02846] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01424] =  I8a0037ad2845a3fbba9da380a8b8a576['h02848] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01425] =  I8a0037ad2845a3fbba9da380a8b8a576['h0284a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01426] =  I8a0037ad2845a3fbba9da380a8b8a576['h0284c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01427] =  I8a0037ad2845a3fbba9da380a8b8a576['h0284e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01428] =  I8a0037ad2845a3fbba9da380a8b8a576['h02850] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01429] =  I8a0037ad2845a3fbba9da380a8b8a576['h02852] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0142a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02854] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0142b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02856] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0142c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02858] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0142d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0285a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0142e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0285c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0142f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0285e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01430] =  I8a0037ad2845a3fbba9da380a8b8a576['h02860] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01431] =  I8a0037ad2845a3fbba9da380a8b8a576['h02862] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01432] =  I8a0037ad2845a3fbba9da380a8b8a576['h02864] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01433] =  I8a0037ad2845a3fbba9da380a8b8a576['h02866] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01434] =  I8a0037ad2845a3fbba9da380a8b8a576['h02868] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01435] =  I8a0037ad2845a3fbba9da380a8b8a576['h0286a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01436] =  I8a0037ad2845a3fbba9da380a8b8a576['h0286c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01437] =  I8a0037ad2845a3fbba9da380a8b8a576['h0286e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01438] =  I8a0037ad2845a3fbba9da380a8b8a576['h02870] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01439] =  I8a0037ad2845a3fbba9da380a8b8a576['h02872] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0143a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02874] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0143b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02876] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0143c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02878] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0143d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0287a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0143e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0287c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0143f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0287e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01440] =  I8a0037ad2845a3fbba9da380a8b8a576['h02880] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01441] =  I8a0037ad2845a3fbba9da380a8b8a576['h02882] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01442] =  I8a0037ad2845a3fbba9da380a8b8a576['h02884] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01443] =  I8a0037ad2845a3fbba9da380a8b8a576['h02886] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01444] =  I8a0037ad2845a3fbba9da380a8b8a576['h02888] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01445] =  I8a0037ad2845a3fbba9da380a8b8a576['h0288a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01446] =  I8a0037ad2845a3fbba9da380a8b8a576['h0288c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01447] =  I8a0037ad2845a3fbba9da380a8b8a576['h0288e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01448] =  I8a0037ad2845a3fbba9da380a8b8a576['h02890] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01449] =  I8a0037ad2845a3fbba9da380a8b8a576['h02892] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0144a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02894] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0144b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02896] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0144c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02898] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0144d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0289a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0144e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0289c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0144f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0289e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01450] =  I8a0037ad2845a3fbba9da380a8b8a576['h028a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01451] =  I8a0037ad2845a3fbba9da380a8b8a576['h028a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01452] =  I8a0037ad2845a3fbba9da380a8b8a576['h028a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01453] =  I8a0037ad2845a3fbba9da380a8b8a576['h028a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01454] =  I8a0037ad2845a3fbba9da380a8b8a576['h028a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01455] =  I8a0037ad2845a3fbba9da380a8b8a576['h028aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01456] =  I8a0037ad2845a3fbba9da380a8b8a576['h028ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01457] =  I8a0037ad2845a3fbba9da380a8b8a576['h028ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01458] =  I8a0037ad2845a3fbba9da380a8b8a576['h028b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01459] =  I8a0037ad2845a3fbba9da380a8b8a576['h028b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0145a] =  I8a0037ad2845a3fbba9da380a8b8a576['h028b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0145b] =  I8a0037ad2845a3fbba9da380a8b8a576['h028b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0145c] =  I8a0037ad2845a3fbba9da380a8b8a576['h028b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0145d] =  I8a0037ad2845a3fbba9da380a8b8a576['h028ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0145e] =  I8a0037ad2845a3fbba9da380a8b8a576['h028bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0145f] =  I8a0037ad2845a3fbba9da380a8b8a576['h028be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01460] =  I8a0037ad2845a3fbba9da380a8b8a576['h028c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01461] =  I8a0037ad2845a3fbba9da380a8b8a576['h028c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01462] =  I8a0037ad2845a3fbba9da380a8b8a576['h028c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01463] =  I8a0037ad2845a3fbba9da380a8b8a576['h028c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01464] =  I8a0037ad2845a3fbba9da380a8b8a576['h028c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01465] =  I8a0037ad2845a3fbba9da380a8b8a576['h028ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01466] =  I8a0037ad2845a3fbba9da380a8b8a576['h028cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01467] =  I8a0037ad2845a3fbba9da380a8b8a576['h028ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01468] =  I8a0037ad2845a3fbba9da380a8b8a576['h028d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01469] =  I8a0037ad2845a3fbba9da380a8b8a576['h028d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0146a] =  I8a0037ad2845a3fbba9da380a8b8a576['h028d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0146b] =  I8a0037ad2845a3fbba9da380a8b8a576['h028d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0146c] =  I8a0037ad2845a3fbba9da380a8b8a576['h028d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0146d] =  I8a0037ad2845a3fbba9da380a8b8a576['h028da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0146e] =  I8a0037ad2845a3fbba9da380a8b8a576['h028dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0146f] =  I8a0037ad2845a3fbba9da380a8b8a576['h028de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01470] =  I8a0037ad2845a3fbba9da380a8b8a576['h028e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01471] =  I8a0037ad2845a3fbba9da380a8b8a576['h028e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01472] =  I8a0037ad2845a3fbba9da380a8b8a576['h028e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01473] =  I8a0037ad2845a3fbba9da380a8b8a576['h028e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01474] =  I8a0037ad2845a3fbba9da380a8b8a576['h028e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01475] =  I8a0037ad2845a3fbba9da380a8b8a576['h028ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01476] =  I8a0037ad2845a3fbba9da380a8b8a576['h028ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01477] =  I8a0037ad2845a3fbba9da380a8b8a576['h028ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01478] =  I8a0037ad2845a3fbba9da380a8b8a576['h028f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01479] =  I8a0037ad2845a3fbba9da380a8b8a576['h028f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0147a] =  I8a0037ad2845a3fbba9da380a8b8a576['h028f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0147b] =  I8a0037ad2845a3fbba9da380a8b8a576['h028f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0147c] =  I8a0037ad2845a3fbba9da380a8b8a576['h028f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0147d] =  I8a0037ad2845a3fbba9da380a8b8a576['h028fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0147e] =  I8a0037ad2845a3fbba9da380a8b8a576['h028fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0147f] =  I8a0037ad2845a3fbba9da380a8b8a576['h028fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01480] =  I8a0037ad2845a3fbba9da380a8b8a576['h02900] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01481] =  I8a0037ad2845a3fbba9da380a8b8a576['h02902] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01482] =  I8a0037ad2845a3fbba9da380a8b8a576['h02904] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01483] =  I8a0037ad2845a3fbba9da380a8b8a576['h02906] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01484] =  I8a0037ad2845a3fbba9da380a8b8a576['h02908] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01485] =  I8a0037ad2845a3fbba9da380a8b8a576['h0290a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01486] =  I8a0037ad2845a3fbba9da380a8b8a576['h0290c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01487] =  I8a0037ad2845a3fbba9da380a8b8a576['h0290e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01488] =  I8a0037ad2845a3fbba9da380a8b8a576['h02910] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01489] =  I8a0037ad2845a3fbba9da380a8b8a576['h02912] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0148a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02914] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0148b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02916] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0148c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02918] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0148d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0291a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0148e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0291c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0148f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0291e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01490] =  I8a0037ad2845a3fbba9da380a8b8a576['h02920] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01491] =  I8a0037ad2845a3fbba9da380a8b8a576['h02922] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01492] =  I8a0037ad2845a3fbba9da380a8b8a576['h02924] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01493] =  I8a0037ad2845a3fbba9da380a8b8a576['h02926] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01494] =  I8a0037ad2845a3fbba9da380a8b8a576['h02928] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01495] =  I8a0037ad2845a3fbba9da380a8b8a576['h0292a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01496] =  I8a0037ad2845a3fbba9da380a8b8a576['h0292c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01497] =  I8a0037ad2845a3fbba9da380a8b8a576['h0292e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01498] =  I8a0037ad2845a3fbba9da380a8b8a576['h02930] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01499] =  I8a0037ad2845a3fbba9da380a8b8a576['h02932] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0149a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02934] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0149b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02936] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0149c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02938] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0149d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0293a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0149e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0293c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0149f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0293e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02940] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02942] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02944] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02946] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02948] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0294a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0294c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0294e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02950] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02952] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h02954] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h02956] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h02958] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0295a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0295c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014af] =  I8a0037ad2845a3fbba9da380a8b8a576['h0295e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02960] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02962] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02964] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02966] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02968] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0296a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0296c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0296e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02970] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02972] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h02974] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h02976] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h02978] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0297a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014be] =  I8a0037ad2845a3fbba9da380a8b8a576['h0297c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0297e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02980] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02982] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02984] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02986] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02988] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0298a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0298c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0298e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02990] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02992] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h02994] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h02996] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h02998] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0299a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0299c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0299e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h029a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h029a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h029a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h029a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h029a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h029aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h029ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h029ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h029b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h029b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014da] =  I8a0037ad2845a3fbba9da380a8b8a576['h029b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014db] =  I8a0037ad2845a3fbba9da380a8b8a576['h029b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h029b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h029ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014de] =  I8a0037ad2845a3fbba9da380a8b8a576['h029bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014df] =  I8a0037ad2845a3fbba9da380a8b8a576['h029be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h029c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h029c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h029c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h029c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h029c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h029ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h029cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h029ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h029d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h029d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h029d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h029d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h029d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h029da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h029dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h029de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h029e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h029e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h029e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h029e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h029e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h029ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h029ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h029ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h029f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h029f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h029f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h029f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h029f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h029fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h029fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h014ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h029fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01500] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01501] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01502] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01503] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01504] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01505] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01506] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01507] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01508] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01509] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0150a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0150b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0150c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0150d] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0150e] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0150f] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01510] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01511] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01512] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01513] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01514] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01515] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01516] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01517] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01518] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01519] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0151a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0151b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0151c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0151d] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0151e] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0151f] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01520] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01521] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01522] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01523] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01524] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01525] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01526] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01527] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01528] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01529] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0152a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0152b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0152c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0152d] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0152e] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0152f] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01530] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01531] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01532] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01533] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01534] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01535] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01536] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01537] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01538] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01539] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0153a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0153b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0153c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0153d] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0153e] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0153f] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01540] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01541] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01542] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01543] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01544] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01545] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01546] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01547] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01548] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01549] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0154a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0154b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0154c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0154d] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0154e] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0154f] =  I8a0037ad2845a3fbba9da380a8b8a576['h02a9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01550] =  I8a0037ad2845a3fbba9da380a8b8a576['h02aa0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01551] =  I8a0037ad2845a3fbba9da380a8b8a576['h02aa2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01552] =  I8a0037ad2845a3fbba9da380a8b8a576['h02aa4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01553] =  I8a0037ad2845a3fbba9da380a8b8a576['h02aa6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01554] =  I8a0037ad2845a3fbba9da380a8b8a576['h02aa8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01555] =  I8a0037ad2845a3fbba9da380a8b8a576['h02aaa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01556] =  I8a0037ad2845a3fbba9da380a8b8a576['h02aac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01557] =  I8a0037ad2845a3fbba9da380a8b8a576['h02aae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01558] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ab0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01559] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ab2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0155a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ab4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0155b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ab6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0155c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ab8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0155d] =  I8a0037ad2845a3fbba9da380a8b8a576['h02aba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0155e] =  I8a0037ad2845a3fbba9da380a8b8a576['h02abc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0155f] =  I8a0037ad2845a3fbba9da380a8b8a576['h02abe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01560] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ac0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01561] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ac2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01562] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ac4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01563] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ac6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01564] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ac8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01565] =  I8a0037ad2845a3fbba9da380a8b8a576['h02aca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01566] =  I8a0037ad2845a3fbba9da380a8b8a576['h02acc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01567] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ace] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01568] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ad0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01569] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ad2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0156a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ad4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0156b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ad6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0156c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ad8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0156d] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ada] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0156e] =  I8a0037ad2845a3fbba9da380a8b8a576['h02adc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0156f] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ade] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01570] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ae0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01571] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ae2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01572] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ae4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01573] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ae6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01574] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ae8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01575] =  I8a0037ad2845a3fbba9da380a8b8a576['h02aea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01576] =  I8a0037ad2845a3fbba9da380a8b8a576['h02aec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01577] =  I8a0037ad2845a3fbba9da380a8b8a576['h02aee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01578] =  I8a0037ad2845a3fbba9da380a8b8a576['h02af0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01579] =  I8a0037ad2845a3fbba9da380a8b8a576['h02af2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0157a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02af4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0157b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02af6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0157c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02af8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0157d] =  I8a0037ad2845a3fbba9da380a8b8a576['h02afa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0157e] =  I8a0037ad2845a3fbba9da380a8b8a576['h02afc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0157f] =  I8a0037ad2845a3fbba9da380a8b8a576['h02afe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01580] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01581] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01582] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01583] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01584] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01585] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01586] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01587] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01588] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01589] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0158a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0158b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0158c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0158d] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0158e] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0158f] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01590] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01591] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01592] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01593] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01594] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01595] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01596] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01597] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01598] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01599] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0159a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0159b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0159c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0159d] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0159e] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0159f] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015af] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015be] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h02b9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ba0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ba2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ba4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ba6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ba8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h02baa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015da] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015db] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015de] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015df] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bcc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bdc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02be0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02be2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02be4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02be6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02be8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bf0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bf2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bf4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bf6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bf8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bfa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bfc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h015ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h02bfe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01600] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01601] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01602] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01603] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01604] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01605] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01606] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01607] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01608] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01609] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0160a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0160b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0160c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0160d] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0160e] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0160f] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01610] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01611] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01612] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01613] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01614] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01615] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01616] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01617] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01618] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01619] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0161a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0161b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0161c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0161d] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0161e] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0161f] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01620] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01621] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01622] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01623] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01624] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01625] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01626] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01627] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01628] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01629] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0162a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0162b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0162c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0162d] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0162e] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0162f] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01630] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01631] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01632] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01633] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01634] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01635] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01636] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01637] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01638] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01639] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0163a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0163b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0163c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0163d] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0163e] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0163f] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01640] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01641] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01642] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01643] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01644] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01645] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01646] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01647] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01648] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01649] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0164a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0164b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0164c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0164d] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0164e] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0164f] =  I8a0037ad2845a3fbba9da380a8b8a576['h02c9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01650] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ca0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01651] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ca2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01652] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ca4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01653] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ca6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01654] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ca8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01655] =  I8a0037ad2845a3fbba9da380a8b8a576['h02caa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01656] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01657] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01658] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01659] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0165a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0165b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0165c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0165d] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0165e] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0165f] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01660] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01661] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01662] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01663] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01664] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01665] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01666] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ccc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01667] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01668] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01669] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0166a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0166b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0166c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0166d] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0166e] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cdc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0166f] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01670] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ce0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01671] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ce2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01672] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ce4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01673] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ce6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01674] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ce8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01675] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01676] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01677] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01678] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cf0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01679] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cf2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0167a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cf4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0167b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cf6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0167c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cf8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0167d] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cfa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0167e] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cfc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0167f] =  I8a0037ad2845a3fbba9da380a8b8a576['h02cfe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01680] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01681] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01682] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01683] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01684] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01685] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01686] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01687] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01688] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01689] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0168a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0168b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0168c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0168d] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0168e] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0168f] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01690] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01691] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01692] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01693] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01694] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01695] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01696] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01697] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01698] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01699] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0169a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0169b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0169c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0169d] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0169e] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0169f] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016af] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016be] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h02d9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02da0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02da2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02da4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02da6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02da8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h02daa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h02dac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h02dae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02db0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02db2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016da] =  I8a0037ad2845a3fbba9da380a8b8a576['h02db4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016db] =  I8a0037ad2845a3fbba9da380a8b8a576['h02db6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h02db8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h02dba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016de] =  I8a0037ad2845a3fbba9da380a8b8a576['h02dbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016df] =  I8a0037ad2845a3fbba9da380a8b8a576['h02dbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02dc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02dc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02dc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02dc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02dc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h02dca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h02dcc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h02dce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02dd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02dd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h02dd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h02dd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h02dd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h02dda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ddc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h02dde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02de0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02de2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02de4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02de6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02de8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h02dea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h02dec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h02dee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02df0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02df2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h02df4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h02df6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h02df8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h02dfa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h02dfc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h016ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h02dfe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01700] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01701] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01702] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01703] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01704] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01705] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01706] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01707] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01708] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01709] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0170a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0170b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0170c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0170d] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0170e] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0170f] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01710] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01711] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01712] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01713] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01714] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01715] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01716] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01717] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01718] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01719] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0171a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0171b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0171c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0171d] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0171e] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0171f] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01720] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01721] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01722] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01723] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01724] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01725] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01726] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01727] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01728] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01729] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0172a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0172b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0172c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0172d] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0172e] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0172f] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01730] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01731] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01732] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01733] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01734] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01735] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01736] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01737] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01738] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01739] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0173a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0173b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0173c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0173d] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0173e] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0173f] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01740] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01741] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01742] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01743] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01744] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01745] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01746] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01747] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01748] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01749] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0174a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0174b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0174c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0174d] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0174e] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0174f] =  I8a0037ad2845a3fbba9da380a8b8a576['h02e9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01750] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ea0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01751] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ea2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01752] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ea4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01753] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ea6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01754] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ea8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01755] =  I8a0037ad2845a3fbba9da380a8b8a576['h02eaa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01756] =  I8a0037ad2845a3fbba9da380a8b8a576['h02eac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01757] =  I8a0037ad2845a3fbba9da380a8b8a576['h02eae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01758] =  I8a0037ad2845a3fbba9da380a8b8a576['h02eb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01759] =  I8a0037ad2845a3fbba9da380a8b8a576['h02eb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0175a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02eb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0175b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02eb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0175c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02eb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0175d] =  I8a0037ad2845a3fbba9da380a8b8a576['h02eba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0175e] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ebc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0175f] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ebe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01760] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ec0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01761] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ec2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01762] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ec4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01763] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ec6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01764] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ec8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01765] =  I8a0037ad2845a3fbba9da380a8b8a576['h02eca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01766] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ecc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01767] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ece] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01768] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ed0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01769] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ed2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0176a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ed4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0176b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ed6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0176c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ed8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0176d] =  I8a0037ad2845a3fbba9da380a8b8a576['h02eda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0176e] =  I8a0037ad2845a3fbba9da380a8b8a576['h02edc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0176f] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ede] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01770] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ee0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01771] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ee2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01772] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ee4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01773] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ee6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01774] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ee8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01775] =  I8a0037ad2845a3fbba9da380a8b8a576['h02eea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01776] =  I8a0037ad2845a3fbba9da380a8b8a576['h02eec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01777] =  I8a0037ad2845a3fbba9da380a8b8a576['h02eee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01778] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ef0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01779] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ef2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0177a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ef4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0177b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ef6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0177c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ef8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0177d] =  I8a0037ad2845a3fbba9da380a8b8a576['h02efa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0177e] =  I8a0037ad2845a3fbba9da380a8b8a576['h02efc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0177f] =  I8a0037ad2845a3fbba9da380a8b8a576['h02efe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01780] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01781] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01782] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01783] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01784] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01785] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01786] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01787] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01788] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01789] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0178a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0178b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0178c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0178d] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0178e] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0178f] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01790] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01791] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01792] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01793] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01794] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01795] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01796] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01797] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01798] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01799] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0179a] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0179b] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0179c] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0179d] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0179e] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0179f] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017af] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017be] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h02f9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fa0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fa2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fa4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fa6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fa8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h02faa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017da] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017db] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017de] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017df] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fcc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fdc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fe0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fe2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fe4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fe6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fe8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h02fee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ff0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ff2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ff4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ff6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ff8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ffa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ffc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h017ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h02ffe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01800] =  I8a0037ad2845a3fbba9da380a8b8a576['h03000] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01801] =  I8a0037ad2845a3fbba9da380a8b8a576['h03002] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01802] =  I8a0037ad2845a3fbba9da380a8b8a576['h03004] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01803] =  I8a0037ad2845a3fbba9da380a8b8a576['h03006] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01804] =  I8a0037ad2845a3fbba9da380a8b8a576['h03008] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01805] =  I8a0037ad2845a3fbba9da380a8b8a576['h0300a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01806] =  I8a0037ad2845a3fbba9da380a8b8a576['h0300c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01807] =  I8a0037ad2845a3fbba9da380a8b8a576['h0300e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01808] =  I8a0037ad2845a3fbba9da380a8b8a576['h03010] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01809] =  I8a0037ad2845a3fbba9da380a8b8a576['h03012] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0180a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03014] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0180b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03016] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0180c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03018] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0180d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0301a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0180e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0301c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0180f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0301e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01810] =  I8a0037ad2845a3fbba9da380a8b8a576['h03020] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01811] =  I8a0037ad2845a3fbba9da380a8b8a576['h03022] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01812] =  I8a0037ad2845a3fbba9da380a8b8a576['h03024] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01813] =  I8a0037ad2845a3fbba9da380a8b8a576['h03026] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01814] =  I8a0037ad2845a3fbba9da380a8b8a576['h03028] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01815] =  I8a0037ad2845a3fbba9da380a8b8a576['h0302a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01816] =  I8a0037ad2845a3fbba9da380a8b8a576['h0302c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01817] =  I8a0037ad2845a3fbba9da380a8b8a576['h0302e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01818] =  I8a0037ad2845a3fbba9da380a8b8a576['h03030] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01819] =  I8a0037ad2845a3fbba9da380a8b8a576['h03032] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0181a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03034] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0181b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03036] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0181c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03038] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0181d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0303a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0181e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0303c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0181f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0303e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01820] =  I8a0037ad2845a3fbba9da380a8b8a576['h03040] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01821] =  I8a0037ad2845a3fbba9da380a8b8a576['h03042] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01822] =  I8a0037ad2845a3fbba9da380a8b8a576['h03044] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01823] =  I8a0037ad2845a3fbba9da380a8b8a576['h03046] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01824] =  I8a0037ad2845a3fbba9da380a8b8a576['h03048] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01825] =  I8a0037ad2845a3fbba9da380a8b8a576['h0304a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01826] =  I8a0037ad2845a3fbba9da380a8b8a576['h0304c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01827] =  I8a0037ad2845a3fbba9da380a8b8a576['h0304e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01828] =  I8a0037ad2845a3fbba9da380a8b8a576['h03050] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01829] =  I8a0037ad2845a3fbba9da380a8b8a576['h03052] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0182a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03054] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0182b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03056] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0182c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03058] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0182d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0305a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0182e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0305c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0182f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0305e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01830] =  I8a0037ad2845a3fbba9da380a8b8a576['h03060] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01831] =  I8a0037ad2845a3fbba9da380a8b8a576['h03062] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01832] =  I8a0037ad2845a3fbba9da380a8b8a576['h03064] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01833] =  I8a0037ad2845a3fbba9da380a8b8a576['h03066] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01834] =  I8a0037ad2845a3fbba9da380a8b8a576['h03068] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01835] =  I8a0037ad2845a3fbba9da380a8b8a576['h0306a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01836] =  I8a0037ad2845a3fbba9da380a8b8a576['h0306c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01837] =  I8a0037ad2845a3fbba9da380a8b8a576['h0306e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01838] =  I8a0037ad2845a3fbba9da380a8b8a576['h03070] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01839] =  I8a0037ad2845a3fbba9da380a8b8a576['h03072] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0183a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03074] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0183b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03076] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0183c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03078] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0183d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0307a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0183e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0307c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0183f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0307e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01840] =  I8a0037ad2845a3fbba9da380a8b8a576['h03080] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01841] =  I8a0037ad2845a3fbba9da380a8b8a576['h03082] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01842] =  I8a0037ad2845a3fbba9da380a8b8a576['h03084] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01843] =  I8a0037ad2845a3fbba9da380a8b8a576['h03086] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01844] =  I8a0037ad2845a3fbba9da380a8b8a576['h03088] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01845] =  I8a0037ad2845a3fbba9da380a8b8a576['h0308a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01846] =  I8a0037ad2845a3fbba9da380a8b8a576['h0308c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01847] =  I8a0037ad2845a3fbba9da380a8b8a576['h0308e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01848] =  I8a0037ad2845a3fbba9da380a8b8a576['h03090] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01849] =  I8a0037ad2845a3fbba9da380a8b8a576['h03092] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0184a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03094] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0184b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03096] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0184c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03098] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0184d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0309a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0184e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0309c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0184f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0309e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01850] =  I8a0037ad2845a3fbba9da380a8b8a576['h030a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01851] =  I8a0037ad2845a3fbba9da380a8b8a576['h030a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01852] =  I8a0037ad2845a3fbba9da380a8b8a576['h030a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01853] =  I8a0037ad2845a3fbba9da380a8b8a576['h030a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01854] =  I8a0037ad2845a3fbba9da380a8b8a576['h030a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01855] =  I8a0037ad2845a3fbba9da380a8b8a576['h030aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01856] =  I8a0037ad2845a3fbba9da380a8b8a576['h030ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01857] =  I8a0037ad2845a3fbba9da380a8b8a576['h030ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01858] =  I8a0037ad2845a3fbba9da380a8b8a576['h030b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01859] =  I8a0037ad2845a3fbba9da380a8b8a576['h030b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0185a] =  I8a0037ad2845a3fbba9da380a8b8a576['h030b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0185b] =  I8a0037ad2845a3fbba9da380a8b8a576['h030b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0185c] =  I8a0037ad2845a3fbba9da380a8b8a576['h030b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0185d] =  I8a0037ad2845a3fbba9da380a8b8a576['h030ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0185e] =  I8a0037ad2845a3fbba9da380a8b8a576['h030bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0185f] =  I8a0037ad2845a3fbba9da380a8b8a576['h030be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01860] =  I8a0037ad2845a3fbba9da380a8b8a576['h030c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01861] =  I8a0037ad2845a3fbba9da380a8b8a576['h030c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01862] =  I8a0037ad2845a3fbba9da380a8b8a576['h030c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01863] =  I8a0037ad2845a3fbba9da380a8b8a576['h030c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01864] =  I8a0037ad2845a3fbba9da380a8b8a576['h030c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01865] =  I8a0037ad2845a3fbba9da380a8b8a576['h030ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01866] =  I8a0037ad2845a3fbba9da380a8b8a576['h030cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01867] =  I8a0037ad2845a3fbba9da380a8b8a576['h030ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01868] =  I8a0037ad2845a3fbba9da380a8b8a576['h030d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01869] =  I8a0037ad2845a3fbba9da380a8b8a576['h030d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0186a] =  I8a0037ad2845a3fbba9da380a8b8a576['h030d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0186b] =  I8a0037ad2845a3fbba9da380a8b8a576['h030d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0186c] =  I8a0037ad2845a3fbba9da380a8b8a576['h030d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0186d] =  I8a0037ad2845a3fbba9da380a8b8a576['h030da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0186e] =  I8a0037ad2845a3fbba9da380a8b8a576['h030dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0186f] =  I8a0037ad2845a3fbba9da380a8b8a576['h030de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01870] =  I8a0037ad2845a3fbba9da380a8b8a576['h030e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01871] =  I8a0037ad2845a3fbba9da380a8b8a576['h030e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01872] =  I8a0037ad2845a3fbba9da380a8b8a576['h030e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01873] =  I8a0037ad2845a3fbba9da380a8b8a576['h030e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01874] =  I8a0037ad2845a3fbba9da380a8b8a576['h030e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01875] =  I8a0037ad2845a3fbba9da380a8b8a576['h030ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01876] =  I8a0037ad2845a3fbba9da380a8b8a576['h030ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01877] =  I8a0037ad2845a3fbba9da380a8b8a576['h030ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01878] =  I8a0037ad2845a3fbba9da380a8b8a576['h030f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01879] =  I8a0037ad2845a3fbba9da380a8b8a576['h030f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0187a] =  I8a0037ad2845a3fbba9da380a8b8a576['h030f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0187b] =  I8a0037ad2845a3fbba9da380a8b8a576['h030f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0187c] =  I8a0037ad2845a3fbba9da380a8b8a576['h030f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0187d] =  I8a0037ad2845a3fbba9da380a8b8a576['h030fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0187e] =  I8a0037ad2845a3fbba9da380a8b8a576['h030fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0187f] =  I8a0037ad2845a3fbba9da380a8b8a576['h030fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01880] =  I8a0037ad2845a3fbba9da380a8b8a576['h03100] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01881] =  I8a0037ad2845a3fbba9da380a8b8a576['h03102] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01882] =  I8a0037ad2845a3fbba9da380a8b8a576['h03104] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01883] =  I8a0037ad2845a3fbba9da380a8b8a576['h03106] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01884] =  I8a0037ad2845a3fbba9da380a8b8a576['h03108] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01885] =  I8a0037ad2845a3fbba9da380a8b8a576['h0310a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01886] =  I8a0037ad2845a3fbba9da380a8b8a576['h0310c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01887] =  I8a0037ad2845a3fbba9da380a8b8a576['h0310e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01888] =  I8a0037ad2845a3fbba9da380a8b8a576['h03110] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01889] =  I8a0037ad2845a3fbba9da380a8b8a576['h03112] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0188a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03114] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0188b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03116] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0188c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03118] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0188d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0311a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0188e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0311c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0188f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0311e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01890] =  I8a0037ad2845a3fbba9da380a8b8a576['h03120] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01891] =  I8a0037ad2845a3fbba9da380a8b8a576['h03122] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01892] =  I8a0037ad2845a3fbba9da380a8b8a576['h03124] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01893] =  I8a0037ad2845a3fbba9da380a8b8a576['h03126] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01894] =  I8a0037ad2845a3fbba9da380a8b8a576['h03128] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01895] =  I8a0037ad2845a3fbba9da380a8b8a576['h0312a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01896] =  I8a0037ad2845a3fbba9da380a8b8a576['h0312c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01897] =  I8a0037ad2845a3fbba9da380a8b8a576['h0312e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01898] =  I8a0037ad2845a3fbba9da380a8b8a576['h03130] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01899] =  I8a0037ad2845a3fbba9da380a8b8a576['h03132] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0189a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03134] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0189b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03136] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0189c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03138] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0189d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0313a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0189e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0313c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0189f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0313e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03140] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03142] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03144] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03146] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03148] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0314a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0314c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0314e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03150] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03152] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h03154] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h03156] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h03158] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0315a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0315c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018af] =  I8a0037ad2845a3fbba9da380a8b8a576['h0315e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03160] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03162] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03164] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03166] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03168] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0316a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0316c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0316e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03170] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03172] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h03174] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h03176] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h03178] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0317a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018be] =  I8a0037ad2845a3fbba9da380a8b8a576['h0317c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0317e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03180] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03182] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03184] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03186] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03188] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0318a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0318c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0318e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03190] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03192] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h03194] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h03196] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h03198] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0319a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0319c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0319e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h031a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h031a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h031a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h031a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h031a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h031aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h031ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h031ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h031b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h031b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018da] =  I8a0037ad2845a3fbba9da380a8b8a576['h031b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018db] =  I8a0037ad2845a3fbba9da380a8b8a576['h031b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h031b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h031ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018de] =  I8a0037ad2845a3fbba9da380a8b8a576['h031bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018df] =  I8a0037ad2845a3fbba9da380a8b8a576['h031be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h031c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h031c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h031c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h031c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h031c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h031ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h031cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h031ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h031d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h031d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h031d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h031d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h031d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h031da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h031dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h031de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h031e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h031e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h031e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h031e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h031e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h031ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h031ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h031ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h031f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h031f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h031f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h031f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h031f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h031fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h031fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h018ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h031fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01900] =  I8a0037ad2845a3fbba9da380a8b8a576['h03200] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01901] =  I8a0037ad2845a3fbba9da380a8b8a576['h03202] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01902] =  I8a0037ad2845a3fbba9da380a8b8a576['h03204] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01903] =  I8a0037ad2845a3fbba9da380a8b8a576['h03206] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01904] =  I8a0037ad2845a3fbba9da380a8b8a576['h03208] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01905] =  I8a0037ad2845a3fbba9da380a8b8a576['h0320a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01906] =  I8a0037ad2845a3fbba9da380a8b8a576['h0320c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01907] =  I8a0037ad2845a3fbba9da380a8b8a576['h0320e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01908] =  I8a0037ad2845a3fbba9da380a8b8a576['h03210] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01909] =  I8a0037ad2845a3fbba9da380a8b8a576['h03212] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0190a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03214] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0190b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03216] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0190c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03218] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0190d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0321a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0190e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0321c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0190f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0321e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01910] =  I8a0037ad2845a3fbba9da380a8b8a576['h03220] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01911] =  I8a0037ad2845a3fbba9da380a8b8a576['h03222] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01912] =  I8a0037ad2845a3fbba9da380a8b8a576['h03224] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01913] =  I8a0037ad2845a3fbba9da380a8b8a576['h03226] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01914] =  I8a0037ad2845a3fbba9da380a8b8a576['h03228] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01915] =  I8a0037ad2845a3fbba9da380a8b8a576['h0322a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01916] =  I8a0037ad2845a3fbba9da380a8b8a576['h0322c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01917] =  I8a0037ad2845a3fbba9da380a8b8a576['h0322e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01918] =  I8a0037ad2845a3fbba9da380a8b8a576['h03230] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01919] =  I8a0037ad2845a3fbba9da380a8b8a576['h03232] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0191a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03234] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0191b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03236] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0191c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03238] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0191d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0323a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0191e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0323c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0191f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0323e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01920] =  I8a0037ad2845a3fbba9da380a8b8a576['h03240] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01921] =  I8a0037ad2845a3fbba9da380a8b8a576['h03242] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01922] =  I8a0037ad2845a3fbba9da380a8b8a576['h03244] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01923] =  I8a0037ad2845a3fbba9da380a8b8a576['h03246] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01924] =  I8a0037ad2845a3fbba9da380a8b8a576['h03248] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01925] =  I8a0037ad2845a3fbba9da380a8b8a576['h0324a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01926] =  I8a0037ad2845a3fbba9da380a8b8a576['h0324c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01927] =  I8a0037ad2845a3fbba9da380a8b8a576['h0324e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01928] =  I8a0037ad2845a3fbba9da380a8b8a576['h03250] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01929] =  I8a0037ad2845a3fbba9da380a8b8a576['h03252] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0192a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03254] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0192b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03256] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0192c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03258] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0192d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0325a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0192e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0325c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0192f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0325e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01930] =  I8a0037ad2845a3fbba9da380a8b8a576['h03260] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01931] =  I8a0037ad2845a3fbba9da380a8b8a576['h03262] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01932] =  I8a0037ad2845a3fbba9da380a8b8a576['h03264] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01933] =  I8a0037ad2845a3fbba9da380a8b8a576['h03266] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01934] =  I8a0037ad2845a3fbba9da380a8b8a576['h03268] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01935] =  I8a0037ad2845a3fbba9da380a8b8a576['h0326a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01936] =  I8a0037ad2845a3fbba9da380a8b8a576['h0326c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01937] =  I8a0037ad2845a3fbba9da380a8b8a576['h0326e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01938] =  I8a0037ad2845a3fbba9da380a8b8a576['h03270] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01939] =  I8a0037ad2845a3fbba9da380a8b8a576['h03272] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0193a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03274] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0193b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03276] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0193c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03278] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0193d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0327a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0193e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0327c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0193f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0327e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01940] =  I8a0037ad2845a3fbba9da380a8b8a576['h03280] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01941] =  I8a0037ad2845a3fbba9da380a8b8a576['h03282] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01942] =  I8a0037ad2845a3fbba9da380a8b8a576['h03284] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01943] =  I8a0037ad2845a3fbba9da380a8b8a576['h03286] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01944] =  I8a0037ad2845a3fbba9da380a8b8a576['h03288] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01945] =  I8a0037ad2845a3fbba9da380a8b8a576['h0328a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01946] =  I8a0037ad2845a3fbba9da380a8b8a576['h0328c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01947] =  I8a0037ad2845a3fbba9da380a8b8a576['h0328e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01948] =  I8a0037ad2845a3fbba9da380a8b8a576['h03290] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01949] =  I8a0037ad2845a3fbba9da380a8b8a576['h03292] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0194a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03294] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0194b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03296] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0194c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03298] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0194d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0329a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0194e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0329c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0194f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0329e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01950] =  I8a0037ad2845a3fbba9da380a8b8a576['h032a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01951] =  I8a0037ad2845a3fbba9da380a8b8a576['h032a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01952] =  I8a0037ad2845a3fbba9da380a8b8a576['h032a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01953] =  I8a0037ad2845a3fbba9da380a8b8a576['h032a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01954] =  I8a0037ad2845a3fbba9da380a8b8a576['h032a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01955] =  I8a0037ad2845a3fbba9da380a8b8a576['h032aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01956] =  I8a0037ad2845a3fbba9da380a8b8a576['h032ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01957] =  I8a0037ad2845a3fbba9da380a8b8a576['h032ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01958] =  I8a0037ad2845a3fbba9da380a8b8a576['h032b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01959] =  I8a0037ad2845a3fbba9da380a8b8a576['h032b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0195a] =  I8a0037ad2845a3fbba9da380a8b8a576['h032b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0195b] =  I8a0037ad2845a3fbba9da380a8b8a576['h032b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0195c] =  I8a0037ad2845a3fbba9da380a8b8a576['h032b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0195d] =  I8a0037ad2845a3fbba9da380a8b8a576['h032ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0195e] =  I8a0037ad2845a3fbba9da380a8b8a576['h032bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0195f] =  I8a0037ad2845a3fbba9da380a8b8a576['h032be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01960] =  I8a0037ad2845a3fbba9da380a8b8a576['h032c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01961] =  I8a0037ad2845a3fbba9da380a8b8a576['h032c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01962] =  I8a0037ad2845a3fbba9da380a8b8a576['h032c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01963] =  I8a0037ad2845a3fbba9da380a8b8a576['h032c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01964] =  I8a0037ad2845a3fbba9da380a8b8a576['h032c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01965] =  I8a0037ad2845a3fbba9da380a8b8a576['h032ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01966] =  I8a0037ad2845a3fbba9da380a8b8a576['h032cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01967] =  I8a0037ad2845a3fbba9da380a8b8a576['h032ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01968] =  I8a0037ad2845a3fbba9da380a8b8a576['h032d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01969] =  I8a0037ad2845a3fbba9da380a8b8a576['h032d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0196a] =  I8a0037ad2845a3fbba9da380a8b8a576['h032d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0196b] =  I8a0037ad2845a3fbba9da380a8b8a576['h032d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0196c] =  I8a0037ad2845a3fbba9da380a8b8a576['h032d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0196d] =  I8a0037ad2845a3fbba9da380a8b8a576['h032da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0196e] =  I8a0037ad2845a3fbba9da380a8b8a576['h032dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0196f] =  I8a0037ad2845a3fbba9da380a8b8a576['h032de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01970] =  I8a0037ad2845a3fbba9da380a8b8a576['h032e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01971] =  I8a0037ad2845a3fbba9da380a8b8a576['h032e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01972] =  I8a0037ad2845a3fbba9da380a8b8a576['h032e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01973] =  I8a0037ad2845a3fbba9da380a8b8a576['h032e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01974] =  I8a0037ad2845a3fbba9da380a8b8a576['h032e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01975] =  I8a0037ad2845a3fbba9da380a8b8a576['h032ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01976] =  I8a0037ad2845a3fbba9da380a8b8a576['h032ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01977] =  I8a0037ad2845a3fbba9da380a8b8a576['h032ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01978] =  I8a0037ad2845a3fbba9da380a8b8a576['h032f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01979] =  I8a0037ad2845a3fbba9da380a8b8a576['h032f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0197a] =  I8a0037ad2845a3fbba9da380a8b8a576['h032f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0197b] =  I8a0037ad2845a3fbba9da380a8b8a576['h032f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0197c] =  I8a0037ad2845a3fbba9da380a8b8a576['h032f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0197d] =  I8a0037ad2845a3fbba9da380a8b8a576['h032fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0197e] =  I8a0037ad2845a3fbba9da380a8b8a576['h032fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0197f] =  I8a0037ad2845a3fbba9da380a8b8a576['h032fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01980] =  I8a0037ad2845a3fbba9da380a8b8a576['h03300] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01981] =  I8a0037ad2845a3fbba9da380a8b8a576['h03302] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01982] =  I8a0037ad2845a3fbba9da380a8b8a576['h03304] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01983] =  I8a0037ad2845a3fbba9da380a8b8a576['h03306] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01984] =  I8a0037ad2845a3fbba9da380a8b8a576['h03308] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01985] =  I8a0037ad2845a3fbba9da380a8b8a576['h0330a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01986] =  I8a0037ad2845a3fbba9da380a8b8a576['h0330c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01987] =  I8a0037ad2845a3fbba9da380a8b8a576['h0330e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01988] =  I8a0037ad2845a3fbba9da380a8b8a576['h03310] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01989] =  I8a0037ad2845a3fbba9da380a8b8a576['h03312] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0198a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03314] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0198b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03316] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0198c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03318] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0198d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0331a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0198e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0331c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0198f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0331e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01990] =  I8a0037ad2845a3fbba9da380a8b8a576['h03320] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01991] =  I8a0037ad2845a3fbba9da380a8b8a576['h03322] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01992] =  I8a0037ad2845a3fbba9da380a8b8a576['h03324] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01993] =  I8a0037ad2845a3fbba9da380a8b8a576['h03326] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01994] =  I8a0037ad2845a3fbba9da380a8b8a576['h03328] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01995] =  I8a0037ad2845a3fbba9da380a8b8a576['h0332a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01996] =  I8a0037ad2845a3fbba9da380a8b8a576['h0332c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01997] =  I8a0037ad2845a3fbba9da380a8b8a576['h0332e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01998] =  I8a0037ad2845a3fbba9da380a8b8a576['h03330] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01999] =  I8a0037ad2845a3fbba9da380a8b8a576['h03332] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0199a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03334] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0199b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03336] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0199c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03338] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0199d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0333a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0199e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0333c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0199f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0333e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03340] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03342] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03344] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03346] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03348] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0334a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0334c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0334e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03350] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03352] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h03354] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h03356] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h03358] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0335a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0335c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019af] =  I8a0037ad2845a3fbba9da380a8b8a576['h0335e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03360] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03362] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03364] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03366] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03368] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0336a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0336c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0336e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03370] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03372] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h03374] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h03376] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h03378] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0337a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019be] =  I8a0037ad2845a3fbba9da380a8b8a576['h0337c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0337e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03380] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03382] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03384] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03386] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03388] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0338a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0338c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0338e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03390] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03392] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h03394] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h03396] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h03398] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0339a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0339c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0339e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h033a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h033a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h033a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h033a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h033a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h033aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h033ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h033ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h033b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h033b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019da] =  I8a0037ad2845a3fbba9da380a8b8a576['h033b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019db] =  I8a0037ad2845a3fbba9da380a8b8a576['h033b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h033b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h033ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019de] =  I8a0037ad2845a3fbba9da380a8b8a576['h033bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019df] =  I8a0037ad2845a3fbba9da380a8b8a576['h033be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h033c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h033c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h033c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h033c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h033c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h033ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h033cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h033ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h033d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h033d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h033d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h033d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h033d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h033da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h033dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h033de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h033e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h033e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h033e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h033e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h033e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h033ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h033ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h033ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h033f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h033f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h033f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h033f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h033f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h033fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h033fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h019ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h033fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a00] =  I8a0037ad2845a3fbba9da380a8b8a576['h03400] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a01] =  I8a0037ad2845a3fbba9da380a8b8a576['h03402] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a02] =  I8a0037ad2845a3fbba9da380a8b8a576['h03404] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a03] =  I8a0037ad2845a3fbba9da380a8b8a576['h03406] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a04] =  I8a0037ad2845a3fbba9da380a8b8a576['h03408] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a05] =  I8a0037ad2845a3fbba9da380a8b8a576['h0340a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a06] =  I8a0037ad2845a3fbba9da380a8b8a576['h0340c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a07] =  I8a0037ad2845a3fbba9da380a8b8a576['h0340e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a08] =  I8a0037ad2845a3fbba9da380a8b8a576['h03410] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a09] =  I8a0037ad2845a3fbba9da380a8b8a576['h03412] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a0a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03414] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a0b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03416] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a0c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03418] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a0d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0341a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a0e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0341c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a0f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0341e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a10] =  I8a0037ad2845a3fbba9da380a8b8a576['h03420] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a11] =  I8a0037ad2845a3fbba9da380a8b8a576['h03422] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a12] =  I8a0037ad2845a3fbba9da380a8b8a576['h03424] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a13] =  I8a0037ad2845a3fbba9da380a8b8a576['h03426] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a14] =  I8a0037ad2845a3fbba9da380a8b8a576['h03428] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a15] =  I8a0037ad2845a3fbba9da380a8b8a576['h0342a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a16] =  I8a0037ad2845a3fbba9da380a8b8a576['h0342c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a17] =  I8a0037ad2845a3fbba9da380a8b8a576['h0342e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a18] =  I8a0037ad2845a3fbba9da380a8b8a576['h03430] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a19] =  I8a0037ad2845a3fbba9da380a8b8a576['h03432] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a1a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03434] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a1b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03436] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a1c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03438] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a1d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0343a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a1e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0343c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a1f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0343e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a20] =  I8a0037ad2845a3fbba9da380a8b8a576['h03440] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a21] =  I8a0037ad2845a3fbba9da380a8b8a576['h03442] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a22] =  I8a0037ad2845a3fbba9da380a8b8a576['h03444] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a23] =  I8a0037ad2845a3fbba9da380a8b8a576['h03446] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a24] =  I8a0037ad2845a3fbba9da380a8b8a576['h03448] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a25] =  I8a0037ad2845a3fbba9da380a8b8a576['h0344a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a26] =  I8a0037ad2845a3fbba9da380a8b8a576['h0344c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a27] =  I8a0037ad2845a3fbba9da380a8b8a576['h0344e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a28] =  I8a0037ad2845a3fbba9da380a8b8a576['h03450] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a29] =  I8a0037ad2845a3fbba9da380a8b8a576['h03452] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a2a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03454] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a2b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03456] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a2c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03458] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a2d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0345a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a2e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0345c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a2f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0345e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a30] =  I8a0037ad2845a3fbba9da380a8b8a576['h03460] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a31] =  I8a0037ad2845a3fbba9da380a8b8a576['h03462] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a32] =  I8a0037ad2845a3fbba9da380a8b8a576['h03464] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a33] =  I8a0037ad2845a3fbba9da380a8b8a576['h03466] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a34] =  I8a0037ad2845a3fbba9da380a8b8a576['h03468] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a35] =  I8a0037ad2845a3fbba9da380a8b8a576['h0346a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a36] =  I8a0037ad2845a3fbba9da380a8b8a576['h0346c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a37] =  I8a0037ad2845a3fbba9da380a8b8a576['h0346e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a38] =  I8a0037ad2845a3fbba9da380a8b8a576['h03470] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a39] =  I8a0037ad2845a3fbba9da380a8b8a576['h03472] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a3a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03474] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a3b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03476] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a3c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03478] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a3d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0347a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a3e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0347c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a3f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0347e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a40] =  I8a0037ad2845a3fbba9da380a8b8a576['h03480] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a41] =  I8a0037ad2845a3fbba9da380a8b8a576['h03482] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a42] =  I8a0037ad2845a3fbba9da380a8b8a576['h03484] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a43] =  I8a0037ad2845a3fbba9da380a8b8a576['h03486] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a44] =  I8a0037ad2845a3fbba9da380a8b8a576['h03488] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a45] =  I8a0037ad2845a3fbba9da380a8b8a576['h0348a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a46] =  I8a0037ad2845a3fbba9da380a8b8a576['h0348c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a47] =  I8a0037ad2845a3fbba9da380a8b8a576['h0348e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a48] =  I8a0037ad2845a3fbba9da380a8b8a576['h03490] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a49] =  I8a0037ad2845a3fbba9da380a8b8a576['h03492] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a4a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03494] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a4b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03496] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a4c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03498] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a4d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0349a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a4e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0349c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a4f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0349e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a50] =  I8a0037ad2845a3fbba9da380a8b8a576['h034a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a51] =  I8a0037ad2845a3fbba9da380a8b8a576['h034a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a52] =  I8a0037ad2845a3fbba9da380a8b8a576['h034a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a53] =  I8a0037ad2845a3fbba9da380a8b8a576['h034a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a54] =  I8a0037ad2845a3fbba9da380a8b8a576['h034a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a55] =  I8a0037ad2845a3fbba9da380a8b8a576['h034aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a56] =  I8a0037ad2845a3fbba9da380a8b8a576['h034ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a57] =  I8a0037ad2845a3fbba9da380a8b8a576['h034ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a58] =  I8a0037ad2845a3fbba9da380a8b8a576['h034b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a59] =  I8a0037ad2845a3fbba9da380a8b8a576['h034b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a5a] =  I8a0037ad2845a3fbba9da380a8b8a576['h034b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a5b] =  I8a0037ad2845a3fbba9da380a8b8a576['h034b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a5c] =  I8a0037ad2845a3fbba9da380a8b8a576['h034b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a5d] =  I8a0037ad2845a3fbba9da380a8b8a576['h034ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a5e] =  I8a0037ad2845a3fbba9da380a8b8a576['h034bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a5f] =  I8a0037ad2845a3fbba9da380a8b8a576['h034be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a60] =  I8a0037ad2845a3fbba9da380a8b8a576['h034c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a61] =  I8a0037ad2845a3fbba9da380a8b8a576['h034c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a62] =  I8a0037ad2845a3fbba9da380a8b8a576['h034c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a63] =  I8a0037ad2845a3fbba9da380a8b8a576['h034c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a64] =  I8a0037ad2845a3fbba9da380a8b8a576['h034c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a65] =  I8a0037ad2845a3fbba9da380a8b8a576['h034ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a66] =  I8a0037ad2845a3fbba9da380a8b8a576['h034cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a67] =  I8a0037ad2845a3fbba9da380a8b8a576['h034ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a68] =  I8a0037ad2845a3fbba9da380a8b8a576['h034d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a69] =  I8a0037ad2845a3fbba9da380a8b8a576['h034d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a6a] =  I8a0037ad2845a3fbba9da380a8b8a576['h034d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a6b] =  I8a0037ad2845a3fbba9da380a8b8a576['h034d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a6c] =  I8a0037ad2845a3fbba9da380a8b8a576['h034d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a6d] =  I8a0037ad2845a3fbba9da380a8b8a576['h034da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a6e] =  I8a0037ad2845a3fbba9da380a8b8a576['h034dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a6f] =  I8a0037ad2845a3fbba9da380a8b8a576['h034de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a70] =  I8a0037ad2845a3fbba9da380a8b8a576['h034e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a71] =  I8a0037ad2845a3fbba9da380a8b8a576['h034e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a72] =  I8a0037ad2845a3fbba9da380a8b8a576['h034e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a73] =  I8a0037ad2845a3fbba9da380a8b8a576['h034e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a74] =  I8a0037ad2845a3fbba9da380a8b8a576['h034e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a75] =  I8a0037ad2845a3fbba9da380a8b8a576['h034ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a76] =  I8a0037ad2845a3fbba9da380a8b8a576['h034ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a77] =  I8a0037ad2845a3fbba9da380a8b8a576['h034ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a78] =  I8a0037ad2845a3fbba9da380a8b8a576['h034f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a79] =  I8a0037ad2845a3fbba9da380a8b8a576['h034f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a7a] =  I8a0037ad2845a3fbba9da380a8b8a576['h034f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a7b] =  I8a0037ad2845a3fbba9da380a8b8a576['h034f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a7c] =  I8a0037ad2845a3fbba9da380a8b8a576['h034f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a7d] =  I8a0037ad2845a3fbba9da380a8b8a576['h034fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a7e] =  I8a0037ad2845a3fbba9da380a8b8a576['h034fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a7f] =  I8a0037ad2845a3fbba9da380a8b8a576['h034fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a80] =  I8a0037ad2845a3fbba9da380a8b8a576['h03500] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a81] =  I8a0037ad2845a3fbba9da380a8b8a576['h03502] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a82] =  I8a0037ad2845a3fbba9da380a8b8a576['h03504] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a83] =  I8a0037ad2845a3fbba9da380a8b8a576['h03506] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a84] =  I8a0037ad2845a3fbba9da380a8b8a576['h03508] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a85] =  I8a0037ad2845a3fbba9da380a8b8a576['h0350a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a86] =  I8a0037ad2845a3fbba9da380a8b8a576['h0350c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a87] =  I8a0037ad2845a3fbba9da380a8b8a576['h0350e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a88] =  I8a0037ad2845a3fbba9da380a8b8a576['h03510] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a89] =  I8a0037ad2845a3fbba9da380a8b8a576['h03512] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a8a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03514] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a8b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03516] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a8c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03518] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a8d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0351a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a8e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0351c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a8f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0351e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a90] =  I8a0037ad2845a3fbba9da380a8b8a576['h03520] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a91] =  I8a0037ad2845a3fbba9da380a8b8a576['h03522] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a92] =  I8a0037ad2845a3fbba9da380a8b8a576['h03524] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a93] =  I8a0037ad2845a3fbba9da380a8b8a576['h03526] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a94] =  I8a0037ad2845a3fbba9da380a8b8a576['h03528] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a95] =  I8a0037ad2845a3fbba9da380a8b8a576['h0352a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a96] =  I8a0037ad2845a3fbba9da380a8b8a576['h0352c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a97] =  I8a0037ad2845a3fbba9da380a8b8a576['h0352e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a98] =  I8a0037ad2845a3fbba9da380a8b8a576['h03530] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a99] =  I8a0037ad2845a3fbba9da380a8b8a576['h03532] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a9a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03534] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a9b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03536] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a9c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03538] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a9d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0353a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a9e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0353c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01a9f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0353e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01aa0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03540] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01aa1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03542] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01aa2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03544] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01aa3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03546] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01aa4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03548] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01aa5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0354a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01aa6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0354c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01aa7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0354e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01aa8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03550] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01aa9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03552] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01aaa] =  I8a0037ad2845a3fbba9da380a8b8a576['h03554] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01aab] =  I8a0037ad2845a3fbba9da380a8b8a576['h03556] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01aac] =  I8a0037ad2845a3fbba9da380a8b8a576['h03558] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01aad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0355a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01aae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0355c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01aaf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0355e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ab0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03560] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ab1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03562] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ab2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03564] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ab3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03566] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ab4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03568] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ab5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0356a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ab6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0356c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ab7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0356e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ab8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03570] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ab9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03572] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01aba] =  I8a0037ad2845a3fbba9da380a8b8a576['h03574] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01abb] =  I8a0037ad2845a3fbba9da380a8b8a576['h03576] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01abc] =  I8a0037ad2845a3fbba9da380a8b8a576['h03578] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01abd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0357a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01abe] =  I8a0037ad2845a3fbba9da380a8b8a576['h0357c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01abf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0357e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ac0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03580] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ac1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03582] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ac2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03584] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ac3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03586] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ac4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03588] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ac5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0358a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ac6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0358c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ac7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0358e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ac8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03590] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ac9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03592] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01aca] =  I8a0037ad2845a3fbba9da380a8b8a576['h03594] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01acb] =  I8a0037ad2845a3fbba9da380a8b8a576['h03596] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01acc] =  I8a0037ad2845a3fbba9da380a8b8a576['h03598] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01acd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0359a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ace] =  I8a0037ad2845a3fbba9da380a8b8a576['h0359c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01acf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0359e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ad0] =  I8a0037ad2845a3fbba9da380a8b8a576['h035a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ad1] =  I8a0037ad2845a3fbba9da380a8b8a576['h035a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ad2] =  I8a0037ad2845a3fbba9da380a8b8a576['h035a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ad3] =  I8a0037ad2845a3fbba9da380a8b8a576['h035a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ad4] =  I8a0037ad2845a3fbba9da380a8b8a576['h035a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ad5] =  I8a0037ad2845a3fbba9da380a8b8a576['h035aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ad6] =  I8a0037ad2845a3fbba9da380a8b8a576['h035ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ad7] =  I8a0037ad2845a3fbba9da380a8b8a576['h035ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ad8] =  I8a0037ad2845a3fbba9da380a8b8a576['h035b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ad9] =  I8a0037ad2845a3fbba9da380a8b8a576['h035b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ada] =  I8a0037ad2845a3fbba9da380a8b8a576['h035b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01adb] =  I8a0037ad2845a3fbba9da380a8b8a576['h035b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01adc] =  I8a0037ad2845a3fbba9da380a8b8a576['h035b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01add] =  I8a0037ad2845a3fbba9da380a8b8a576['h035ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ade] =  I8a0037ad2845a3fbba9da380a8b8a576['h035bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01adf] =  I8a0037ad2845a3fbba9da380a8b8a576['h035be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ae0] =  I8a0037ad2845a3fbba9da380a8b8a576['h035c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ae1] =  I8a0037ad2845a3fbba9da380a8b8a576['h035c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ae2] =  I8a0037ad2845a3fbba9da380a8b8a576['h035c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ae3] =  I8a0037ad2845a3fbba9da380a8b8a576['h035c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ae4] =  I8a0037ad2845a3fbba9da380a8b8a576['h035c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ae5] =  I8a0037ad2845a3fbba9da380a8b8a576['h035ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ae6] =  I8a0037ad2845a3fbba9da380a8b8a576['h035cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ae7] =  I8a0037ad2845a3fbba9da380a8b8a576['h035ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ae8] =  I8a0037ad2845a3fbba9da380a8b8a576['h035d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ae9] =  I8a0037ad2845a3fbba9da380a8b8a576['h035d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01aea] =  I8a0037ad2845a3fbba9da380a8b8a576['h035d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01aeb] =  I8a0037ad2845a3fbba9da380a8b8a576['h035d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01aec] =  I8a0037ad2845a3fbba9da380a8b8a576['h035d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01aed] =  I8a0037ad2845a3fbba9da380a8b8a576['h035da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01aee] =  I8a0037ad2845a3fbba9da380a8b8a576['h035dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01aef] =  I8a0037ad2845a3fbba9da380a8b8a576['h035de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01af0] =  I8a0037ad2845a3fbba9da380a8b8a576['h035e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01af1] =  I8a0037ad2845a3fbba9da380a8b8a576['h035e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01af2] =  I8a0037ad2845a3fbba9da380a8b8a576['h035e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01af3] =  I8a0037ad2845a3fbba9da380a8b8a576['h035e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01af4] =  I8a0037ad2845a3fbba9da380a8b8a576['h035e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01af5] =  I8a0037ad2845a3fbba9da380a8b8a576['h035ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01af6] =  I8a0037ad2845a3fbba9da380a8b8a576['h035ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01af7] =  I8a0037ad2845a3fbba9da380a8b8a576['h035ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01af8] =  I8a0037ad2845a3fbba9da380a8b8a576['h035f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01af9] =  I8a0037ad2845a3fbba9da380a8b8a576['h035f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01afa] =  I8a0037ad2845a3fbba9da380a8b8a576['h035f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01afb] =  I8a0037ad2845a3fbba9da380a8b8a576['h035f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01afc] =  I8a0037ad2845a3fbba9da380a8b8a576['h035f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01afd] =  I8a0037ad2845a3fbba9da380a8b8a576['h035fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01afe] =  I8a0037ad2845a3fbba9da380a8b8a576['h035fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01aff] =  I8a0037ad2845a3fbba9da380a8b8a576['h035fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b00] =  I8a0037ad2845a3fbba9da380a8b8a576['h03600] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b01] =  I8a0037ad2845a3fbba9da380a8b8a576['h03602] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b02] =  I8a0037ad2845a3fbba9da380a8b8a576['h03604] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b03] =  I8a0037ad2845a3fbba9da380a8b8a576['h03606] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b04] =  I8a0037ad2845a3fbba9da380a8b8a576['h03608] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b05] =  I8a0037ad2845a3fbba9da380a8b8a576['h0360a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b06] =  I8a0037ad2845a3fbba9da380a8b8a576['h0360c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b07] =  I8a0037ad2845a3fbba9da380a8b8a576['h0360e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b08] =  I8a0037ad2845a3fbba9da380a8b8a576['h03610] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b09] =  I8a0037ad2845a3fbba9da380a8b8a576['h03612] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b0a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03614] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b0b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03616] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b0c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03618] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b0d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0361a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b0e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0361c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b0f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0361e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b10] =  I8a0037ad2845a3fbba9da380a8b8a576['h03620] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b11] =  I8a0037ad2845a3fbba9da380a8b8a576['h03622] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b12] =  I8a0037ad2845a3fbba9da380a8b8a576['h03624] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b13] =  I8a0037ad2845a3fbba9da380a8b8a576['h03626] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b14] =  I8a0037ad2845a3fbba9da380a8b8a576['h03628] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b15] =  I8a0037ad2845a3fbba9da380a8b8a576['h0362a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b16] =  I8a0037ad2845a3fbba9da380a8b8a576['h0362c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b17] =  I8a0037ad2845a3fbba9da380a8b8a576['h0362e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b18] =  I8a0037ad2845a3fbba9da380a8b8a576['h03630] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b19] =  I8a0037ad2845a3fbba9da380a8b8a576['h03632] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b1a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03634] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b1b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03636] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b1c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03638] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b1d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0363a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b1e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0363c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b1f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0363e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b20] =  I8a0037ad2845a3fbba9da380a8b8a576['h03640] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b21] =  I8a0037ad2845a3fbba9da380a8b8a576['h03642] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b22] =  I8a0037ad2845a3fbba9da380a8b8a576['h03644] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b23] =  I8a0037ad2845a3fbba9da380a8b8a576['h03646] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b24] =  I8a0037ad2845a3fbba9da380a8b8a576['h03648] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b25] =  I8a0037ad2845a3fbba9da380a8b8a576['h0364a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b26] =  I8a0037ad2845a3fbba9da380a8b8a576['h0364c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b27] =  I8a0037ad2845a3fbba9da380a8b8a576['h0364e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b28] =  I8a0037ad2845a3fbba9da380a8b8a576['h03650] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b29] =  I8a0037ad2845a3fbba9da380a8b8a576['h03652] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b2a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03654] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b2b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03656] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b2c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03658] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b2d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0365a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b2e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0365c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b2f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0365e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b30] =  I8a0037ad2845a3fbba9da380a8b8a576['h03660] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b31] =  I8a0037ad2845a3fbba9da380a8b8a576['h03662] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b32] =  I8a0037ad2845a3fbba9da380a8b8a576['h03664] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b33] =  I8a0037ad2845a3fbba9da380a8b8a576['h03666] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b34] =  I8a0037ad2845a3fbba9da380a8b8a576['h03668] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b35] =  I8a0037ad2845a3fbba9da380a8b8a576['h0366a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b36] =  I8a0037ad2845a3fbba9da380a8b8a576['h0366c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b37] =  I8a0037ad2845a3fbba9da380a8b8a576['h0366e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b38] =  I8a0037ad2845a3fbba9da380a8b8a576['h03670] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b39] =  I8a0037ad2845a3fbba9da380a8b8a576['h03672] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b3a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03674] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b3b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03676] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b3c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03678] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b3d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0367a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b3e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0367c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b3f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0367e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b40] =  I8a0037ad2845a3fbba9da380a8b8a576['h03680] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b41] =  I8a0037ad2845a3fbba9da380a8b8a576['h03682] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b42] =  I8a0037ad2845a3fbba9da380a8b8a576['h03684] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b43] =  I8a0037ad2845a3fbba9da380a8b8a576['h03686] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b44] =  I8a0037ad2845a3fbba9da380a8b8a576['h03688] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b45] =  I8a0037ad2845a3fbba9da380a8b8a576['h0368a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b46] =  I8a0037ad2845a3fbba9da380a8b8a576['h0368c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b47] =  I8a0037ad2845a3fbba9da380a8b8a576['h0368e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b48] =  I8a0037ad2845a3fbba9da380a8b8a576['h03690] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b49] =  I8a0037ad2845a3fbba9da380a8b8a576['h03692] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b4a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03694] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b4b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03696] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b4c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03698] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b4d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0369a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b4e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0369c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b4f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0369e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b50] =  I8a0037ad2845a3fbba9da380a8b8a576['h036a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b51] =  I8a0037ad2845a3fbba9da380a8b8a576['h036a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b52] =  I8a0037ad2845a3fbba9da380a8b8a576['h036a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b53] =  I8a0037ad2845a3fbba9da380a8b8a576['h036a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b54] =  I8a0037ad2845a3fbba9da380a8b8a576['h036a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b55] =  I8a0037ad2845a3fbba9da380a8b8a576['h036aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b56] =  I8a0037ad2845a3fbba9da380a8b8a576['h036ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b57] =  I8a0037ad2845a3fbba9da380a8b8a576['h036ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b58] =  I8a0037ad2845a3fbba9da380a8b8a576['h036b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b59] =  I8a0037ad2845a3fbba9da380a8b8a576['h036b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b5a] =  I8a0037ad2845a3fbba9da380a8b8a576['h036b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b5b] =  I8a0037ad2845a3fbba9da380a8b8a576['h036b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b5c] =  I8a0037ad2845a3fbba9da380a8b8a576['h036b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b5d] =  I8a0037ad2845a3fbba9da380a8b8a576['h036ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b5e] =  I8a0037ad2845a3fbba9da380a8b8a576['h036bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b5f] =  I8a0037ad2845a3fbba9da380a8b8a576['h036be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b60] =  I8a0037ad2845a3fbba9da380a8b8a576['h036c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b61] =  I8a0037ad2845a3fbba9da380a8b8a576['h036c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b62] =  I8a0037ad2845a3fbba9da380a8b8a576['h036c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b63] =  I8a0037ad2845a3fbba9da380a8b8a576['h036c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b64] =  I8a0037ad2845a3fbba9da380a8b8a576['h036c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b65] =  I8a0037ad2845a3fbba9da380a8b8a576['h036ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b66] =  I8a0037ad2845a3fbba9da380a8b8a576['h036cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b67] =  I8a0037ad2845a3fbba9da380a8b8a576['h036ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b68] =  I8a0037ad2845a3fbba9da380a8b8a576['h036d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b69] =  I8a0037ad2845a3fbba9da380a8b8a576['h036d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b6a] =  I8a0037ad2845a3fbba9da380a8b8a576['h036d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b6b] =  I8a0037ad2845a3fbba9da380a8b8a576['h036d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b6c] =  I8a0037ad2845a3fbba9da380a8b8a576['h036d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b6d] =  I8a0037ad2845a3fbba9da380a8b8a576['h036da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b6e] =  I8a0037ad2845a3fbba9da380a8b8a576['h036dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b6f] =  I8a0037ad2845a3fbba9da380a8b8a576['h036de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b70] =  I8a0037ad2845a3fbba9da380a8b8a576['h036e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b71] =  I8a0037ad2845a3fbba9da380a8b8a576['h036e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b72] =  I8a0037ad2845a3fbba9da380a8b8a576['h036e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b73] =  I8a0037ad2845a3fbba9da380a8b8a576['h036e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b74] =  I8a0037ad2845a3fbba9da380a8b8a576['h036e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b75] =  I8a0037ad2845a3fbba9da380a8b8a576['h036ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b76] =  I8a0037ad2845a3fbba9da380a8b8a576['h036ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b77] =  I8a0037ad2845a3fbba9da380a8b8a576['h036ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b78] =  I8a0037ad2845a3fbba9da380a8b8a576['h036f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b79] =  I8a0037ad2845a3fbba9da380a8b8a576['h036f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b7a] =  I8a0037ad2845a3fbba9da380a8b8a576['h036f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b7b] =  I8a0037ad2845a3fbba9da380a8b8a576['h036f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b7c] =  I8a0037ad2845a3fbba9da380a8b8a576['h036f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b7d] =  I8a0037ad2845a3fbba9da380a8b8a576['h036fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b7e] =  I8a0037ad2845a3fbba9da380a8b8a576['h036fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b7f] =  I8a0037ad2845a3fbba9da380a8b8a576['h036fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b80] =  I8a0037ad2845a3fbba9da380a8b8a576['h03700] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b81] =  I8a0037ad2845a3fbba9da380a8b8a576['h03702] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b82] =  I8a0037ad2845a3fbba9da380a8b8a576['h03704] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b83] =  I8a0037ad2845a3fbba9da380a8b8a576['h03706] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b84] =  I8a0037ad2845a3fbba9da380a8b8a576['h03708] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b85] =  I8a0037ad2845a3fbba9da380a8b8a576['h0370a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b86] =  I8a0037ad2845a3fbba9da380a8b8a576['h0370c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b87] =  I8a0037ad2845a3fbba9da380a8b8a576['h0370e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b88] =  I8a0037ad2845a3fbba9da380a8b8a576['h03710] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b89] =  I8a0037ad2845a3fbba9da380a8b8a576['h03712] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b8a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03714] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b8b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03716] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b8c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03718] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b8d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0371a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b8e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0371c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b8f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0371e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b90] =  I8a0037ad2845a3fbba9da380a8b8a576['h03720] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b91] =  I8a0037ad2845a3fbba9da380a8b8a576['h03722] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b92] =  I8a0037ad2845a3fbba9da380a8b8a576['h03724] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b93] =  I8a0037ad2845a3fbba9da380a8b8a576['h03726] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b94] =  I8a0037ad2845a3fbba9da380a8b8a576['h03728] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b95] =  I8a0037ad2845a3fbba9da380a8b8a576['h0372a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b96] =  I8a0037ad2845a3fbba9da380a8b8a576['h0372c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b97] =  I8a0037ad2845a3fbba9da380a8b8a576['h0372e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b98] =  I8a0037ad2845a3fbba9da380a8b8a576['h03730] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b99] =  I8a0037ad2845a3fbba9da380a8b8a576['h03732] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b9a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03734] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b9b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03736] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b9c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03738] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b9d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0373a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b9e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0373c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01b9f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0373e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ba0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03740] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ba1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03742] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ba2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03744] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ba3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03746] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ba4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03748] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ba5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0374a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ba6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0374c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ba7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0374e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ba8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03750] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ba9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03752] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01baa] =  I8a0037ad2845a3fbba9da380a8b8a576['h03754] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bab] =  I8a0037ad2845a3fbba9da380a8b8a576['h03756] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bac] =  I8a0037ad2845a3fbba9da380a8b8a576['h03758] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0375a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0375c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01baf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0375e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bb0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03760] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bb1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03762] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bb2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03764] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bb3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03766] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bb4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03768] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bb5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0376a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bb6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0376c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bb7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0376e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bb8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03770] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bb9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03772] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bba] =  I8a0037ad2845a3fbba9da380a8b8a576['h03774] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bbb] =  I8a0037ad2845a3fbba9da380a8b8a576['h03776] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bbc] =  I8a0037ad2845a3fbba9da380a8b8a576['h03778] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bbd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0377a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bbe] =  I8a0037ad2845a3fbba9da380a8b8a576['h0377c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bbf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0377e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bc0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03780] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bc1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03782] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bc2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03784] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bc3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03786] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bc4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03788] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bc5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0378a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bc6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0378c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bc7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0378e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bc8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03790] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bc9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03792] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bca] =  I8a0037ad2845a3fbba9da380a8b8a576['h03794] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bcb] =  I8a0037ad2845a3fbba9da380a8b8a576['h03796] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bcc] =  I8a0037ad2845a3fbba9da380a8b8a576['h03798] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bcd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0379a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0379c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bcf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0379e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bd0] =  I8a0037ad2845a3fbba9da380a8b8a576['h037a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bd1] =  I8a0037ad2845a3fbba9da380a8b8a576['h037a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bd2] =  I8a0037ad2845a3fbba9da380a8b8a576['h037a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bd3] =  I8a0037ad2845a3fbba9da380a8b8a576['h037a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bd4] =  I8a0037ad2845a3fbba9da380a8b8a576['h037a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bd5] =  I8a0037ad2845a3fbba9da380a8b8a576['h037aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bd6] =  I8a0037ad2845a3fbba9da380a8b8a576['h037ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bd7] =  I8a0037ad2845a3fbba9da380a8b8a576['h037ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bd8] =  I8a0037ad2845a3fbba9da380a8b8a576['h037b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bd9] =  I8a0037ad2845a3fbba9da380a8b8a576['h037b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bda] =  I8a0037ad2845a3fbba9da380a8b8a576['h037b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bdb] =  I8a0037ad2845a3fbba9da380a8b8a576['h037b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bdc] =  I8a0037ad2845a3fbba9da380a8b8a576['h037b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bdd] =  I8a0037ad2845a3fbba9da380a8b8a576['h037ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bde] =  I8a0037ad2845a3fbba9da380a8b8a576['h037bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bdf] =  I8a0037ad2845a3fbba9da380a8b8a576['h037be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01be0] =  I8a0037ad2845a3fbba9da380a8b8a576['h037c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01be1] =  I8a0037ad2845a3fbba9da380a8b8a576['h037c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01be2] =  I8a0037ad2845a3fbba9da380a8b8a576['h037c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01be3] =  I8a0037ad2845a3fbba9da380a8b8a576['h037c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01be4] =  I8a0037ad2845a3fbba9da380a8b8a576['h037c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01be5] =  I8a0037ad2845a3fbba9da380a8b8a576['h037ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01be6] =  I8a0037ad2845a3fbba9da380a8b8a576['h037cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01be7] =  I8a0037ad2845a3fbba9da380a8b8a576['h037ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01be8] =  I8a0037ad2845a3fbba9da380a8b8a576['h037d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01be9] =  I8a0037ad2845a3fbba9da380a8b8a576['h037d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bea] =  I8a0037ad2845a3fbba9da380a8b8a576['h037d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01beb] =  I8a0037ad2845a3fbba9da380a8b8a576['h037d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bec] =  I8a0037ad2845a3fbba9da380a8b8a576['h037d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bed] =  I8a0037ad2845a3fbba9da380a8b8a576['h037da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bee] =  I8a0037ad2845a3fbba9da380a8b8a576['h037dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bef] =  I8a0037ad2845a3fbba9da380a8b8a576['h037de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bf0] =  I8a0037ad2845a3fbba9da380a8b8a576['h037e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bf1] =  I8a0037ad2845a3fbba9da380a8b8a576['h037e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bf2] =  I8a0037ad2845a3fbba9da380a8b8a576['h037e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bf3] =  I8a0037ad2845a3fbba9da380a8b8a576['h037e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bf4] =  I8a0037ad2845a3fbba9da380a8b8a576['h037e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bf5] =  I8a0037ad2845a3fbba9da380a8b8a576['h037ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bf6] =  I8a0037ad2845a3fbba9da380a8b8a576['h037ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bf7] =  I8a0037ad2845a3fbba9da380a8b8a576['h037ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bf8] =  I8a0037ad2845a3fbba9da380a8b8a576['h037f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bf9] =  I8a0037ad2845a3fbba9da380a8b8a576['h037f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bfa] =  I8a0037ad2845a3fbba9da380a8b8a576['h037f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bfb] =  I8a0037ad2845a3fbba9da380a8b8a576['h037f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bfc] =  I8a0037ad2845a3fbba9da380a8b8a576['h037f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bfd] =  I8a0037ad2845a3fbba9da380a8b8a576['h037fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bfe] =  I8a0037ad2845a3fbba9da380a8b8a576['h037fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01bff] =  I8a0037ad2845a3fbba9da380a8b8a576['h037fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c00] =  I8a0037ad2845a3fbba9da380a8b8a576['h03800] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c01] =  I8a0037ad2845a3fbba9da380a8b8a576['h03802] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c02] =  I8a0037ad2845a3fbba9da380a8b8a576['h03804] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c03] =  I8a0037ad2845a3fbba9da380a8b8a576['h03806] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c04] =  I8a0037ad2845a3fbba9da380a8b8a576['h03808] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c05] =  I8a0037ad2845a3fbba9da380a8b8a576['h0380a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c06] =  I8a0037ad2845a3fbba9da380a8b8a576['h0380c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c07] =  I8a0037ad2845a3fbba9da380a8b8a576['h0380e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c08] =  I8a0037ad2845a3fbba9da380a8b8a576['h03810] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c09] =  I8a0037ad2845a3fbba9da380a8b8a576['h03812] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c0a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03814] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c0b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03816] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c0c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03818] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c0d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0381a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c0e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0381c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c0f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0381e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c10] =  I8a0037ad2845a3fbba9da380a8b8a576['h03820] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c11] =  I8a0037ad2845a3fbba9da380a8b8a576['h03822] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c12] =  I8a0037ad2845a3fbba9da380a8b8a576['h03824] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c13] =  I8a0037ad2845a3fbba9da380a8b8a576['h03826] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c14] =  I8a0037ad2845a3fbba9da380a8b8a576['h03828] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c15] =  I8a0037ad2845a3fbba9da380a8b8a576['h0382a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c16] =  I8a0037ad2845a3fbba9da380a8b8a576['h0382c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c17] =  I8a0037ad2845a3fbba9da380a8b8a576['h0382e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c18] =  I8a0037ad2845a3fbba9da380a8b8a576['h03830] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c19] =  I8a0037ad2845a3fbba9da380a8b8a576['h03832] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c1a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03834] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c1b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03836] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c1c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03838] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c1d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0383a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c1e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0383c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c1f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0383e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c20] =  I8a0037ad2845a3fbba9da380a8b8a576['h03840] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c21] =  I8a0037ad2845a3fbba9da380a8b8a576['h03842] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c22] =  I8a0037ad2845a3fbba9da380a8b8a576['h03844] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c23] =  I8a0037ad2845a3fbba9da380a8b8a576['h03846] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c24] =  I8a0037ad2845a3fbba9da380a8b8a576['h03848] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c25] =  I8a0037ad2845a3fbba9da380a8b8a576['h0384a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c26] =  I8a0037ad2845a3fbba9da380a8b8a576['h0384c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c27] =  I8a0037ad2845a3fbba9da380a8b8a576['h0384e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c28] =  I8a0037ad2845a3fbba9da380a8b8a576['h03850] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c29] =  I8a0037ad2845a3fbba9da380a8b8a576['h03852] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c2a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03854] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c2b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03856] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c2c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03858] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c2d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0385a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c2e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0385c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c2f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0385e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c30] =  I8a0037ad2845a3fbba9da380a8b8a576['h03860] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c31] =  I8a0037ad2845a3fbba9da380a8b8a576['h03862] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c32] =  I8a0037ad2845a3fbba9da380a8b8a576['h03864] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c33] =  I8a0037ad2845a3fbba9da380a8b8a576['h03866] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c34] =  I8a0037ad2845a3fbba9da380a8b8a576['h03868] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c35] =  I8a0037ad2845a3fbba9da380a8b8a576['h0386a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c36] =  I8a0037ad2845a3fbba9da380a8b8a576['h0386c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c37] =  I8a0037ad2845a3fbba9da380a8b8a576['h0386e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c38] =  I8a0037ad2845a3fbba9da380a8b8a576['h03870] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c39] =  I8a0037ad2845a3fbba9da380a8b8a576['h03872] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c3a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03874] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c3b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03876] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c3c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03878] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c3d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0387a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c3e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0387c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c3f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0387e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c40] =  I8a0037ad2845a3fbba9da380a8b8a576['h03880] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c41] =  I8a0037ad2845a3fbba9da380a8b8a576['h03882] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c42] =  I8a0037ad2845a3fbba9da380a8b8a576['h03884] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c43] =  I8a0037ad2845a3fbba9da380a8b8a576['h03886] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c44] =  I8a0037ad2845a3fbba9da380a8b8a576['h03888] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c45] =  I8a0037ad2845a3fbba9da380a8b8a576['h0388a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c46] =  I8a0037ad2845a3fbba9da380a8b8a576['h0388c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c47] =  I8a0037ad2845a3fbba9da380a8b8a576['h0388e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c48] =  I8a0037ad2845a3fbba9da380a8b8a576['h03890] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c49] =  I8a0037ad2845a3fbba9da380a8b8a576['h03892] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c4a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03894] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c4b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03896] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c4c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03898] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c4d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0389a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c4e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0389c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c4f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0389e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c50] =  I8a0037ad2845a3fbba9da380a8b8a576['h038a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c51] =  I8a0037ad2845a3fbba9da380a8b8a576['h038a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c52] =  I8a0037ad2845a3fbba9da380a8b8a576['h038a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c53] =  I8a0037ad2845a3fbba9da380a8b8a576['h038a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c54] =  I8a0037ad2845a3fbba9da380a8b8a576['h038a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c55] =  I8a0037ad2845a3fbba9da380a8b8a576['h038aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c56] =  I8a0037ad2845a3fbba9da380a8b8a576['h038ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c57] =  I8a0037ad2845a3fbba9da380a8b8a576['h038ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c58] =  I8a0037ad2845a3fbba9da380a8b8a576['h038b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c59] =  I8a0037ad2845a3fbba9da380a8b8a576['h038b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c5a] =  I8a0037ad2845a3fbba9da380a8b8a576['h038b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c5b] =  I8a0037ad2845a3fbba9da380a8b8a576['h038b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c5c] =  I8a0037ad2845a3fbba9da380a8b8a576['h038b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c5d] =  I8a0037ad2845a3fbba9da380a8b8a576['h038ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c5e] =  I8a0037ad2845a3fbba9da380a8b8a576['h038bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c5f] =  I8a0037ad2845a3fbba9da380a8b8a576['h038be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c60] =  I8a0037ad2845a3fbba9da380a8b8a576['h038c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c61] =  I8a0037ad2845a3fbba9da380a8b8a576['h038c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c62] =  I8a0037ad2845a3fbba9da380a8b8a576['h038c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c63] =  I8a0037ad2845a3fbba9da380a8b8a576['h038c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c64] =  I8a0037ad2845a3fbba9da380a8b8a576['h038c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c65] =  I8a0037ad2845a3fbba9da380a8b8a576['h038ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c66] =  I8a0037ad2845a3fbba9da380a8b8a576['h038cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c67] =  I8a0037ad2845a3fbba9da380a8b8a576['h038ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c68] =  I8a0037ad2845a3fbba9da380a8b8a576['h038d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c69] =  I8a0037ad2845a3fbba9da380a8b8a576['h038d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c6a] =  I8a0037ad2845a3fbba9da380a8b8a576['h038d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c6b] =  I8a0037ad2845a3fbba9da380a8b8a576['h038d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c6c] =  I8a0037ad2845a3fbba9da380a8b8a576['h038d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c6d] =  I8a0037ad2845a3fbba9da380a8b8a576['h038da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c6e] =  I8a0037ad2845a3fbba9da380a8b8a576['h038dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c6f] =  I8a0037ad2845a3fbba9da380a8b8a576['h038de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c70] =  I8a0037ad2845a3fbba9da380a8b8a576['h038e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c71] =  I8a0037ad2845a3fbba9da380a8b8a576['h038e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c72] =  I8a0037ad2845a3fbba9da380a8b8a576['h038e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c73] =  I8a0037ad2845a3fbba9da380a8b8a576['h038e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c74] =  I8a0037ad2845a3fbba9da380a8b8a576['h038e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c75] =  I8a0037ad2845a3fbba9da380a8b8a576['h038ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c76] =  I8a0037ad2845a3fbba9da380a8b8a576['h038ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c77] =  I8a0037ad2845a3fbba9da380a8b8a576['h038ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c78] =  I8a0037ad2845a3fbba9da380a8b8a576['h038f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c79] =  I8a0037ad2845a3fbba9da380a8b8a576['h038f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c7a] =  I8a0037ad2845a3fbba9da380a8b8a576['h038f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c7b] =  I8a0037ad2845a3fbba9da380a8b8a576['h038f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c7c] =  I8a0037ad2845a3fbba9da380a8b8a576['h038f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c7d] =  I8a0037ad2845a3fbba9da380a8b8a576['h038fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c7e] =  I8a0037ad2845a3fbba9da380a8b8a576['h038fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c7f] =  I8a0037ad2845a3fbba9da380a8b8a576['h038fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c80] =  I8a0037ad2845a3fbba9da380a8b8a576['h03900] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c81] =  I8a0037ad2845a3fbba9da380a8b8a576['h03902] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c82] =  I8a0037ad2845a3fbba9da380a8b8a576['h03904] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c83] =  I8a0037ad2845a3fbba9da380a8b8a576['h03906] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c84] =  I8a0037ad2845a3fbba9da380a8b8a576['h03908] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c85] =  I8a0037ad2845a3fbba9da380a8b8a576['h0390a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c86] =  I8a0037ad2845a3fbba9da380a8b8a576['h0390c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c87] =  I8a0037ad2845a3fbba9da380a8b8a576['h0390e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c88] =  I8a0037ad2845a3fbba9da380a8b8a576['h03910] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c89] =  I8a0037ad2845a3fbba9da380a8b8a576['h03912] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c8a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03914] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c8b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03916] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c8c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03918] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c8d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0391a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c8e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0391c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c8f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0391e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c90] =  I8a0037ad2845a3fbba9da380a8b8a576['h03920] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c91] =  I8a0037ad2845a3fbba9da380a8b8a576['h03922] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c92] =  I8a0037ad2845a3fbba9da380a8b8a576['h03924] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c93] =  I8a0037ad2845a3fbba9da380a8b8a576['h03926] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c94] =  I8a0037ad2845a3fbba9da380a8b8a576['h03928] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c95] =  I8a0037ad2845a3fbba9da380a8b8a576['h0392a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c96] =  I8a0037ad2845a3fbba9da380a8b8a576['h0392c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c97] =  I8a0037ad2845a3fbba9da380a8b8a576['h0392e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c98] =  I8a0037ad2845a3fbba9da380a8b8a576['h03930] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c99] =  I8a0037ad2845a3fbba9da380a8b8a576['h03932] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c9a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03934] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c9b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03936] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c9c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03938] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c9d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0393a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c9e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0393c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01c9f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0393e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ca0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03940] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ca1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03942] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ca2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03944] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ca3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03946] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ca4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03948] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ca5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0394a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ca6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0394c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ca7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0394e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ca8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03950] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ca9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03952] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01caa] =  I8a0037ad2845a3fbba9da380a8b8a576['h03954] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cab] =  I8a0037ad2845a3fbba9da380a8b8a576['h03956] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cac] =  I8a0037ad2845a3fbba9da380a8b8a576['h03958] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0395a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0395c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01caf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0395e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cb0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03960] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cb1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03962] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cb2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03964] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cb3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03966] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cb4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03968] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cb5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0396a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cb6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0396c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cb7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0396e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cb8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03970] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cb9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03972] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cba] =  I8a0037ad2845a3fbba9da380a8b8a576['h03974] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cbb] =  I8a0037ad2845a3fbba9da380a8b8a576['h03976] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cbc] =  I8a0037ad2845a3fbba9da380a8b8a576['h03978] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cbd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0397a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cbe] =  I8a0037ad2845a3fbba9da380a8b8a576['h0397c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cbf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0397e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cc0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03980] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cc1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03982] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cc2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03984] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cc3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03986] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cc4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03988] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cc5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0398a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cc6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0398c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cc7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0398e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cc8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03990] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cc9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03992] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cca] =  I8a0037ad2845a3fbba9da380a8b8a576['h03994] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ccb] =  I8a0037ad2845a3fbba9da380a8b8a576['h03996] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ccc] =  I8a0037ad2845a3fbba9da380a8b8a576['h03998] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ccd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0399a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0399c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ccf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0399e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cd0] =  I8a0037ad2845a3fbba9da380a8b8a576['h039a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cd1] =  I8a0037ad2845a3fbba9da380a8b8a576['h039a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cd2] =  I8a0037ad2845a3fbba9da380a8b8a576['h039a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cd3] =  I8a0037ad2845a3fbba9da380a8b8a576['h039a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cd4] =  I8a0037ad2845a3fbba9da380a8b8a576['h039a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cd5] =  I8a0037ad2845a3fbba9da380a8b8a576['h039aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cd6] =  I8a0037ad2845a3fbba9da380a8b8a576['h039ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cd7] =  I8a0037ad2845a3fbba9da380a8b8a576['h039ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cd8] =  I8a0037ad2845a3fbba9da380a8b8a576['h039b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cd9] =  I8a0037ad2845a3fbba9da380a8b8a576['h039b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cda] =  I8a0037ad2845a3fbba9da380a8b8a576['h039b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cdb] =  I8a0037ad2845a3fbba9da380a8b8a576['h039b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cdc] =  I8a0037ad2845a3fbba9da380a8b8a576['h039b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cdd] =  I8a0037ad2845a3fbba9da380a8b8a576['h039ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cde] =  I8a0037ad2845a3fbba9da380a8b8a576['h039bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cdf] =  I8a0037ad2845a3fbba9da380a8b8a576['h039be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ce0] =  I8a0037ad2845a3fbba9da380a8b8a576['h039c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ce1] =  I8a0037ad2845a3fbba9da380a8b8a576['h039c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ce2] =  I8a0037ad2845a3fbba9da380a8b8a576['h039c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ce3] =  I8a0037ad2845a3fbba9da380a8b8a576['h039c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ce4] =  I8a0037ad2845a3fbba9da380a8b8a576['h039c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ce5] =  I8a0037ad2845a3fbba9da380a8b8a576['h039ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ce6] =  I8a0037ad2845a3fbba9da380a8b8a576['h039cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ce7] =  I8a0037ad2845a3fbba9da380a8b8a576['h039ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ce8] =  I8a0037ad2845a3fbba9da380a8b8a576['h039d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ce9] =  I8a0037ad2845a3fbba9da380a8b8a576['h039d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cea] =  I8a0037ad2845a3fbba9da380a8b8a576['h039d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ceb] =  I8a0037ad2845a3fbba9da380a8b8a576['h039d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cec] =  I8a0037ad2845a3fbba9da380a8b8a576['h039d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ced] =  I8a0037ad2845a3fbba9da380a8b8a576['h039da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cee] =  I8a0037ad2845a3fbba9da380a8b8a576['h039dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cef] =  I8a0037ad2845a3fbba9da380a8b8a576['h039de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cf0] =  I8a0037ad2845a3fbba9da380a8b8a576['h039e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cf1] =  I8a0037ad2845a3fbba9da380a8b8a576['h039e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cf2] =  I8a0037ad2845a3fbba9da380a8b8a576['h039e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cf3] =  I8a0037ad2845a3fbba9da380a8b8a576['h039e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cf4] =  I8a0037ad2845a3fbba9da380a8b8a576['h039e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cf5] =  I8a0037ad2845a3fbba9da380a8b8a576['h039ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cf6] =  I8a0037ad2845a3fbba9da380a8b8a576['h039ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cf7] =  I8a0037ad2845a3fbba9da380a8b8a576['h039ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cf8] =  I8a0037ad2845a3fbba9da380a8b8a576['h039f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cf9] =  I8a0037ad2845a3fbba9da380a8b8a576['h039f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cfa] =  I8a0037ad2845a3fbba9da380a8b8a576['h039f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cfb] =  I8a0037ad2845a3fbba9da380a8b8a576['h039f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cfc] =  I8a0037ad2845a3fbba9da380a8b8a576['h039f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cfd] =  I8a0037ad2845a3fbba9da380a8b8a576['h039fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cfe] =  I8a0037ad2845a3fbba9da380a8b8a576['h039fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01cff] =  I8a0037ad2845a3fbba9da380a8b8a576['h039fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d00] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d01] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d02] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d03] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d04] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d05] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d06] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d07] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d08] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d09] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d0a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d0b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d0c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d0d] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d0e] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d0f] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d10] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d11] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d12] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d13] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d14] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d15] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d16] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d17] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d18] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d19] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d1a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d1b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d1c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d1d] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d1e] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d1f] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d20] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d21] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d22] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d23] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d24] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d25] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d26] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d27] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d28] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d29] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d2a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d2b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d2c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d2d] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d2e] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d2f] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d30] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d31] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d32] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d33] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d34] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d35] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d36] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d37] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d38] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d39] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d3a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d3b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d3c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d3d] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d3e] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d3f] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d40] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d41] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d42] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d43] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d44] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d45] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d46] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d47] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d48] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d49] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d4a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d4b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d4c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d4d] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d4e] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d4f] =  I8a0037ad2845a3fbba9da380a8b8a576['h03a9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d50] =  I8a0037ad2845a3fbba9da380a8b8a576['h03aa0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d51] =  I8a0037ad2845a3fbba9da380a8b8a576['h03aa2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d52] =  I8a0037ad2845a3fbba9da380a8b8a576['h03aa4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d53] =  I8a0037ad2845a3fbba9da380a8b8a576['h03aa6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d54] =  I8a0037ad2845a3fbba9da380a8b8a576['h03aa8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d55] =  I8a0037ad2845a3fbba9da380a8b8a576['h03aaa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d56] =  I8a0037ad2845a3fbba9da380a8b8a576['h03aac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d57] =  I8a0037ad2845a3fbba9da380a8b8a576['h03aae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d58] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ab0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d59] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ab2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d5a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ab4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d5b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ab6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d5c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ab8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d5d] =  I8a0037ad2845a3fbba9da380a8b8a576['h03aba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d5e] =  I8a0037ad2845a3fbba9da380a8b8a576['h03abc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d5f] =  I8a0037ad2845a3fbba9da380a8b8a576['h03abe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d60] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ac0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d61] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ac2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d62] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ac4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d63] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ac6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d64] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ac8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d65] =  I8a0037ad2845a3fbba9da380a8b8a576['h03aca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d66] =  I8a0037ad2845a3fbba9da380a8b8a576['h03acc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d67] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ace] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d68] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ad0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d69] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ad2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d6a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ad4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d6b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ad6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d6c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ad8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d6d] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ada] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d6e] =  I8a0037ad2845a3fbba9da380a8b8a576['h03adc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d6f] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ade] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d70] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ae0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d71] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ae2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d72] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ae4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d73] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ae6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d74] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ae8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d75] =  I8a0037ad2845a3fbba9da380a8b8a576['h03aea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d76] =  I8a0037ad2845a3fbba9da380a8b8a576['h03aec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d77] =  I8a0037ad2845a3fbba9da380a8b8a576['h03aee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d78] =  I8a0037ad2845a3fbba9da380a8b8a576['h03af0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d79] =  I8a0037ad2845a3fbba9da380a8b8a576['h03af2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d7a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03af4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d7b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03af6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d7c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03af8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d7d] =  I8a0037ad2845a3fbba9da380a8b8a576['h03afa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d7e] =  I8a0037ad2845a3fbba9da380a8b8a576['h03afc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d7f] =  I8a0037ad2845a3fbba9da380a8b8a576['h03afe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d80] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d81] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d82] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d83] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d84] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d85] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d86] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d87] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d88] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d89] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d8a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d8b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d8c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d8d] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d8e] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d8f] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d90] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d91] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d92] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d93] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d94] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d95] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d96] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d97] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d98] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d99] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d9a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d9b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d9c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d9d] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d9e] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01d9f] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01da0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01da1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01da2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01da3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01da4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01da5] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01da6] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01da7] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01da8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01da9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01daa] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dab] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dac] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dad] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dae] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01daf] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01db0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01db1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01db2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01db3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01db4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01db5] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01db6] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01db7] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01db8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01db9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dba] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dbb] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dbc] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dbd] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dbe] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dbf] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dc0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dc1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dc2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dc3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dc4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dc5] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dc6] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dc7] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dc8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dc9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dca] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dcb] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dcc] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dcd] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dce] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dcf] =  I8a0037ad2845a3fbba9da380a8b8a576['h03b9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dd0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ba0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dd1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ba2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dd2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ba4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dd3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ba6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dd4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ba8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dd5] =  I8a0037ad2845a3fbba9da380a8b8a576['h03baa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dd6] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dd7] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dd8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dd9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dda] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ddb] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ddc] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ddd] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dde] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ddf] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01de0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01de1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01de2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01de3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01de4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01de5] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01de6] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bcc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01de7] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01de8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01de9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dea] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01deb] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dec] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ded] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dee] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bdc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01def] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01df0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03be0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01df1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03be2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01df2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03be4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01df3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03be6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01df4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03be8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01df5] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01df6] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01df7] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01df8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bf0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01df9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bf2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dfa] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bf4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dfb] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bf6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dfc] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bf8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dfd] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bfa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dfe] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bfc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01dff] =  I8a0037ad2845a3fbba9da380a8b8a576['h03bfe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e00] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e01] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e02] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e03] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e04] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e05] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e06] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e07] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e08] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e09] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e0a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e0b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e0c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e0d] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e0e] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e0f] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e10] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e11] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e12] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e13] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e14] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e15] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e16] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e17] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e18] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e19] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e1a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e1b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e1c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e1d] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e1e] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e1f] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e20] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e21] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e22] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e23] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e24] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e25] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e26] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e27] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e28] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e29] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e2a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e2b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e2c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e2d] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e2e] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e2f] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e30] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e31] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e32] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e33] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e34] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e35] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e36] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e37] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e38] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e39] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e3a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e3b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e3c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e3d] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e3e] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e3f] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e40] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e41] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e42] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e43] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e44] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e45] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e46] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e47] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e48] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e49] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e4a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e4b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e4c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e4d] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e4e] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e4f] =  I8a0037ad2845a3fbba9da380a8b8a576['h03c9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e50] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ca0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e51] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ca2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e52] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ca4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e53] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ca6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e54] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ca8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e55] =  I8a0037ad2845a3fbba9da380a8b8a576['h03caa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e56] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e57] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e58] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e59] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e5a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e5b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e5c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e5d] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e5e] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e5f] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e60] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e61] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e62] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e63] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e64] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e65] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e66] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ccc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e67] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e68] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e69] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e6a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e6b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e6c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e6d] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e6e] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cdc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e6f] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e70] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ce0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e71] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ce2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e72] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ce4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e73] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ce6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e74] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ce8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e75] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e76] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e77] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e78] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cf0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e79] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cf2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e7a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cf4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e7b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cf6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e7c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cf8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e7d] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cfa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e7e] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cfc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e7f] =  I8a0037ad2845a3fbba9da380a8b8a576['h03cfe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e80] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e81] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e82] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e83] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e84] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e85] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e86] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e87] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e88] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e89] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e8a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e8b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e8c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e8d] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e8e] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e8f] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e90] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e91] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e92] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e93] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e94] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e95] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e96] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e97] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e98] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e99] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e9a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e9b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e9c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e9d] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e9e] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01e9f] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ea0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ea1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ea2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ea3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ea4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ea5] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ea6] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ea7] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ea8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ea9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01eaa] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01eab] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01eac] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ead] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01eae] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01eaf] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01eb0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01eb1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01eb2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01eb3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01eb4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01eb5] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01eb6] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01eb7] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01eb8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01eb9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01eba] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ebb] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ebc] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ebd] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ebe] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ebf] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ec0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ec1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ec2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ec3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ec4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ec5] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ec6] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ec7] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ec8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ec9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01eca] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ecb] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ecc] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ecd] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ece] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ecf] =  I8a0037ad2845a3fbba9da380a8b8a576['h03d9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ed0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03da0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ed1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03da2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ed2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03da4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ed3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03da6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ed4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03da8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ed5] =  I8a0037ad2845a3fbba9da380a8b8a576['h03daa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ed6] =  I8a0037ad2845a3fbba9da380a8b8a576['h03dac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ed7] =  I8a0037ad2845a3fbba9da380a8b8a576['h03dae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ed8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03db0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ed9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03db2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01eda] =  I8a0037ad2845a3fbba9da380a8b8a576['h03db4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01edb] =  I8a0037ad2845a3fbba9da380a8b8a576['h03db6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01edc] =  I8a0037ad2845a3fbba9da380a8b8a576['h03db8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01edd] =  I8a0037ad2845a3fbba9da380a8b8a576['h03dba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ede] =  I8a0037ad2845a3fbba9da380a8b8a576['h03dbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01edf] =  I8a0037ad2845a3fbba9da380a8b8a576['h03dbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ee0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03dc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ee1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03dc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ee2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03dc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ee3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03dc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ee4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03dc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ee5] =  I8a0037ad2845a3fbba9da380a8b8a576['h03dca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ee6] =  I8a0037ad2845a3fbba9da380a8b8a576['h03dcc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ee7] =  I8a0037ad2845a3fbba9da380a8b8a576['h03dce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ee8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03dd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ee9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03dd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01eea] =  I8a0037ad2845a3fbba9da380a8b8a576['h03dd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01eeb] =  I8a0037ad2845a3fbba9da380a8b8a576['h03dd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01eec] =  I8a0037ad2845a3fbba9da380a8b8a576['h03dd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01eed] =  I8a0037ad2845a3fbba9da380a8b8a576['h03dda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01eee] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ddc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01eef] =  I8a0037ad2845a3fbba9da380a8b8a576['h03dde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ef0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03de0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ef1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03de2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ef2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03de4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ef3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03de6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ef4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03de8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ef5] =  I8a0037ad2845a3fbba9da380a8b8a576['h03dea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ef6] =  I8a0037ad2845a3fbba9da380a8b8a576['h03dec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ef7] =  I8a0037ad2845a3fbba9da380a8b8a576['h03dee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ef8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03df0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ef9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03df2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01efa] =  I8a0037ad2845a3fbba9da380a8b8a576['h03df4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01efb] =  I8a0037ad2845a3fbba9da380a8b8a576['h03df6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01efc] =  I8a0037ad2845a3fbba9da380a8b8a576['h03df8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01efd] =  I8a0037ad2845a3fbba9da380a8b8a576['h03dfa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01efe] =  I8a0037ad2845a3fbba9da380a8b8a576['h03dfc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01eff] =  I8a0037ad2845a3fbba9da380a8b8a576['h03dfe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f00] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f01] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f02] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f03] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f04] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f05] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f06] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f07] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f08] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f09] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f0a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f0b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f0c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f0d] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f0e] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f0f] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f10] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f11] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f12] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f13] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f14] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f15] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f16] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f17] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f18] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f19] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f1a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f1b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f1c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f1d] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f1e] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f1f] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f20] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f21] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f22] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f23] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f24] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f25] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f26] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f27] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f28] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f29] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f2a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f2b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f2c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f2d] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f2e] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f2f] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f30] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f31] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f32] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f33] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f34] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f35] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f36] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f37] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f38] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f39] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f3a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f3b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f3c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f3d] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f3e] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f3f] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f40] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f41] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f42] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f43] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f44] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f45] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f46] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f47] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f48] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f49] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f4a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f4b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f4c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f4d] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f4e] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f4f] =  I8a0037ad2845a3fbba9da380a8b8a576['h03e9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f50] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ea0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f51] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ea2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f52] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ea4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f53] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ea6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f54] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ea8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f55] =  I8a0037ad2845a3fbba9da380a8b8a576['h03eaa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f56] =  I8a0037ad2845a3fbba9da380a8b8a576['h03eac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f57] =  I8a0037ad2845a3fbba9da380a8b8a576['h03eae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f58] =  I8a0037ad2845a3fbba9da380a8b8a576['h03eb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f59] =  I8a0037ad2845a3fbba9da380a8b8a576['h03eb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f5a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03eb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f5b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03eb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f5c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03eb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f5d] =  I8a0037ad2845a3fbba9da380a8b8a576['h03eba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f5e] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ebc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f5f] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ebe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f60] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ec0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f61] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ec2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f62] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ec4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f63] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ec6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f64] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ec8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f65] =  I8a0037ad2845a3fbba9da380a8b8a576['h03eca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f66] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ecc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f67] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ece] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f68] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ed0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f69] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ed2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f6a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ed4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f6b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ed6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f6c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ed8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f6d] =  I8a0037ad2845a3fbba9da380a8b8a576['h03eda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f6e] =  I8a0037ad2845a3fbba9da380a8b8a576['h03edc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f6f] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ede] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f70] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ee0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f71] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ee2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f72] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ee4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f73] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ee6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f74] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ee8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f75] =  I8a0037ad2845a3fbba9da380a8b8a576['h03eea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f76] =  I8a0037ad2845a3fbba9da380a8b8a576['h03eec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f77] =  I8a0037ad2845a3fbba9da380a8b8a576['h03eee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f78] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ef0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f79] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ef2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f7a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ef4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f7b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ef6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f7c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ef8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f7d] =  I8a0037ad2845a3fbba9da380a8b8a576['h03efa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f7e] =  I8a0037ad2845a3fbba9da380a8b8a576['h03efc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f7f] =  I8a0037ad2845a3fbba9da380a8b8a576['h03efe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f80] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f81] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f82] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f83] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f84] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f85] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f86] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f87] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f88] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f89] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f8a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f8b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f8c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f8d] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f8e] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f8f] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f90] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f91] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f92] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f93] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f94] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f95] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f96] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f97] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f98] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f99] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f9a] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f9b] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f9c] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f9d] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f9e] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01f9f] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fa0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fa1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fa2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fa3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fa4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fa5] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fa6] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fa7] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fa8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fa9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01faa] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fab] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fac] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fad] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fae] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01faf] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fb0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fb1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fb2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fb3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fb4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fb5] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fb6] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fb7] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fb8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fb9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fba] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fbb] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fbc] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fbd] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fbe] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fbf] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fc0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fc1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fc2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fc3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fc4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fc5] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fc6] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fc7] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fc8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fc9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fca] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fcb] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fcc] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fcd] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fce] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fcf] =  I8a0037ad2845a3fbba9da380a8b8a576['h03f9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fd0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fa0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fd1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fa2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fd2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fa4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fd3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fa6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fd4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fa8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fd5] =  I8a0037ad2845a3fbba9da380a8b8a576['h03faa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fd6] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fd7] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fd8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fd9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fda] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fdb] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fdc] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fdd] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fde] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fdf] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fe0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fe1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fe2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fe3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fe4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fe5] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fe6] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fcc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fe7] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fe8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fe9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fea] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01feb] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fec] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fed] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fee] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fdc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fef] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ff0] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fe0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ff1] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fe2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ff2] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fe4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ff3] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fe6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ff4] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fe8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ff5] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ff6] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ff7] =  I8a0037ad2845a3fbba9da380a8b8a576['h03fee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ff8] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ff0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ff9] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ff2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ffa] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ff4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ffb] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ff6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ffc] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ff8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ffd] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ffa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01ffe] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ffc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h01fff] =  I8a0037ad2845a3fbba9da380a8b8a576['h03ffe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02000] =  I8a0037ad2845a3fbba9da380a8b8a576['h04000] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02001] =  I8a0037ad2845a3fbba9da380a8b8a576['h04002] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02002] =  I8a0037ad2845a3fbba9da380a8b8a576['h04004] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02003] =  I8a0037ad2845a3fbba9da380a8b8a576['h04006] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02004] =  I8a0037ad2845a3fbba9da380a8b8a576['h04008] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02005] =  I8a0037ad2845a3fbba9da380a8b8a576['h0400a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02006] =  I8a0037ad2845a3fbba9da380a8b8a576['h0400c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02007] =  I8a0037ad2845a3fbba9da380a8b8a576['h0400e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02008] =  I8a0037ad2845a3fbba9da380a8b8a576['h04010] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02009] =  I8a0037ad2845a3fbba9da380a8b8a576['h04012] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0200a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04014] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0200b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04016] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0200c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04018] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0200d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0401a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0200e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0401c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0200f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0401e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02010] =  I8a0037ad2845a3fbba9da380a8b8a576['h04020] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02011] =  I8a0037ad2845a3fbba9da380a8b8a576['h04022] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02012] =  I8a0037ad2845a3fbba9da380a8b8a576['h04024] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02013] =  I8a0037ad2845a3fbba9da380a8b8a576['h04026] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02014] =  I8a0037ad2845a3fbba9da380a8b8a576['h04028] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02015] =  I8a0037ad2845a3fbba9da380a8b8a576['h0402a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02016] =  I8a0037ad2845a3fbba9da380a8b8a576['h0402c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02017] =  I8a0037ad2845a3fbba9da380a8b8a576['h0402e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02018] =  I8a0037ad2845a3fbba9da380a8b8a576['h04030] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02019] =  I8a0037ad2845a3fbba9da380a8b8a576['h04032] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0201a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04034] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0201b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04036] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0201c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04038] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0201d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0403a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0201e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0403c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0201f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0403e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02020] =  I8a0037ad2845a3fbba9da380a8b8a576['h04040] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02021] =  I8a0037ad2845a3fbba9da380a8b8a576['h04042] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02022] =  I8a0037ad2845a3fbba9da380a8b8a576['h04044] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02023] =  I8a0037ad2845a3fbba9da380a8b8a576['h04046] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02024] =  I8a0037ad2845a3fbba9da380a8b8a576['h04048] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02025] =  I8a0037ad2845a3fbba9da380a8b8a576['h0404a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02026] =  I8a0037ad2845a3fbba9da380a8b8a576['h0404c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02027] =  I8a0037ad2845a3fbba9da380a8b8a576['h0404e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02028] =  I8a0037ad2845a3fbba9da380a8b8a576['h04050] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02029] =  I8a0037ad2845a3fbba9da380a8b8a576['h04052] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0202a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04054] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0202b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04056] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0202c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04058] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0202d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0405a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0202e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0405c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0202f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0405e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02030] =  I8a0037ad2845a3fbba9da380a8b8a576['h04060] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02031] =  I8a0037ad2845a3fbba9da380a8b8a576['h04062] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02032] =  I8a0037ad2845a3fbba9da380a8b8a576['h04064] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02033] =  I8a0037ad2845a3fbba9da380a8b8a576['h04066] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02034] =  I8a0037ad2845a3fbba9da380a8b8a576['h04068] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02035] =  I8a0037ad2845a3fbba9da380a8b8a576['h0406a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02036] =  I8a0037ad2845a3fbba9da380a8b8a576['h0406c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02037] =  I8a0037ad2845a3fbba9da380a8b8a576['h0406e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02038] =  I8a0037ad2845a3fbba9da380a8b8a576['h04070] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02039] =  I8a0037ad2845a3fbba9da380a8b8a576['h04072] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0203a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04074] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0203b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04076] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0203c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04078] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0203d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0407a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0203e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0407c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0203f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0407e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02040] =  I8a0037ad2845a3fbba9da380a8b8a576['h04080] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02041] =  I8a0037ad2845a3fbba9da380a8b8a576['h04082] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02042] =  I8a0037ad2845a3fbba9da380a8b8a576['h04084] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02043] =  I8a0037ad2845a3fbba9da380a8b8a576['h04086] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02044] =  I8a0037ad2845a3fbba9da380a8b8a576['h04088] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02045] =  I8a0037ad2845a3fbba9da380a8b8a576['h0408a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02046] =  I8a0037ad2845a3fbba9da380a8b8a576['h0408c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02047] =  I8a0037ad2845a3fbba9da380a8b8a576['h0408e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02048] =  I8a0037ad2845a3fbba9da380a8b8a576['h04090] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02049] =  I8a0037ad2845a3fbba9da380a8b8a576['h04092] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0204a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04094] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0204b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04096] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0204c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04098] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0204d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0409a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0204e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0409c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0204f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0409e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02050] =  I8a0037ad2845a3fbba9da380a8b8a576['h040a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02051] =  I8a0037ad2845a3fbba9da380a8b8a576['h040a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02052] =  I8a0037ad2845a3fbba9da380a8b8a576['h040a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02053] =  I8a0037ad2845a3fbba9da380a8b8a576['h040a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02054] =  I8a0037ad2845a3fbba9da380a8b8a576['h040a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02055] =  I8a0037ad2845a3fbba9da380a8b8a576['h040aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02056] =  I8a0037ad2845a3fbba9da380a8b8a576['h040ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02057] =  I8a0037ad2845a3fbba9da380a8b8a576['h040ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02058] =  I8a0037ad2845a3fbba9da380a8b8a576['h040b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02059] =  I8a0037ad2845a3fbba9da380a8b8a576['h040b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0205a] =  I8a0037ad2845a3fbba9da380a8b8a576['h040b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0205b] =  I8a0037ad2845a3fbba9da380a8b8a576['h040b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0205c] =  I8a0037ad2845a3fbba9da380a8b8a576['h040b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0205d] =  I8a0037ad2845a3fbba9da380a8b8a576['h040ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0205e] =  I8a0037ad2845a3fbba9da380a8b8a576['h040bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0205f] =  I8a0037ad2845a3fbba9da380a8b8a576['h040be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02060] =  I8a0037ad2845a3fbba9da380a8b8a576['h040c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02061] =  I8a0037ad2845a3fbba9da380a8b8a576['h040c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02062] =  I8a0037ad2845a3fbba9da380a8b8a576['h040c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02063] =  I8a0037ad2845a3fbba9da380a8b8a576['h040c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02064] =  I8a0037ad2845a3fbba9da380a8b8a576['h040c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02065] =  I8a0037ad2845a3fbba9da380a8b8a576['h040ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02066] =  I8a0037ad2845a3fbba9da380a8b8a576['h040cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02067] =  I8a0037ad2845a3fbba9da380a8b8a576['h040ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02068] =  I8a0037ad2845a3fbba9da380a8b8a576['h040d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02069] =  I8a0037ad2845a3fbba9da380a8b8a576['h040d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0206a] =  I8a0037ad2845a3fbba9da380a8b8a576['h040d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0206b] =  I8a0037ad2845a3fbba9da380a8b8a576['h040d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0206c] =  I8a0037ad2845a3fbba9da380a8b8a576['h040d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0206d] =  I8a0037ad2845a3fbba9da380a8b8a576['h040da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0206e] =  I8a0037ad2845a3fbba9da380a8b8a576['h040dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0206f] =  I8a0037ad2845a3fbba9da380a8b8a576['h040de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02070] =  I8a0037ad2845a3fbba9da380a8b8a576['h040e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02071] =  I8a0037ad2845a3fbba9da380a8b8a576['h040e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02072] =  I8a0037ad2845a3fbba9da380a8b8a576['h040e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02073] =  I8a0037ad2845a3fbba9da380a8b8a576['h040e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02074] =  I8a0037ad2845a3fbba9da380a8b8a576['h040e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02075] =  I8a0037ad2845a3fbba9da380a8b8a576['h040ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02076] =  I8a0037ad2845a3fbba9da380a8b8a576['h040ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02077] =  I8a0037ad2845a3fbba9da380a8b8a576['h040ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02078] =  I8a0037ad2845a3fbba9da380a8b8a576['h040f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02079] =  I8a0037ad2845a3fbba9da380a8b8a576['h040f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0207a] =  I8a0037ad2845a3fbba9da380a8b8a576['h040f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0207b] =  I8a0037ad2845a3fbba9da380a8b8a576['h040f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0207c] =  I8a0037ad2845a3fbba9da380a8b8a576['h040f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0207d] =  I8a0037ad2845a3fbba9da380a8b8a576['h040fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0207e] =  I8a0037ad2845a3fbba9da380a8b8a576['h040fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0207f] =  I8a0037ad2845a3fbba9da380a8b8a576['h040fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02080] =  I8a0037ad2845a3fbba9da380a8b8a576['h04100] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02081] =  I8a0037ad2845a3fbba9da380a8b8a576['h04102] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02082] =  I8a0037ad2845a3fbba9da380a8b8a576['h04104] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02083] =  I8a0037ad2845a3fbba9da380a8b8a576['h04106] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02084] =  I8a0037ad2845a3fbba9da380a8b8a576['h04108] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02085] =  I8a0037ad2845a3fbba9da380a8b8a576['h0410a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02086] =  I8a0037ad2845a3fbba9da380a8b8a576['h0410c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02087] =  I8a0037ad2845a3fbba9da380a8b8a576['h0410e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02088] =  I8a0037ad2845a3fbba9da380a8b8a576['h04110] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02089] =  I8a0037ad2845a3fbba9da380a8b8a576['h04112] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0208a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04114] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0208b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04116] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0208c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04118] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0208d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0411a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0208e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0411c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0208f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0411e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02090] =  I8a0037ad2845a3fbba9da380a8b8a576['h04120] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02091] =  I8a0037ad2845a3fbba9da380a8b8a576['h04122] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02092] =  I8a0037ad2845a3fbba9da380a8b8a576['h04124] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02093] =  I8a0037ad2845a3fbba9da380a8b8a576['h04126] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02094] =  I8a0037ad2845a3fbba9da380a8b8a576['h04128] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02095] =  I8a0037ad2845a3fbba9da380a8b8a576['h0412a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02096] =  I8a0037ad2845a3fbba9da380a8b8a576['h0412c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02097] =  I8a0037ad2845a3fbba9da380a8b8a576['h0412e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02098] =  I8a0037ad2845a3fbba9da380a8b8a576['h04130] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02099] =  I8a0037ad2845a3fbba9da380a8b8a576['h04132] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0209a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04134] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0209b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04136] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0209c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04138] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0209d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0413a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0209e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0413c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0209f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0413e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04140] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04142] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04144] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04146] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04148] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0414a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0414c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0414e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04150] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04152] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h04154] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h04156] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h04158] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0415a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0415c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020af] =  I8a0037ad2845a3fbba9da380a8b8a576['h0415e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04160] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04162] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04164] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04166] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04168] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0416a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0416c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0416e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04170] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04172] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h04174] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h04176] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h04178] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0417a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020be] =  I8a0037ad2845a3fbba9da380a8b8a576['h0417c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0417e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04180] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04182] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04184] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04186] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04188] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0418a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0418c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0418e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04190] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04192] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h04194] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h04196] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h04198] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0419a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0419c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0419e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h041a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h041a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h041a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h041a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h041a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h041aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h041ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h041ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h041b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h041b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020da] =  I8a0037ad2845a3fbba9da380a8b8a576['h041b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020db] =  I8a0037ad2845a3fbba9da380a8b8a576['h041b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h041b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h041ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020de] =  I8a0037ad2845a3fbba9da380a8b8a576['h041bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020df] =  I8a0037ad2845a3fbba9da380a8b8a576['h041be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h041c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h041c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h041c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h041c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h041c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h041ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h041cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h041ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h041d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h041d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h041d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h041d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h041d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h041da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h041dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h041de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h041e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h041e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h041e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h041e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h041e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h041ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h041ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h041ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h041f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h041f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h041f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h041f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h041f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h041fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h041fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h020ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h041fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02100] =  I8a0037ad2845a3fbba9da380a8b8a576['h04200] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02101] =  I8a0037ad2845a3fbba9da380a8b8a576['h04202] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02102] =  I8a0037ad2845a3fbba9da380a8b8a576['h04204] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02103] =  I8a0037ad2845a3fbba9da380a8b8a576['h04206] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02104] =  I8a0037ad2845a3fbba9da380a8b8a576['h04208] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02105] =  I8a0037ad2845a3fbba9da380a8b8a576['h0420a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02106] =  I8a0037ad2845a3fbba9da380a8b8a576['h0420c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02107] =  I8a0037ad2845a3fbba9da380a8b8a576['h0420e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02108] =  I8a0037ad2845a3fbba9da380a8b8a576['h04210] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02109] =  I8a0037ad2845a3fbba9da380a8b8a576['h04212] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0210a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04214] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0210b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04216] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0210c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04218] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0210d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0421a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0210e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0421c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0210f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0421e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02110] =  I8a0037ad2845a3fbba9da380a8b8a576['h04220] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02111] =  I8a0037ad2845a3fbba9da380a8b8a576['h04222] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02112] =  I8a0037ad2845a3fbba9da380a8b8a576['h04224] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02113] =  I8a0037ad2845a3fbba9da380a8b8a576['h04226] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02114] =  I8a0037ad2845a3fbba9da380a8b8a576['h04228] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02115] =  I8a0037ad2845a3fbba9da380a8b8a576['h0422a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02116] =  I8a0037ad2845a3fbba9da380a8b8a576['h0422c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02117] =  I8a0037ad2845a3fbba9da380a8b8a576['h0422e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02118] =  I8a0037ad2845a3fbba9da380a8b8a576['h04230] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02119] =  I8a0037ad2845a3fbba9da380a8b8a576['h04232] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0211a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04234] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0211b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04236] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0211c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04238] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0211d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0423a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0211e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0423c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0211f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0423e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02120] =  I8a0037ad2845a3fbba9da380a8b8a576['h04240] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02121] =  I8a0037ad2845a3fbba9da380a8b8a576['h04242] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02122] =  I8a0037ad2845a3fbba9da380a8b8a576['h04244] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02123] =  I8a0037ad2845a3fbba9da380a8b8a576['h04246] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02124] =  I8a0037ad2845a3fbba9da380a8b8a576['h04248] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02125] =  I8a0037ad2845a3fbba9da380a8b8a576['h0424a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02126] =  I8a0037ad2845a3fbba9da380a8b8a576['h0424c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02127] =  I8a0037ad2845a3fbba9da380a8b8a576['h0424e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02128] =  I8a0037ad2845a3fbba9da380a8b8a576['h04250] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02129] =  I8a0037ad2845a3fbba9da380a8b8a576['h04252] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0212a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04254] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0212b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04256] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0212c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04258] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0212d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0425a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0212e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0425c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0212f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0425e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02130] =  I8a0037ad2845a3fbba9da380a8b8a576['h04260] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02131] =  I8a0037ad2845a3fbba9da380a8b8a576['h04262] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02132] =  I8a0037ad2845a3fbba9da380a8b8a576['h04264] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02133] =  I8a0037ad2845a3fbba9da380a8b8a576['h04266] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02134] =  I8a0037ad2845a3fbba9da380a8b8a576['h04268] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02135] =  I8a0037ad2845a3fbba9da380a8b8a576['h0426a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02136] =  I8a0037ad2845a3fbba9da380a8b8a576['h0426c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02137] =  I8a0037ad2845a3fbba9da380a8b8a576['h0426e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02138] =  I8a0037ad2845a3fbba9da380a8b8a576['h04270] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02139] =  I8a0037ad2845a3fbba9da380a8b8a576['h04272] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0213a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04274] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0213b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04276] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0213c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04278] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0213d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0427a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0213e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0427c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0213f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0427e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02140] =  I8a0037ad2845a3fbba9da380a8b8a576['h04280] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02141] =  I8a0037ad2845a3fbba9da380a8b8a576['h04282] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02142] =  I8a0037ad2845a3fbba9da380a8b8a576['h04284] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02143] =  I8a0037ad2845a3fbba9da380a8b8a576['h04286] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02144] =  I8a0037ad2845a3fbba9da380a8b8a576['h04288] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02145] =  I8a0037ad2845a3fbba9da380a8b8a576['h0428a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02146] =  I8a0037ad2845a3fbba9da380a8b8a576['h0428c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02147] =  I8a0037ad2845a3fbba9da380a8b8a576['h0428e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02148] =  I8a0037ad2845a3fbba9da380a8b8a576['h04290] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02149] =  I8a0037ad2845a3fbba9da380a8b8a576['h04292] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0214a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04294] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0214b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04296] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0214c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04298] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0214d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0429a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0214e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0429c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0214f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0429e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02150] =  I8a0037ad2845a3fbba9da380a8b8a576['h042a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02151] =  I8a0037ad2845a3fbba9da380a8b8a576['h042a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02152] =  I8a0037ad2845a3fbba9da380a8b8a576['h042a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02153] =  I8a0037ad2845a3fbba9da380a8b8a576['h042a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02154] =  I8a0037ad2845a3fbba9da380a8b8a576['h042a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02155] =  I8a0037ad2845a3fbba9da380a8b8a576['h042aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02156] =  I8a0037ad2845a3fbba9da380a8b8a576['h042ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02157] =  I8a0037ad2845a3fbba9da380a8b8a576['h042ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02158] =  I8a0037ad2845a3fbba9da380a8b8a576['h042b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02159] =  I8a0037ad2845a3fbba9da380a8b8a576['h042b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0215a] =  I8a0037ad2845a3fbba9da380a8b8a576['h042b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0215b] =  I8a0037ad2845a3fbba9da380a8b8a576['h042b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0215c] =  I8a0037ad2845a3fbba9da380a8b8a576['h042b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0215d] =  I8a0037ad2845a3fbba9da380a8b8a576['h042ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0215e] =  I8a0037ad2845a3fbba9da380a8b8a576['h042bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0215f] =  I8a0037ad2845a3fbba9da380a8b8a576['h042be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02160] =  I8a0037ad2845a3fbba9da380a8b8a576['h042c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02161] =  I8a0037ad2845a3fbba9da380a8b8a576['h042c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02162] =  I8a0037ad2845a3fbba9da380a8b8a576['h042c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02163] =  I8a0037ad2845a3fbba9da380a8b8a576['h042c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02164] =  I8a0037ad2845a3fbba9da380a8b8a576['h042c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02165] =  I8a0037ad2845a3fbba9da380a8b8a576['h042ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02166] =  I8a0037ad2845a3fbba9da380a8b8a576['h042cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02167] =  I8a0037ad2845a3fbba9da380a8b8a576['h042ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02168] =  I8a0037ad2845a3fbba9da380a8b8a576['h042d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02169] =  I8a0037ad2845a3fbba9da380a8b8a576['h042d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0216a] =  I8a0037ad2845a3fbba9da380a8b8a576['h042d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0216b] =  I8a0037ad2845a3fbba9da380a8b8a576['h042d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0216c] =  I8a0037ad2845a3fbba9da380a8b8a576['h042d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0216d] =  I8a0037ad2845a3fbba9da380a8b8a576['h042da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0216e] =  I8a0037ad2845a3fbba9da380a8b8a576['h042dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0216f] =  I8a0037ad2845a3fbba9da380a8b8a576['h042de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02170] =  I8a0037ad2845a3fbba9da380a8b8a576['h042e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02171] =  I8a0037ad2845a3fbba9da380a8b8a576['h042e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02172] =  I8a0037ad2845a3fbba9da380a8b8a576['h042e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02173] =  I8a0037ad2845a3fbba9da380a8b8a576['h042e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02174] =  I8a0037ad2845a3fbba9da380a8b8a576['h042e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02175] =  I8a0037ad2845a3fbba9da380a8b8a576['h042ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02176] =  I8a0037ad2845a3fbba9da380a8b8a576['h042ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02177] =  I8a0037ad2845a3fbba9da380a8b8a576['h042ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02178] =  I8a0037ad2845a3fbba9da380a8b8a576['h042f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02179] =  I8a0037ad2845a3fbba9da380a8b8a576['h042f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0217a] =  I8a0037ad2845a3fbba9da380a8b8a576['h042f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0217b] =  I8a0037ad2845a3fbba9da380a8b8a576['h042f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0217c] =  I8a0037ad2845a3fbba9da380a8b8a576['h042f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0217d] =  I8a0037ad2845a3fbba9da380a8b8a576['h042fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0217e] =  I8a0037ad2845a3fbba9da380a8b8a576['h042fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0217f] =  I8a0037ad2845a3fbba9da380a8b8a576['h042fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02180] =  I8a0037ad2845a3fbba9da380a8b8a576['h04300] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02181] =  I8a0037ad2845a3fbba9da380a8b8a576['h04302] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02182] =  I8a0037ad2845a3fbba9da380a8b8a576['h04304] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02183] =  I8a0037ad2845a3fbba9da380a8b8a576['h04306] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02184] =  I8a0037ad2845a3fbba9da380a8b8a576['h04308] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02185] =  I8a0037ad2845a3fbba9da380a8b8a576['h0430a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02186] =  I8a0037ad2845a3fbba9da380a8b8a576['h0430c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02187] =  I8a0037ad2845a3fbba9da380a8b8a576['h0430e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02188] =  I8a0037ad2845a3fbba9da380a8b8a576['h04310] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02189] =  I8a0037ad2845a3fbba9da380a8b8a576['h04312] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0218a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04314] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0218b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04316] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0218c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04318] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0218d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0431a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0218e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0431c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0218f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0431e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02190] =  I8a0037ad2845a3fbba9da380a8b8a576['h04320] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02191] =  I8a0037ad2845a3fbba9da380a8b8a576['h04322] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02192] =  I8a0037ad2845a3fbba9da380a8b8a576['h04324] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02193] =  I8a0037ad2845a3fbba9da380a8b8a576['h04326] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02194] =  I8a0037ad2845a3fbba9da380a8b8a576['h04328] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02195] =  I8a0037ad2845a3fbba9da380a8b8a576['h0432a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02196] =  I8a0037ad2845a3fbba9da380a8b8a576['h0432c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02197] =  I8a0037ad2845a3fbba9da380a8b8a576['h0432e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02198] =  I8a0037ad2845a3fbba9da380a8b8a576['h04330] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02199] =  I8a0037ad2845a3fbba9da380a8b8a576['h04332] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0219a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04334] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0219b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04336] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0219c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04338] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0219d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0433a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0219e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0433c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0219f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0433e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04340] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04342] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04344] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04346] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04348] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0434a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0434c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0434e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04350] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04352] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h04354] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h04356] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h04358] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0435a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0435c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021af] =  I8a0037ad2845a3fbba9da380a8b8a576['h0435e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04360] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04362] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04364] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04366] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04368] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0436a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0436c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0436e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04370] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04372] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h04374] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h04376] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h04378] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0437a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021be] =  I8a0037ad2845a3fbba9da380a8b8a576['h0437c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0437e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04380] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04382] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04384] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04386] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04388] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0438a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0438c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0438e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04390] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04392] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h04394] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h04396] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h04398] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0439a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0439c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0439e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h043a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h043a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h043a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h043a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h043a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h043aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h043ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h043ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h043b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h043b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021da] =  I8a0037ad2845a3fbba9da380a8b8a576['h043b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021db] =  I8a0037ad2845a3fbba9da380a8b8a576['h043b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h043b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h043ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021de] =  I8a0037ad2845a3fbba9da380a8b8a576['h043bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021df] =  I8a0037ad2845a3fbba9da380a8b8a576['h043be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h043c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h043c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h043c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h043c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h043c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h043ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h043cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h043ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h043d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h043d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h043d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h043d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h043d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h043da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h043dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h043de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h043e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h043e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h043e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h043e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h043e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h043ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h043ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h043ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h043f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h043f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h043f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h043f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h043f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h043fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h043fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h021ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h043fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02200] =  I8a0037ad2845a3fbba9da380a8b8a576['h04400] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02201] =  I8a0037ad2845a3fbba9da380a8b8a576['h04402] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02202] =  I8a0037ad2845a3fbba9da380a8b8a576['h04404] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02203] =  I8a0037ad2845a3fbba9da380a8b8a576['h04406] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02204] =  I8a0037ad2845a3fbba9da380a8b8a576['h04408] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02205] =  I8a0037ad2845a3fbba9da380a8b8a576['h0440a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02206] =  I8a0037ad2845a3fbba9da380a8b8a576['h0440c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02207] =  I8a0037ad2845a3fbba9da380a8b8a576['h0440e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02208] =  I8a0037ad2845a3fbba9da380a8b8a576['h04410] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02209] =  I8a0037ad2845a3fbba9da380a8b8a576['h04412] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0220a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04414] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0220b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04416] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0220c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04418] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0220d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0441a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0220e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0441c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0220f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0441e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02210] =  I8a0037ad2845a3fbba9da380a8b8a576['h04420] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02211] =  I8a0037ad2845a3fbba9da380a8b8a576['h04422] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02212] =  I8a0037ad2845a3fbba9da380a8b8a576['h04424] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02213] =  I8a0037ad2845a3fbba9da380a8b8a576['h04426] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02214] =  I8a0037ad2845a3fbba9da380a8b8a576['h04428] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02215] =  I8a0037ad2845a3fbba9da380a8b8a576['h0442a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02216] =  I8a0037ad2845a3fbba9da380a8b8a576['h0442c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02217] =  I8a0037ad2845a3fbba9da380a8b8a576['h0442e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02218] =  I8a0037ad2845a3fbba9da380a8b8a576['h04430] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02219] =  I8a0037ad2845a3fbba9da380a8b8a576['h04432] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0221a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04434] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0221b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04436] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0221c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04438] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0221d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0443a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0221e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0443c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0221f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0443e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02220] =  I8a0037ad2845a3fbba9da380a8b8a576['h04440] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02221] =  I8a0037ad2845a3fbba9da380a8b8a576['h04442] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02222] =  I8a0037ad2845a3fbba9da380a8b8a576['h04444] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02223] =  I8a0037ad2845a3fbba9da380a8b8a576['h04446] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02224] =  I8a0037ad2845a3fbba9da380a8b8a576['h04448] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02225] =  I8a0037ad2845a3fbba9da380a8b8a576['h0444a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02226] =  I8a0037ad2845a3fbba9da380a8b8a576['h0444c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02227] =  I8a0037ad2845a3fbba9da380a8b8a576['h0444e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02228] =  I8a0037ad2845a3fbba9da380a8b8a576['h04450] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02229] =  I8a0037ad2845a3fbba9da380a8b8a576['h04452] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0222a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04454] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0222b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04456] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0222c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04458] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0222d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0445a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0222e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0445c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0222f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0445e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02230] =  I8a0037ad2845a3fbba9da380a8b8a576['h04460] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02231] =  I8a0037ad2845a3fbba9da380a8b8a576['h04462] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02232] =  I8a0037ad2845a3fbba9da380a8b8a576['h04464] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02233] =  I8a0037ad2845a3fbba9da380a8b8a576['h04466] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02234] =  I8a0037ad2845a3fbba9da380a8b8a576['h04468] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02235] =  I8a0037ad2845a3fbba9da380a8b8a576['h0446a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02236] =  I8a0037ad2845a3fbba9da380a8b8a576['h0446c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02237] =  I8a0037ad2845a3fbba9da380a8b8a576['h0446e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02238] =  I8a0037ad2845a3fbba9da380a8b8a576['h04470] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02239] =  I8a0037ad2845a3fbba9da380a8b8a576['h04472] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0223a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04474] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0223b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04476] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0223c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04478] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0223d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0447a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0223e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0447c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0223f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0447e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02240] =  I8a0037ad2845a3fbba9da380a8b8a576['h04480] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02241] =  I8a0037ad2845a3fbba9da380a8b8a576['h04482] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02242] =  I8a0037ad2845a3fbba9da380a8b8a576['h04484] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02243] =  I8a0037ad2845a3fbba9da380a8b8a576['h04486] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02244] =  I8a0037ad2845a3fbba9da380a8b8a576['h04488] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02245] =  I8a0037ad2845a3fbba9da380a8b8a576['h0448a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02246] =  I8a0037ad2845a3fbba9da380a8b8a576['h0448c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02247] =  I8a0037ad2845a3fbba9da380a8b8a576['h0448e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02248] =  I8a0037ad2845a3fbba9da380a8b8a576['h04490] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02249] =  I8a0037ad2845a3fbba9da380a8b8a576['h04492] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0224a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04494] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0224b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04496] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0224c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04498] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0224d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0449a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0224e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0449c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0224f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0449e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02250] =  I8a0037ad2845a3fbba9da380a8b8a576['h044a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02251] =  I8a0037ad2845a3fbba9da380a8b8a576['h044a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02252] =  I8a0037ad2845a3fbba9da380a8b8a576['h044a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02253] =  I8a0037ad2845a3fbba9da380a8b8a576['h044a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02254] =  I8a0037ad2845a3fbba9da380a8b8a576['h044a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02255] =  I8a0037ad2845a3fbba9da380a8b8a576['h044aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02256] =  I8a0037ad2845a3fbba9da380a8b8a576['h044ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02257] =  I8a0037ad2845a3fbba9da380a8b8a576['h044ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02258] =  I8a0037ad2845a3fbba9da380a8b8a576['h044b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02259] =  I8a0037ad2845a3fbba9da380a8b8a576['h044b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0225a] =  I8a0037ad2845a3fbba9da380a8b8a576['h044b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0225b] =  I8a0037ad2845a3fbba9da380a8b8a576['h044b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0225c] =  I8a0037ad2845a3fbba9da380a8b8a576['h044b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0225d] =  I8a0037ad2845a3fbba9da380a8b8a576['h044ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0225e] =  I8a0037ad2845a3fbba9da380a8b8a576['h044bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0225f] =  I8a0037ad2845a3fbba9da380a8b8a576['h044be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02260] =  I8a0037ad2845a3fbba9da380a8b8a576['h044c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02261] =  I8a0037ad2845a3fbba9da380a8b8a576['h044c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02262] =  I8a0037ad2845a3fbba9da380a8b8a576['h044c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02263] =  I8a0037ad2845a3fbba9da380a8b8a576['h044c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02264] =  I8a0037ad2845a3fbba9da380a8b8a576['h044c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02265] =  I8a0037ad2845a3fbba9da380a8b8a576['h044ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02266] =  I8a0037ad2845a3fbba9da380a8b8a576['h044cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02267] =  I8a0037ad2845a3fbba9da380a8b8a576['h044ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02268] =  I8a0037ad2845a3fbba9da380a8b8a576['h044d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02269] =  I8a0037ad2845a3fbba9da380a8b8a576['h044d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0226a] =  I8a0037ad2845a3fbba9da380a8b8a576['h044d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0226b] =  I8a0037ad2845a3fbba9da380a8b8a576['h044d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0226c] =  I8a0037ad2845a3fbba9da380a8b8a576['h044d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0226d] =  I8a0037ad2845a3fbba9da380a8b8a576['h044da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0226e] =  I8a0037ad2845a3fbba9da380a8b8a576['h044dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0226f] =  I8a0037ad2845a3fbba9da380a8b8a576['h044de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02270] =  I8a0037ad2845a3fbba9da380a8b8a576['h044e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02271] =  I8a0037ad2845a3fbba9da380a8b8a576['h044e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02272] =  I8a0037ad2845a3fbba9da380a8b8a576['h044e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02273] =  I8a0037ad2845a3fbba9da380a8b8a576['h044e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02274] =  I8a0037ad2845a3fbba9da380a8b8a576['h044e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02275] =  I8a0037ad2845a3fbba9da380a8b8a576['h044ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02276] =  I8a0037ad2845a3fbba9da380a8b8a576['h044ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02277] =  I8a0037ad2845a3fbba9da380a8b8a576['h044ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02278] =  I8a0037ad2845a3fbba9da380a8b8a576['h044f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02279] =  I8a0037ad2845a3fbba9da380a8b8a576['h044f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0227a] =  I8a0037ad2845a3fbba9da380a8b8a576['h044f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0227b] =  I8a0037ad2845a3fbba9da380a8b8a576['h044f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0227c] =  I8a0037ad2845a3fbba9da380a8b8a576['h044f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0227d] =  I8a0037ad2845a3fbba9da380a8b8a576['h044fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0227e] =  I8a0037ad2845a3fbba9da380a8b8a576['h044fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0227f] =  I8a0037ad2845a3fbba9da380a8b8a576['h044fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02280] =  I8a0037ad2845a3fbba9da380a8b8a576['h04500] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02281] =  I8a0037ad2845a3fbba9da380a8b8a576['h04502] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02282] =  I8a0037ad2845a3fbba9da380a8b8a576['h04504] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02283] =  I8a0037ad2845a3fbba9da380a8b8a576['h04506] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02284] =  I8a0037ad2845a3fbba9da380a8b8a576['h04508] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02285] =  I8a0037ad2845a3fbba9da380a8b8a576['h0450a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02286] =  I8a0037ad2845a3fbba9da380a8b8a576['h0450c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02287] =  I8a0037ad2845a3fbba9da380a8b8a576['h0450e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02288] =  I8a0037ad2845a3fbba9da380a8b8a576['h04510] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02289] =  I8a0037ad2845a3fbba9da380a8b8a576['h04512] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0228a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04514] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0228b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04516] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0228c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04518] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0228d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0451a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0228e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0451c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0228f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0451e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02290] =  I8a0037ad2845a3fbba9da380a8b8a576['h04520] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02291] =  I8a0037ad2845a3fbba9da380a8b8a576['h04522] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02292] =  I8a0037ad2845a3fbba9da380a8b8a576['h04524] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02293] =  I8a0037ad2845a3fbba9da380a8b8a576['h04526] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02294] =  I8a0037ad2845a3fbba9da380a8b8a576['h04528] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02295] =  I8a0037ad2845a3fbba9da380a8b8a576['h0452a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02296] =  I8a0037ad2845a3fbba9da380a8b8a576['h0452c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02297] =  I8a0037ad2845a3fbba9da380a8b8a576['h0452e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02298] =  I8a0037ad2845a3fbba9da380a8b8a576['h04530] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02299] =  I8a0037ad2845a3fbba9da380a8b8a576['h04532] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0229a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04534] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0229b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04536] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0229c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04538] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0229d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0453a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0229e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0453c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0229f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0453e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04540] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04542] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04544] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04546] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04548] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0454a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0454c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0454e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04550] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04552] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h04554] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h04556] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h04558] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0455a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0455c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022af] =  I8a0037ad2845a3fbba9da380a8b8a576['h0455e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04560] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04562] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04564] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04566] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04568] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0456a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0456c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0456e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04570] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04572] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h04574] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h04576] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h04578] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0457a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022be] =  I8a0037ad2845a3fbba9da380a8b8a576['h0457c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0457e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04580] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04582] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04584] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04586] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04588] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0458a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0458c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0458e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04590] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04592] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h04594] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h04596] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h04598] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0459a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0459c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0459e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h045a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h045a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h045a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h045a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h045a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h045aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h045ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h045ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h045b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h045b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022da] =  I8a0037ad2845a3fbba9da380a8b8a576['h045b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022db] =  I8a0037ad2845a3fbba9da380a8b8a576['h045b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h045b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h045ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022de] =  I8a0037ad2845a3fbba9da380a8b8a576['h045bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022df] =  I8a0037ad2845a3fbba9da380a8b8a576['h045be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h045c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h045c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h045c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h045c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h045c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h045ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h045cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h045ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h045d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h045d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h045d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h045d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h045d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h045da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h045dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h045de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h045e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h045e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h045e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h045e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h045e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h045ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h045ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h045ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h045f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h045f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h045f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h045f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h045f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h045fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h045fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h022ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h045fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02300] =  I8a0037ad2845a3fbba9da380a8b8a576['h04600] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02301] =  I8a0037ad2845a3fbba9da380a8b8a576['h04602] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02302] =  I8a0037ad2845a3fbba9da380a8b8a576['h04604] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02303] =  I8a0037ad2845a3fbba9da380a8b8a576['h04606] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02304] =  I8a0037ad2845a3fbba9da380a8b8a576['h04608] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02305] =  I8a0037ad2845a3fbba9da380a8b8a576['h0460a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02306] =  I8a0037ad2845a3fbba9da380a8b8a576['h0460c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02307] =  I8a0037ad2845a3fbba9da380a8b8a576['h0460e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02308] =  I8a0037ad2845a3fbba9da380a8b8a576['h04610] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02309] =  I8a0037ad2845a3fbba9da380a8b8a576['h04612] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0230a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04614] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0230b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04616] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0230c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04618] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0230d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0461a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0230e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0461c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0230f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0461e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02310] =  I8a0037ad2845a3fbba9da380a8b8a576['h04620] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02311] =  I8a0037ad2845a3fbba9da380a8b8a576['h04622] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02312] =  I8a0037ad2845a3fbba9da380a8b8a576['h04624] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02313] =  I8a0037ad2845a3fbba9da380a8b8a576['h04626] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02314] =  I8a0037ad2845a3fbba9da380a8b8a576['h04628] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02315] =  I8a0037ad2845a3fbba9da380a8b8a576['h0462a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02316] =  I8a0037ad2845a3fbba9da380a8b8a576['h0462c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02317] =  I8a0037ad2845a3fbba9da380a8b8a576['h0462e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02318] =  I8a0037ad2845a3fbba9da380a8b8a576['h04630] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02319] =  I8a0037ad2845a3fbba9da380a8b8a576['h04632] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0231a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04634] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0231b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04636] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0231c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04638] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0231d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0463a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0231e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0463c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0231f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0463e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02320] =  I8a0037ad2845a3fbba9da380a8b8a576['h04640] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02321] =  I8a0037ad2845a3fbba9da380a8b8a576['h04642] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02322] =  I8a0037ad2845a3fbba9da380a8b8a576['h04644] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02323] =  I8a0037ad2845a3fbba9da380a8b8a576['h04646] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02324] =  I8a0037ad2845a3fbba9da380a8b8a576['h04648] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02325] =  I8a0037ad2845a3fbba9da380a8b8a576['h0464a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02326] =  I8a0037ad2845a3fbba9da380a8b8a576['h0464c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02327] =  I8a0037ad2845a3fbba9da380a8b8a576['h0464e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02328] =  I8a0037ad2845a3fbba9da380a8b8a576['h04650] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02329] =  I8a0037ad2845a3fbba9da380a8b8a576['h04652] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0232a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04654] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0232b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04656] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0232c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04658] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0232d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0465a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0232e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0465c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0232f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0465e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02330] =  I8a0037ad2845a3fbba9da380a8b8a576['h04660] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02331] =  I8a0037ad2845a3fbba9da380a8b8a576['h04662] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02332] =  I8a0037ad2845a3fbba9da380a8b8a576['h04664] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02333] =  I8a0037ad2845a3fbba9da380a8b8a576['h04666] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02334] =  I8a0037ad2845a3fbba9da380a8b8a576['h04668] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02335] =  I8a0037ad2845a3fbba9da380a8b8a576['h0466a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02336] =  I8a0037ad2845a3fbba9da380a8b8a576['h0466c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02337] =  I8a0037ad2845a3fbba9da380a8b8a576['h0466e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02338] =  I8a0037ad2845a3fbba9da380a8b8a576['h04670] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02339] =  I8a0037ad2845a3fbba9da380a8b8a576['h04672] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0233a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04674] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0233b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04676] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0233c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04678] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0233d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0467a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0233e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0467c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0233f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0467e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02340] =  I8a0037ad2845a3fbba9da380a8b8a576['h04680] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02341] =  I8a0037ad2845a3fbba9da380a8b8a576['h04682] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02342] =  I8a0037ad2845a3fbba9da380a8b8a576['h04684] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02343] =  I8a0037ad2845a3fbba9da380a8b8a576['h04686] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02344] =  I8a0037ad2845a3fbba9da380a8b8a576['h04688] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02345] =  I8a0037ad2845a3fbba9da380a8b8a576['h0468a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02346] =  I8a0037ad2845a3fbba9da380a8b8a576['h0468c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02347] =  I8a0037ad2845a3fbba9da380a8b8a576['h0468e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02348] =  I8a0037ad2845a3fbba9da380a8b8a576['h04690] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02349] =  I8a0037ad2845a3fbba9da380a8b8a576['h04692] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0234a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04694] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0234b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04696] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0234c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04698] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0234d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0469a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0234e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0469c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0234f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0469e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02350] =  I8a0037ad2845a3fbba9da380a8b8a576['h046a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02351] =  I8a0037ad2845a3fbba9da380a8b8a576['h046a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02352] =  I8a0037ad2845a3fbba9da380a8b8a576['h046a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02353] =  I8a0037ad2845a3fbba9da380a8b8a576['h046a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02354] =  I8a0037ad2845a3fbba9da380a8b8a576['h046a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02355] =  I8a0037ad2845a3fbba9da380a8b8a576['h046aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02356] =  I8a0037ad2845a3fbba9da380a8b8a576['h046ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02357] =  I8a0037ad2845a3fbba9da380a8b8a576['h046ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02358] =  I8a0037ad2845a3fbba9da380a8b8a576['h046b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02359] =  I8a0037ad2845a3fbba9da380a8b8a576['h046b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0235a] =  I8a0037ad2845a3fbba9da380a8b8a576['h046b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0235b] =  I8a0037ad2845a3fbba9da380a8b8a576['h046b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0235c] =  I8a0037ad2845a3fbba9da380a8b8a576['h046b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0235d] =  I8a0037ad2845a3fbba9da380a8b8a576['h046ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0235e] =  I8a0037ad2845a3fbba9da380a8b8a576['h046bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0235f] =  I8a0037ad2845a3fbba9da380a8b8a576['h046be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02360] =  I8a0037ad2845a3fbba9da380a8b8a576['h046c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02361] =  I8a0037ad2845a3fbba9da380a8b8a576['h046c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02362] =  I8a0037ad2845a3fbba9da380a8b8a576['h046c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02363] =  I8a0037ad2845a3fbba9da380a8b8a576['h046c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02364] =  I8a0037ad2845a3fbba9da380a8b8a576['h046c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02365] =  I8a0037ad2845a3fbba9da380a8b8a576['h046ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02366] =  I8a0037ad2845a3fbba9da380a8b8a576['h046cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02367] =  I8a0037ad2845a3fbba9da380a8b8a576['h046ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02368] =  I8a0037ad2845a3fbba9da380a8b8a576['h046d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02369] =  I8a0037ad2845a3fbba9da380a8b8a576['h046d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0236a] =  I8a0037ad2845a3fbba9da380a8b8a576['h046d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0236b] =  I8a0037ad2845a3fbba9da380a8b8a576['h046d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0236c] =  I8a0037ad2845a3fbba9da380a8b8a576['h046d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0236d] =  I8a0037ad2845a3fbba9da380a8b8a576['h046da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0236e] =  I8a0037ad2845a3fbba9da380a8b8a576['h046dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0236f] =  I8a0037ad2845a3fbba9da380a8b8a576['h046de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02370] =  I8a0037ad2845a3fbba9da380a8b8a576['h046e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02371] =  I8a0037ad2845a3fbba9da380a8b8a576['h046e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02372] =  I8a0037ad2845a3fbba9da380a8b8a576['h046e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02373] =  I8a0037ad2845a3fbba9da380a8b8a576['h046e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02374] =  I8a0037ad2845a3fbba9da380a8b8a576['h046e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02375] =  I8a0037ad2845a3fbba9da380a8b8a576['h046ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02376] =  I8a0037ad2845a3fbba9da380a8b8a576['h046ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02377] =  I8a0037ad2845a3fbba9da380a8b8a576['h046ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02378] =  I8a0037ad2845a3fbba9da380a8b8a576['h046f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02379] =  I8a0037ad2845a3fbba9da380a8b8a576['h046f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0237a] =  I8a0037ad2845a3fbba9da380a8b8a576['h046f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0237b] =  I8a0037ad2845a3fbba9da380a8b8a576['h046f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0237c] =  I8a0037ad2845a3fbba9da380a8b8a576['h046f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0237d] =  I8a0037ad2845a3fbba9da380a8b8a576['h046fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0237e] =  I8a0037ad2845a3fbba9da380a8b8a576['h046fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0237f] =  I8a0037ad2845a3fbba9da380a8b8a576['h046fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02380] =  I8a0037ad2845a3fbba9da380a8b8a576['h04700] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02381] =  I8a0037ad2845a3fbba9da380a8b8a576['h04702] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02382] =  I8a0037ad2845a3fbba9da380a8b8a576['h04704] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02383] =  I8a0037ad2845a3fbba9da380a8b8a576['h04706] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02384] =  I8a0037ad2845a3fbba9da380a8b8a576['h04708] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02385] =  I8a0037ad2845a3fbba9da380a8b8a576['h0470a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02386] =  I8a0037ad2845a3fbba9da380a8b8a576['h0470c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02387] =  I8a0037ad2845a3fbba9da380a8b8a576['h0470e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02388] =  I8a0037ad2845a3fbba9da380a8b8a576['h04710] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02389] =  I8a0037ad2845a3fbba9da380a8b8a576['h04712] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0238a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04714] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0238b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04716] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0238c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04718] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0238d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0471a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0238e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0471c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0238f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0471e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02390] =  I8a0037ad2845a3fbba9da380a8b8a576['h04720] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02391] =  I8a0037ad2845a3fbba9da380a8b8a576['h04722] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02392] =  I8a0037ad2845a3fbba9da380a8b8a576['h04724] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02393] =  I8a0037ad2845a3fbba9da380a8b8a576['h04726] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02394] =  I8a0037ad2845a3fbba9da380a8b8a576['h04728] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02395] =  I8a0037ad2845a3fbba9da380a8b8a576['h0472a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02396] =  I8a0037ad2845a3fbba9da380a8b8a576['h0472c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02397] =  I8a0037ad2845a3fbba9da380a8b8a576['h0472e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02398] =  I8a0037ad2845a3fbba9da380a8b8a576['h04730] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02399] =  I8a0037ad2845a3fbba9da380a8b8a576['h04732] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0239a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04734] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0239b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04736] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0239c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04738] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0239d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0473a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0239e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0473c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0239f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0473e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04740] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04742] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04744] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04746] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04748] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0474a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0474c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0474e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04750] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04752] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h04754] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h04756] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h04758] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0475a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0475c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023af] =  I8a0037ad2845a3fbba9da380a8b8a576['h0475e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04760] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04762] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04764] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04766] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04768] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0476a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0476c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0476e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04770] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04772] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h04774] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h04776] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h04778] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0477a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023be] =  I8a0037ad2845a3fbba9da380a8b8a576['h0477c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0477e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04780] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04782] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04784] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04786] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04788] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0478a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0478c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0478e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04790] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04792] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h04794] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h04796] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h04798] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0479a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0479c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0479e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h047a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h047a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h047a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h047a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h047a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h047aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h047ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h047ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h047b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h047b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023da] =  I8a0037ad2845a3fbba9da380a8b8a576['h047b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023db] =  I8a0037ad2845a3fbba9da380a8b8a576['h047b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h047b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h047ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023de] =  I8a0037ad2845a3fbba9da380a8b8a576['h047bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023df] =  I8a0037ad2845a3fbba9da380a8b8a576['h047be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h047c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h047c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h047c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h047c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h047c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h047ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h047cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h047ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h047d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h047d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h047d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h047d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h047d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h047da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h047dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h047de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h047e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h047e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h047e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h047e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h047e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h047ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h047ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h047ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h047f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h047f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h047f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h047f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h047f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h047fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h047fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h023ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h047fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02400] =  I8a0037ad2845a3fbba9da380a8b8a576['h04800] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02401] =  I8a0037ad2845a3fbba9da380a8b8a576['h04802] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02402] =  I8a0037ad2845a3fbba9da380a8b8a576['h04804] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02403] =  I8a0037ad2845a3fbba9da380a8b8a576['h04806] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02404] =  I8a0037ad2845a3fbba9da380a8b8a576['h04808] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02405] =  I8a0037ad2845a3fbba9da380a8b8a576['h0480a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02406] =  I8a0037ad2845a3fbba9da380a8b8a576['h0480c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02407] =  I8a0037ad2845a3fbba9da380a8b8a576['h0480e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02408] =  I8a0037ad2845a3fbba9da380a8b8a576['h04810] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02409] =  I8a0037ad2845a3fbba9da380a8b8a576['h04812] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0240a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04814] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0240b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04816] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0240c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04818] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0240d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0481a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0240e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0481c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0240f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0481e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02410] =  I8a0037ad2845a3fbba9da380a8b8a576['h04820] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02411] =  I8a0037ad2845a3fbba9da380a8b8a576['h04822] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02412] =  I8a0037ad2845a3fbba9da380a8b8a576['h04824] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02413] =  I8a0037ad2845a3fbba9da380a8b8a576['h04826] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02414] =  I8a0037ad2845a3fbba9da380a8b8a576['h04828] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02415] =  I8a0037ad2845a3fbba9da380a8b8a576['h0482a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02416] =  I8a0037ad2845a3fbba9da380a8b8a576['h0482c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02417] =  I8a0037ad2845a3fbba9da380a8b8a576['h0482e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02418] =  I8a0037ad2845a3fbba9da380a8b8a576['h04830] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02419] =  I8a0037ad2845a3fbba9da380a8b8a576['h04832] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0241a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04834] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0241b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04836] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0241c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04838] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0241d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0483a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0241e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0483c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0241f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0483e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02420] =  I8a0037ad2845a3fbba9da380a8b8a576['h04840] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02421] =  I8a0037ad2845a3fbba9da380a8b8a576['h04842] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02422] =  I8a0037ad2845a3fbba9da380a8b8a576['h04844] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02423] =  I8a0037ad2845a3fbba9da380a8b8a576['h04846] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02424] =  I8a0037ad2845a3fbba9da380a8b8a576['h04848] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02425] =  I8a0037ad2845a3fbba9da380a8b8a576['h0484a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02426] =  I8a0037ad2845a3fbba9da380a8b8a576['h0484c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02427] =  I8a0037ad2845a3fbba9da380a8b8a576['h0484e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02428] =  I8a0037ad2845a3fbba9da380a8b8a576['h04850] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02429] =  I8a0037ad2845a3fbba9da380a8b8a576['h04852] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0242a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04854] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0242b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04856] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0242c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04858] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0242d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0485a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0242e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0485c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0242f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0485e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02430] =  I8a0037ad2845a3fbba9da380a8b8a576['h04860] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02431] =  I8a0037ad2845a3fbba9da380a8b8a576['h04862] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02432] =  I8a0037ad2845a3fbba9da380a8b8a576['h04864] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02433] =  I8a0037ad2845a3fbba9da380a8b8a576['h04866] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02434] =  I8a0037ad2845a3fbba9da380a8b8a576['h04868] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02435] =  I8a0037ad2845a3fbba9da380a8b8a576['h0486a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02436] =  I8a0037ad2845a3fbba9da380a8b8a576['h0486c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02437] =  I8a0037ad2845a3fbba9da380a8b8a576['h0486e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02438] =  I8a0037ad2845a3fbba9da380a8b8a576['h04870] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02439] =  I8a0037ad2845a3fbba9da380a8b8a576['h04872] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0243a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04874] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0243b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04876] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0243c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04878] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0243d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0487a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0243e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0487c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0243f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0487e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02440] =  I8a0037ad2845a3fbba9da380a8b8a576['h04880] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02441] =  I8a0037ad2845a3fbba9da380a8b8a576['h04882] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02442] =  I8a0037ad2845a3fbba9da380a8b8a576['h04884] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02443] =  I8a0037ad2845a3fbba9da380a8b8a576['h04886] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02444] =  I8a0037ad2845a3fbba9da380a8b8a576['h04888] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02445] =  I8a0037ad2845a3fbba9da380a8b8a576['h0488a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02446] =  I8a0037ad2845a3fbba9da380a8b8a576['h0488c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02447] =  I8a0037ad2845a3fbba9da380a8b8a576['h0488e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02448] =  I8a0037ad2845a3fbba9da380a8b8a576['h04890] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02449] =  I8a0037ad2845a3fbba9da380a8b8a576['h04892] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0244a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04894] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0244b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04896] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0244c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04898] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0244d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0489a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0244e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0489c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0244f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0489e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02450] =  I8a0037ad2845a3fbba9da380a8b8a576['h048a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02451] =  I8a0037ad2845a3fbba9da380a8b8a576['h048a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02452] =  I8a0037ad2845a3fbba9da380a8b8a576['h048a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02453] =  I8a0037ad2845a3fbba9da380a8b8a576['h048a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02454] =  I8a0037ad2845a3fbba9da380a8b8a576['h048a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02455] =  I8a0037ad2845a3fbba9da380a8b8a576['h048aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02456] =  I8a0037ad2845a3fbba9da380a8b8a576['h048ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02457] =  I8a0037ad2845a3fbba9da380a8b8a576['h048ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02458] =  I8a0037ad2845a3fbba9da380a8b8a576['h048b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02459] =  I8a0037ad2845a3fbba9da380a8b8a576['h048b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0245a] =  I8a0037ad2845a3fbba9da380a8b8a576['h048b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0245b] =  I8a0037ad2845a3fbba9da380a8b8a576['h048b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0245c] =  I8a0037ad2845a3fbba9da380a8b8a576['h048b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0245d] =  I8a0037ad2845a3fbba9da380a8b8a576['h048ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0245e] =  I8a0037ad2845a3fbba9da380a8b8a576['h048bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0245f] =  I8a0037ad2845a3fbba9da380a8b8a576['h048be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02460] =  I8a0037ad2845a3fbba9da380a8b8a576['h048c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02461] =  I8a0037ad2845a3fbba9da380a8b8a576['h048c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02462] =  I8a0037ad2845a3fbba9da380a8b8a576['h048c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02463] =  I8a0037ad2845a3fbba9da380a8b8a576['h048c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02464] =  I8a0037ad2845a3fbba9da380a8b8a576['h048c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02465] =  I8a0037ad2845a3fbba9da380a8b8a576['h048ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02466] =  I8a0037ad2845a3fbba9da380a8b8a576['h048cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02467] =  I8a0037ad2845a3fbba9da380a8b8a576['h048ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02468] =  I8a0037ad2845a3fbba9da380a8b8a576['h048d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02469] =  I8a0037ad2845a3fbba9da380a8b8a576['h048d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0246a] =  I8a0037ad2845a3fbba9da380a8b8a576['h048d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0246b] =  I8a0037ad2845a3fbba9da380a8b8a576['h048d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0246c] =  I8a0037ad2845a3fbba9da380a8b8a576['h048d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0246d] =  I8a0037ad2845a3fbba9da380a8b8a576['h048da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0246e] =  I8a0037ad2845a3fbba9da380a8b8a576['h048dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0246f] =  I8a0037ad2845a3fbba9da380a8b8a576['h048de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02470] =  I8a0037ad2845a3fbba9da380a8b8a576['h048e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02471] =  I8a0037ad2845a3fbba9da380a8b8a576['h048e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02472] =  I8a0037ad2845a3fbba9da380a8b8a576['h048e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02473] =  I8a0037ad2845a3fbba9da380a8b8a576['h048e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02474] =  I8a0037ad2845a3fbba9da380a8b8a576['h048e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02475] =  I8a0037ad2845a3fbba9da380a8b8a576['h048ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02476] =  I8a0037ad2845a3fbba9da380a8b8a576['h048ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02477] =  I8a0037ad2845a3fbba9da380a8b8a576['h048ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02478] =  I8a0037ad2845a3fbba9da380a8b8a576['h048f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02479] =  I8a0037ad2845a3fbba9da380a8b8a576['h048f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0247a] =  I8a0037ad2845a3fbba9da380a8b8a576['h048f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0247b] =  I8a0037ad2845a3fbba9da380a8b8a576['h048f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0247c] =  I8a0037ad2845a3fbba9da380a8b8a576['h048f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0247d] =  I8a0037ad2845a3fbba9da380a8b8a576['h048fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0247e] =  I8a0037ad2845a3fbba9da380a8b8a576['h048fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0247f] =  I8a0037ad2845a3fbba9da380a8b8a576['h048fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02480] =  I8a0037ad2845a3fbba9da380a8b8a576['h04900] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02481] =  I8a0037ad2845a3fbba9da380a8b8a576['h04902] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02482] =  I8a0037ad2845a3fbba9da380a8b8a576['h04904] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02483] =  I8a0037ad2845a3fbba9da380a8b8a576['h04906] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02484] =  I8a0037ad2845a3fbba9da380a8b8a576['h04908] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02485] =  I8a0037ad2845a3fbba9da380a8b8a576['h0490a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02486] =  I8a0037ad2845a3fbba9da380a8b8a576['h0490c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02487] =  I8a0037ad2845a3fbba9da380a8b8a576['h0490e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02488] =  I8a0037ad2845a3fbba9da380a8b8a576['h04910] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02489] =  I8a0037ad2845a3fbba9da380a8b8a576['h04912] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0248a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04914] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0248b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04916] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0248c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04918] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0248d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0491a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0248e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0491c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0248f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0491e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02490] =  I8a0037ad2845a3fbba9da380a8b8a576['h04920] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02491] =  I8a0037ad2845a3fbba9da380a8b8a576['h04922] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02492] =  I8a0037ad2845a3fbba9da380a8b8a576['h04924] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02493] =  I8a0037ad2845a3fbba9da380a8b8a576['h04926] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02494] =  I8a0037ad2845a3fbba9da380a8b8a576['h04928] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02495] =  I8a0037ad2845a3fbba9da380a8b8a576['h0492a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02496] =  I8a0037ad2845a3fbba9da380a8b8a576['h0492c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02497] =  I8a0037ad2845a3fbba9da380a8b8a576['h0492e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02498] =  I8a0037ad2845a3fbba9da380a8b8a576['h04930] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02499] =  I8a0037ad2845a3fbba9da380a8b8a576['h04932] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0249a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04934] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0249b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04936] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0249c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04938] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0249d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0493a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0249e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0493c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0249f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0493e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04940] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04942] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04944] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04946] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04948] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0494a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0494c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0494e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04950] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04952] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h04954] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h04956] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h04958] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0495a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0495c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024af] =  I8a0037ad2845a3fbba9da380a8b8a576['h0495e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04960] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04962] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04964] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04966] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04968] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0496a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0496c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0496e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04970] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04972] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h04974] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h04976] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h04978] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0497a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024be] =  I8a0037ad2845a3fbba9da380a8b8a576['h0497c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0497e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04980] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04982] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04984] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04986] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04988] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0498a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0498c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0498e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04990] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04992] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h04994] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h04996] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h04998] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0499a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0499c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0499e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h049a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h049a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h049a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h049a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h049a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h049aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h049ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h049ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h049b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h049b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024da] =  I8a0037ad2845a3fbba9da380a8b8a576['h049b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024db] =  I8a0037ad2845a3fbba9da380a8b8a576['h049b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h049b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h049ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024de] =  I8a0037ad2845a3fbba9da380a8b8a576['h049bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024df] =  I8a0037ad2845a3fbba9da380a8b8a576['h049be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h049c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h049c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h049c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h049c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h049c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h049ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h049cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h049ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h049d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h049d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h049d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h049d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h049d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h049da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h049dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h049de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h049e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h049e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h049e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h049e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h049e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h049ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h049ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h049ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h049f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h049f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h049f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h049f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h049f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h049fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h049fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h024ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h049fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02500] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02501] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02502] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02503] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02504] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02505] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02506] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02507] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02508] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02509] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0250a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0250b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0250c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0250d] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0250e] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0250f] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02510] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02511] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02512] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02513] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02514] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02515] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02516] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02517] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02518] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02519] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0251a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0251b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0251c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0251d] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0251e] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0251f] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02520] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02521] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02522] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02523] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02524] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02525] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02526] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02527] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02528] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02529] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0252a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0252b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0252c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0252d] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0252e] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0252f] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02530] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02531] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02532] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02533] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02534] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02535] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02536] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02537] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02538] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02539] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0253a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0253b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0253c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0253d] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0253e] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0253f] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02540] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02541] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02542] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02543] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02544] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02545] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02546] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02547] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02548] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02549] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0254a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0254b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0254c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0254d] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0254e] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0254f] =  I8a0037ad2845a3fbba9da380a8b8a576['h04a9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02550] =  I8a0037ad2845a3fbba9da380a8b8a576['h04aa0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02551] =  I8a0037ad2845a3fbba9da380a8b8a576['h04aa2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02552] =  I8a0037ad2845a3fbba9da380a8b8a576['h04aa4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02553] =  I8a0037ad2845a3fbba9da380a8b8a576['h04aa6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02554] =  I8a0037ad2845a3fbba9da380a8b8a576['h04aa8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02555] =  I8a0037ad2845a3fbba9da380a8b8a576['h04aaa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02556] =  I8a0037ad2845a3fbba9da380a8b8a576['h04aac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02557] =  I8a0037ad2845a3fbba9da380a8b8a576['h04aae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02558] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ab0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02559] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ab2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0255a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ab4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0255b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ab6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0255c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ab8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0255d] =  I8a0037ad2845a3fbba9da380a8b8a576['h04aba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0255e] =  I8a0037ad2845a3fbba9da380a8b8a576['h04abc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0255f] =  I8a0037ad2845a3fbba9da380a8b8a576['h04abe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02560] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ac0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02561] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ac2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02562] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ac4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02563] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ac6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02564] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ac8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02565] =  I8a0037ad2845a3fbba9da380a8b8a576['h04aca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02566] =  I8a0037ad2845a3fbba9da380a8b8a576['h04acc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02567] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ace] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02568] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ad0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02569] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ad2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0256a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ad4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0256b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ad6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0256c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ad8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0256d] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ada] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0256e] =  I8a0037ad2845a3fbba9da380a8b8a576['h04adc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0256f] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ade] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02570] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ae0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02571] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ae2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02572] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ae4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02573] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ae6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02574] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ae8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02575] =  I8a0037ad2845a3fbba9da380a8b8a576['h04aea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02576] =  I8a0037ad2845a3fbba9da380a8b8a576['h04aec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02577] =  I8a0037ad2845a3fbba9da380a8b8a576['h04aee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02578] =  I8a0037ad2845a3fbba9da380a8b8a576['h04af0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02579] =  I8a0037ad2845a3fbba9da380a8b8a576['h04af2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0257a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04af4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0257b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04af6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0257c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04af8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0257d] =  I8a0037ad2845a3fbba9da380a8b8a576['h04afa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0257e] =  I8a0037ad2845a3fbba9da380a8b8a576['h04afc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0257f] =  I8a0037ad2845a3fbba9da380a8b8a576['h04afe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02580] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02581] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02582] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02583] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02584] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02585] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02586] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02587] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02588] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02589] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0258a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0258b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0258c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0258d] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0258e] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0258f] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02590] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02591] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02592] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02593] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02594] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02595] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02596] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02597] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02598] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02599] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0259a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0259b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0259c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0259d] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0259e] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0259f] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025af] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025be] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h04b9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ba0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ba2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ba4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ba6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ba8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h04baa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025da] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025db] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025de] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025df] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bcc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bdc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04be0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04be2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04be4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04be6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04be8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bf0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bf2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bf4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bf6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bf8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bfa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bfc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h025ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h04bfe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02600] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02601] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02602] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02603] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02604] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02605] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02606] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02607] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02608] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02609] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0260a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0260b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0260c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0260d] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0260e] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0260f] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02610] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02611] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02612] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02613] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02614] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02615] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02616] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02617] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02618] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02619] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0261a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0261b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0261c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0261d] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0261e] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0261f] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02620] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02621] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02622] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02623] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02624] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02625] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02626] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02627] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02628] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02629] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0262a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0262b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0262c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0262d] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0262e] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0262f] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02630] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02631] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02632] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02633] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02634] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02635] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02636] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02637] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02638] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02639] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0263a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0263b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0263c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0263d] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0263e] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0263f] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02640] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02641] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02642] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02643] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02644] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02645] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02646] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02647] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02648] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02649] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0264a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0264b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0264c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0264d] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0264e] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0264f] =  I8a0037ad2845a3fbba9da380a8b8a576['h04c9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02650] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ca0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02651] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ca2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02652] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ca4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02653] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ca6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02654] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ca8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02655] =  I8a0037ad2845a3fbba9da380a8b8a576['h04caa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02656] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02657] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02658] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02659] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0265a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0265b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0265c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0265d] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0265e] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0265f] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02660] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02661] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02662] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02663] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02664] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02665] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02666] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ccc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02667] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02668] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02669] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0266a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0266b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0266c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0266d] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0266e] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cdc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0266f] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02670] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ce0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02671] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ce2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02672] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ce4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02673] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ce6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02674] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ce8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02675] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02676] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02677] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02678] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cf0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02679] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cf2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0267a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cf4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0267b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cf6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0267c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cf8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0267d] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cfa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0267e] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cfc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0267f] =  I8a0037ad2845a3fbba9da380a8b8a576['h04cfe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02680] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02681] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02682] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02683] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02684] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02685] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02686] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02687] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02688] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02689] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0268a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0268b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0268c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0268d] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0268e] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0268f] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02690] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02691] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02692] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02693] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02694] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02695] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02696] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02697] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02698] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02699] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0269a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0269b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0269c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0269d] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0269e] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0269f] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026af] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026be] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h04d9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04da0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04da2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04da4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04da6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04da8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h04daa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h04dac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h04dae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04db0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04db2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026da] =  I8a0037ad2845a3fbba9da380a8b8a576['h04db4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026db] =  I8a0037ad2845a3fbba9da380a8b8a576['h04db6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h04db8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h04dba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026de] =  I8a0037ad2845a3fbba9da380a8b8a576['h04dbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026df] =  I8a0037ad2845a3fbba9da380a8b8a576['h04dbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04dc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04dc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04dc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04dc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04dc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h04dca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h04dcc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h04dce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04dd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04dd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h04dd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h04dd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h04dd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h04dda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ddc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h04dde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04de0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04de2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04de4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04de6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04de8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h04dea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h04dec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h04dee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04df0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04df2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h04df4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h04df6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h04df8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h04dfa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h04dfc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h026ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h04dfe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02700] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02701] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02702] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02703] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02704] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02705] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02706] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02707] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02708] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02709] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0270a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0270b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0270c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0270d] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0270e] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0270f] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02710] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02711] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02712] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02713] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02714] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02715] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02716] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02717] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02718] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02719] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0271a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0271b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0271c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0271d] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0271e] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0271f] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02720] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02721] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02722] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02723] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02724] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02725] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02726] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02727] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02728] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02729] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0272a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0272b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0272c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0272d] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0272e] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0272f] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02730] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02731] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02732] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02733] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02734] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02735] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02736] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02737] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02738] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02739] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0273a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0273b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0273c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0273d] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0273e] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0273f] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02740] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02741] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02742] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02743] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02744] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02745] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02746] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02747] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02748] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02749] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0274a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0274b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0274c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0274d] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0274e] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0274f] =  I8a0037ad2845a3fbba9da380a8b8a576['h04e9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02750] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ea0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02751] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ea2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02752] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ea4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02753] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ea6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02754] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ea8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02755] =  I8a0037ad2845a3fbba9da380a8b8a576['h04eaa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02756] =  I8a0037ad2845a3fbba9da380a8b8a576['h04eac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02757] =  I8a0037ad2845a3fbba9da380a8b8a576['h04eae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02758] =  I8a0037ad2845a3fbba9da380a8b8a576['h04eb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02759] =  I8a0037ad2845a3fbba9da380a8b8a576['h04eb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0275a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04eb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0275b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04eb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0275c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04eb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0275d] =  I8a0037ad2845a3fbba9da380a8b8a576['h04eba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0275e] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ebc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0275f] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ebe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02760] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ec0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02761] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ec2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02762] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ec4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02763] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ec6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02764] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ec8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02765] =  I8a0037ad2845a3fbba9da380a8b8a576['h04eca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02766] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ecc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02767] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ece] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02768] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ed0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02769] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ed2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0276a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ed4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0276b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ed6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0276c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ed8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0276d] =  I8a0037ad2845a3fbba9da380a8b8a576['h04eda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0276e] =  I8a0037ad2845a3fbba9da380a8b8a576['h04edc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0276f] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ede] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02770] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ee0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02771] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ee2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02772] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ee4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02773] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ee6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02774] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ee8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02775] =  I8a0037ad2845a3fbba9da380a8b8a576['h04eea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02776] =  I8a0037ad2845a3fbba9da380a8b8a576['h04eec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02777] =  I8a0037ad2845a3fbba9da380a8b8a576['h04eee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02778] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ef0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02779] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ef2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0277a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ef4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0277b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ef6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0277c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ef8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0277d] =  I8a0037ad2845a3fbba9da380a8b8a576['h04efa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0277e] =  I8a0037ad2845a3fbba9da380a8b8a576['h04efc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0277f] =  I8a0037ad2845a3fbba9da380a8b8a576['h04efe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02780] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02781] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02782] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02783] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02784] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02785] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02786] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02787] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02788] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02789] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0278a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0278b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0278c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0278d] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0278e] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0278f] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02790] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02791] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02792] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02793] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02794] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02795] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02796] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02797] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02798] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02799] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0279a] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0279b] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0279c] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0279d] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0279e] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0279f] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027af] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027be] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h04f9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fa0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fa2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fa4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fa6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fa8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h04faa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027da] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027db] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027de] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027df] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fcc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fdc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fe0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fe2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fe4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fe6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fe8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h04fee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ff0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ff2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ff4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ff6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ff8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ffa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ffc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h027ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h04ffe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02800] =  I8a0037ad2845a3fbba9da380a8b8a576['h05000] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02801] =  I8a0037ad2845a3fbba9da380a8b8a576['h05002] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02802] =  I8a0037ad2845a3fbba9da380a8b8a576['h05004] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02803] =  I8a0037ad2845a3fbba9da380a8b8a576['h05006] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02804] =  I8a0037ad2845a3fbba9da380a8b8a576['h05008] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02805] =  I8a0037ad2845a3fbba9da380a8b8a576['h0500a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02806] =  I8a0037ad2845a3fbba9da380a8b8a576['h0500c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02807] =  I8a0037ad2845a3fbba9da380a8b8a576['h0500e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02808] =  I8a0037ad2845a3fbba9da380a8b8a576['h05010] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02809] =  I8a0037ad2845a3fbba9da380a8b8a576['h05012] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0280a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05014] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0280b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05016] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0280c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05018] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0280d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0501a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0280e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0501c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0280f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0501e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02810] =  I8a0037ad2845a3fbba9da380a8b8a576['h05020] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02811] =  I8a0037ad2845a3fbba9da380a8b8a576['h05022] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02812] =  I8a0037ad2845a3fbba9da380a8b8a576['h05024] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02813] =  I8a0037ad2845a3fbba9da380a8b8a576['h05026] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02814] =  I8a0037ad2845a3fbba9da380a8b8a576['h05028] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02815] =  I8a0037ad2845a3fbba9da380a8b8a576['h0502a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02816] =  I8a0037ad2845a3fbba9da380a8b8a576['h0502c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02817] =  I8a0037ad2845a3fbba9da380a8b8a576['h0502e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02818] =  I8a0037ad2845a3fbba9da380a8b8a576['h05030] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02819] =  I8a0037ad2845a3fbba9da380a8b8a576['h05032] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0281a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05034] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0281b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05036] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0281c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05038] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0281d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0503a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0281e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0503c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0281f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0503e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02820] =  I8a0037ad2845a3fbba9da380a8b8a576['h05040] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02821] =  I8a0037ad2845a3fbba9da380a8b8a576['h05042] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02822] =  I8a0037ad2845a3fbba9da380a8b8a576['h05044] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02823] =  I8a0037ad2845a3fbba9da380a8b8a576['h05046] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02824] =  I8a0037ad2845a3fbba9da380a8b8a576['h05048] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02825] =  I8a0037ad2845a3fbba9da380a8b8a576['h0504a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02826] =  I8a0037ad2845a3fbba9da380a8b8a576['h0504c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02827] =  I8a0037ad2845a3fbba9da380a8b8a576['h0504e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02828] =  I8a0037ad2845a3fbba9da380a8b8a576['h05050] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02829] =  I8a0037ad2845a3fbba9da380a8b8a576['h05052] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0282a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05054] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0282b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05056] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0282c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05058] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0282d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0505a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0282e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0505c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0282f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0505e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02830] =  I8a0037ad2845a3fbba9da380a8b8a576['h05060] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02831] =  I8a0037ad2845a3fbba9da380a8b8a576['h05062] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02832] =  I8a0037ad2845a3fbba9da380a8b8a576['h05064] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02833] =  I8a0037ad2845a3fbba9da380a8b8a576['h05066] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02834] =  I8a0037ad2845a3fbba9da380a8b8a576['h05068] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02835] =  I8a0037ad2845a3fbba9da380a8b8a576['h0506a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02836] =  I8a0037ad2845a3fbba9da380a8b8a576['h0506c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02837] =  I8a0037ad2845a3fbba9da380a8b8a576['h0506e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02838] =  I8a0037ad2845a3fbba9da380a8b8a576['h05070] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02839] =  I8a0037ad2845a3fbba9da380a8b8a576['h05072] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0283a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05074] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0283b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05076] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0283c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05078] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0283d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0507a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0283e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0507c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0283f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0507e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02840] =  I8a0037ad2845a3fbba9da380a8b8a576['h05080] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02841] =  I8a0037ad2845a3fbba9da380a8b8a576['h05082] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02842] =  I8a0037ad2845a3fbba9da380a8b8a576['h05084] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02843] =  I8a0037ad2845a3fbba9da380a8b8a576['h05086] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02844] =  I8a0037ad2845a3fbba9da380a8b8a576['h05088] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02845] =  I8a0037ad2845a3fbba9da380a8b8a576['h0508a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02846] =  I8a0037ad2845a3fbba9da380a8b8a576['h0508c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02847] =  I8a0037ad2845a3fbba9da380a8b8a576['h0508e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02848] =  I8a0037ad2845a3fbba9da380a8b8a576['h05090] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02849] =  I8a0037ad2845a3fbba9da380a8b8a576['h05092] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0284a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05094] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0284b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05096] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0284c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05098] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0284d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0509a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0284e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0509c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0284f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0509e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02850] =  I8a0037ad2845a3fbba9da380a8b8a576['h050a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02851] =  I8a0037ad2845a3fbba9da380a8b8a576['h050a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02852] =  I8a0037ad2845a3fbba9da380a8b8a576['h050a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02853] =  I8a0037ad2845a3fbba9da380a8b8a576['h050a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02854] =  I8a0037ad2845a3fbba9da380a8b8a576['h050a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02855] =  I8a0037ad2845a3fbba9da380a8b8a576['h050aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02856] =  I8a0037ad2845a3fbba9da380a8b8a576['h050ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02857] =  I8a0037ad2845a3fbba9da380a8b8a576['h050ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02858] =  I8a0037ad2845a3fbba9da380a8b8a576['h050b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02859] =  I8a0037ad2845a3fbba9da380a8b8a576['h050b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0285a] =  I8a0037ad2845a3fbba9da380a8b8a576['h050b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0285b] =  I8a0037ad2845a3fbba9da380a8b8a576['h050b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0285c] =  I8a0037ad2845a3fbba9da380a8b8a576['h050b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0285d] =  I8a0037ad2845a3fbba9da380a8b8a576['h050ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0285e] =  I8a0037ad2845a3fbba9da380a8b8a576['h050bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0285f] =  I8a0037ad2845a3fbba9da380a8b8a576['h050be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02860] =  I8a0037ad2845a3fbba9da380a8b8a576['h050c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02861] =  I8a0037ad2845a3fbba9da380a8b8a576['h050c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02862] =  I8a0037ad2845a3fbba9da380a8b8a576['h050c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02863] =  I8a0037ad2845a3fbba9da380a8b8a576['h050c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02864] =  I8a0037ad2845a3fbba9da380a8b8a576['h050c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02865] =  I8a0037ad2845a3fbba9da380a8b8a576['h050ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02866] =  I8a0037ad2845a3fbba9da380a8b8a576['h050cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02867] =  I8a0037ad2845a3fbba9da380a8b8a576['h050ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02868] =  I8a0037ad2845a3fbba9da380a8b8a576['h050d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02869] =  I8a0037ad2845a3fbba9da380a8b8a576['h050d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0286a] =  I8a0037ad2845a3fbba9da380a8b8a576['h050d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0286b] =  I8a0037ad2845a3fbba9da380a8b8a576['h050d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0286c] =  I8a0037ad2845a3fbba9da380a8b8a576['h050d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0286d] =  I8a0037ad2845a3fbba9da380a8b8a576['h050da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0286e] =  I8a0037ad2845a3fbba9da380a8b8a576['h050dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0286f] =  I8a0037ad2845a3fbba9da380a8b8a576['h050de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02870] =  I8a0037ad2845a3fbba9da380a8b8a576['h050e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02871] =  I8a0037ad2845a3fbba9da380a8b8a576['h050e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02872] =  I8a0037ad2845a3fbba9da380a8b8a576['h050e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02873] =  I8a0037ad2845a3fbba9da380a8b8a576['h050e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02874] =  I8a0037ad2845a3fbba9da380a8b8a576['h050e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02875] =  I8a0037ad2845a3fbba9da380a8b8a576['h050ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02876] =  I8a0037ad2845a3fbba9da380a8b8a576['h050ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02877] =  I8a0037ad2845a3fbba9da380a8b8a576['h050ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02878] =  I8a0037ad2845a3fbba9da380a8b8a576['h050f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02879] =  I8a0037ad2845a3fbba9da380a8b8a576['h050f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0287a] =  I8a0037ad2845a3fbba9da380a8b8a576['h050f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0287b] =  I8a0037ad2845a3fbba9da380a8b8a576['h050f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0287c] =  I8a0037ad2845a3fbba9da380a8b8a576['h050f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0287d] =  I8a0037ad2845a3fbba9da380a8b8a576['h050fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0287e] =  I8a0037ad2845a3fbba9da380a8b8a576['h050fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0287f] =  I8a0037ad2845a3fbba9da380a8b8a576['h050fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02880] =  I8a0037ad2845a3fbba9da380a8b8a576['h05100] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02881] =  I8a0037ad2845a3fbba9da380a8b8a576['h05102] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02882] =  I8a0037ad2845a3fbba9da380a8b8a576['h05104] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02883] =  I8a0037ad2845a3fbba9da380a8b8a576['h05106] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02884] =  I8a0037ad2845a3fbba9da380a8b8a576['h05108] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02885] =  I8a0037ad2845a3fbba9da380a8b8a576['h0510a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02886] =  I8a0037ad2845a3fbba9da380a8b8a576['h0510c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02887] =  I8a0037ad2845a3fbba9da380a8b8a576['h0510e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02888] =  I8a0037ad2845a3fbba9da380a8b8a576['h05110] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02889] =  I8a0037ad2845a3fbba9da380a8b8a576['h05112] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0288a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05114] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0288b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05116] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0288c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05118] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0288d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0511a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0288e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0511c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0288f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0511e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02890] =  I8a0037ad2845a3fbba9da380a8b8a576['h05120] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02891] =  I8a0037ad2845a3fbba9da380a8b8a576['h05122] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02892] =  I8a0037ad2845a3fbba9da380a8b8a576['h05124] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02893] =  I8a0037ad2845a3fbba9da380a8b8a576['h05126] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02894] =  I8a0037ad2845a3fbba9da380a8b8a576['h05128] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02895] =  I8a0037ad2845a3fbba9da380a8b8a576['h0512a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02896] =  I8a0037ad2845a3fbba9da380a8b8a576['h0512c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02897] =  I8a0037ad2845a3fbba9da380a8b8a576['h0512e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02898] =  I8a0037ad2845a3fbba9da380a8b8a576['h05130] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02899] =  I8a0037ad2845a3fbba9da380a8b8a576['h05132] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0289a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05134] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0289b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05136] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0289c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05138] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0289d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0513a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0289e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0513c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0289f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0513e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05140] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05142] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05144] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05146] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05148] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0514a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0514c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0514e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05150] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05152] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h05154] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h05156] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h05158] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0515a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0515c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028af] =  I8a0037ad2845a3fbba9da380a8b8a576['h0515e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05160] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05162] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05164] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05166] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05168] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0516a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0516c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0516e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05170] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05172] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h05174] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h05176] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h05178] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0517a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028be] =  I8a0037ad2845a3fbba9da380a8b8a576['h0517c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0517e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05180] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05182] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05184] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05186] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05188] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0518a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0518c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0518e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05190] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05192] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h05194] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h05196] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h05198] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0519a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0519c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0519e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h051a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h051a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h051a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h051a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h051a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h051aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h051ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h051ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h051b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h051b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028da] =  I8a0037ad2845a3fbba9da380a8b8a576['h051b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028db] =  I8a0037ad2845a3fbba9da380a8b8a576['h051b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h051b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h051ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028de] =  I8a0037ad2845a3fbba9da380a8b8a576['h051bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028df] =  I8a0037ad2845a3fbba9da380a8b8a576['h051be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h051c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h051c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h051c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h051c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h051c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h051ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h051cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h051ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h051d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h051d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h051d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h051d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h051d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h051da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h051dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h051de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h051e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h051e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h051e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h051e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h051e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h051ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h051ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h051ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h051f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h051f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h051f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h051f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h051f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h051fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h051fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h028ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h051fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02900] =  I8a0037ad2845a3fbba9da380a8b8a576['h05200] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02901] =  I8a0037ad2845a3fbba9da380a8b8a576['h05202] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02902] =  I8a0037ad2845a3fbba9da380a8b8a576['h05204] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02903] =  I8a0037ad2845a3fbba9da380a8b8a576['h05206] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02904] =  I8a0037ad2845a3fbba9da380a8b8a576['h05208] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02905] =  I8a0037ad2845a3fbba9da380a8b8a576['h0520a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02906] =  I8a0037ad2845a3fbba9da380a8b8a576['h0520c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02907] =  I8a0037ad2845a3fbba9da380a8b8a576['h0520e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02908] =  I8a0037ad2845a3fbba9da380a8b8a576['h05210] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02909] =  I8a0037ad2845a3fbba9da380a8b8a576['h05212] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0290a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05214] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0290b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05216] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0290c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05218] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0290d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0521a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0290e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0521c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0290f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0521e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02910] =  I8a0037ad2845a3fbba9da380a8b8a576['h05220] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02911] =  I8a0037ad2845a3fbba9da380a8b8a576['h05222] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02912] =  I8a0037ad2845a3fbba9da380a8b8a576['h05224] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02913] =  I8a0037ad2845a3fbba9da380a8b8a576['h05226] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02914] =  I8a0037ad2845a3fbba9da380a8b8a576['h05228] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02915] =  I8a0037ad2845a3fbba9da380a8b8a576['h0522a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02916] =  I8a0037ad2845a3fbba9da380a8b8a576['h0522c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02917] =  I8a0037ad2845a3fbba9da380a8b8a576['h0522e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02918] =  I8a0037ad2845a3fbba9da380a8b8a576['h05230] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02919] =  I8a0037ad2845a3fbba9da380a8b8a576['h05232] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0291a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05234] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0291b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05236] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0291c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05238] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0291d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0523a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0291e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0523c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0291f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0523e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02920] =  I8a0037ad2845a3fbba9da380a8b8a576['h05240] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02921] =  I8a0037ad2845a3fbba9da380a8b8a576['h05242] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02922] =  I8a0037ad2845a3fbba9da380a8b8a576['h05244] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02923] =  I8a0037ad2845a3fbba9da380a8b8a576['h05246] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02924] =  I8a0037ad2845a3fbba9da380a8b8a576['h05248] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02925] =  I8a0037ad2845a3fbba9da380a8b8a576['h0524a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02926] =  I8a0037ad2845a3fbba9da380a8b8a576['h0524c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02927] =  I8a0037ad2845a3fbba9da380a8b8a576['h0524e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02928] =  I8a0037ad2845a3fbba9da380a8b8a576['h05250] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02929] =  I8a0037ad2845a3fbba9da380a8b8a576['h05252] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0292a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05254] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0292b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05256] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0292c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05258] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0292d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0525a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0292e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0525c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0292f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0525e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02930] =  I8a0037ad2845a3fbba9da380a8b8a576['h05260] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02931] =  I8a0037ad2845a3fbba9da380a8b8a576['h05262] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02932] =  I8a0037ad2845a3fbba9da380a8b8a576['h05264] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02933] =  I8a0037ad2845a3fbba9da380a8b8a576['h05266] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02934] =  I8a0037ad2845a3fbba9da380a8b8a576['h05268] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02935] =  I8a0037ad2845a3fbba9da380a8b8a576['h0526a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02936] =  I8a0037ad2845a3fbba9da380a8b8a576['h0526c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02937] =  I8a0037ad2845a3fbba9da380a8b8a576['h0526e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02938] =  I8a0037ad2845a3fbba9da380a8b8a576['h05270] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02939] =  I8a0037ad2845a3fbba9da380a8b8a576['h05272] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0293a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05274] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0293b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05276] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0293c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05278] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0293d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0527a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0293e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0527c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0293f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0527e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02940] =  I8a0037ad2845a3fbba9da380a8b8a576['h05280] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02941] =  I8a0037ad2845a3fbba9da380a8b8a576['h05282] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02942] =  I8a0037ad2845a3fbba9da380a8b8a576['h05284] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02943] =  I8a0037ad2845a3fbba9da380a8b8a576['h05286] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02944] =  I8a0037ad2845a3fbba9da380a8b8a576['h05288] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02945] =  I8a0037ad2845a3fbba9da380a8b8a576['h0528a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02946] =  I8a0037ad2845a3fbba9da380a8b8a576['h0528c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02947] =  I8a0037ad2845a3fbba9da380a8b8a576['h0528e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02948] =  I8a0037ad2845a3fbba9da380a8b8a576['h05290] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02949] =  I8a0037ad2845a3fbba9da380a8b8a576['h05292] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0294a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05294] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0294b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05296] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0294c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05298] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0294d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0529a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0294e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0529c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0294f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0529e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02950] =  I8a0037ad2845a3fbba9da380a8b8a576['h052a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02951] =  I8a0037ad2845a3fbba9da380a8b8a576['h052a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02952] =  I8a0037ad2845a3fbba9da380a8b8a576['h052a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02953] =  I8a0037ad2845a3fbba9da380a8b8a576['h052a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02954] =  I8a0037ad2845a3fbba9da380a8b8a576['h052a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02955] =  I8a0037ad2845a3fbba9da380a8b8a576['h052aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02956] =  I8a0037ad2845a3fbba9da380a8b8a576['h052ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02957] =  I8a0037ad2845a3fbba9da380a8b8a576['h052ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02958] =  I8a0037ad2845a3fbba9da380a8b8a576['h052b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02959] =  I8a0037ad2845a3fbba9da380a8b8a576['h052b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0295a] =  I8a0037ad2845a3fbba9da380a8b8a576['h052b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0295b] =  I8a0037ad2845a3fbba9da380a8b8a576['h052b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0295c] =  I8a0037ad2845a3fbba9da380a8b8a576['h052b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0295d] =  I8a0037ad2845a3fbba9da380a8b8a576['h052ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0295e] =  I8a0037ad2845a3fbba9da380a8b8a576['h052bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0295f] =  I8a0037ad2845a3fbba9da380a8b8a576['h052be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02960] =  I8a0037ad2845a3fbba9da380a8b8a576['h052c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02961] =  I8a0037ad2845a3fbba9da380a8b8a576['h052c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02962] =  I8a0037ad2845a3fbba9da380a8b8a576['h052c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02963] =  I8a0037ad2845a3fbba9da380a8b8a576['h052c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02964] =  I8a0037ad2845a3fbba9da380a8b8a576['h052c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02965] =  I8a0037ad2845a3fbba9da380a8b8a576['h052ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02966] =  I8a0037ad2845a3fbba9da380a8b8a576['h052cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02967] =  I8a0037ad2845a3fbba9da380a8b8a576['h052ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02968] =  I8a0037ad2845a3fbba9da380a8b8a576['h052d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02969] =  I8a0037ad2845a3fbba9da380a8b8a576['h052d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0296a] =  I8a0037ad2845a3fbba9da380a8b8a576['h052d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0296b] =  I8a0037ad2845a3fbba9da380a8b8a576['h052d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0296c] =  I8a0037ad2845a3fbba9da380a8b8a576['h052d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0296d] =  I8a0037ad2845a3fbba9da380a8b8a576['h052da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0296e] =  I8a0037ad2845a3fbba9da380a8b8a576['h052dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0296f] =  I8a0037ad2845a3fbba9da380a8b8a576['h052de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02970] =  I8a0037ad2845a3fbba9da380a8b8a576['h052e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02971] =  I8a0037ad2845a3fbba9da380a8b8a576['h052e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02972] =  I8a0037ad2845a3fbba9da380a8b8a576['h052e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02973] =  I8a0037ad2845a3fbba9da380a8b8a576['h052e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02974] =  I8a0037ad2845a3fbba9da380a8b8a576['h052e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02975] =  I8a0037ad2845a3fbba9da380a8b8a576['h052ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02976] =  I8a0037ad2845a3fbba9da380a8b8a576['h052ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02977] =  I8a0037ad2845a3fbba9da380a8b8a576['h052ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02978] =  I8a0037ad2845a3fbba9da380a8b8a576['h052f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02979] =  I8a0037ad2845a3fbba9da380a8b8a576['h052f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0297a] =  I8a0037ad2845a3fbba9da380a8b8a576['h052f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0297b] =  I8a0037ad2845a3fbba9da380a8b8a576['h052f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0297c] =  I8a0037ad2845a3fbba9da380a8b8a576['h052f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0297d] =  I8a0037ad2845a3fbba9da380a8b8a576['h052fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0297e] =  I8a0037ad2845a3fbba9da380a8b8a576['h052fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0297f] =  I8a0037ad2845a3fbba9da380a8b8a576['h052fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02980] =  I8a0037ad2845a3fbba9da380a8b8a576['h05300] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02981] =  I8a0037ad2845a3fbba9da380a8b8a576['h05302] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02982] =  I8a0037ad2845a3fbba9da380a8b8a576['h05304] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02983] =  I8a0037ad2845a3fbba9da380a8b8a576['h05306] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02984] =  I8a0037ad2845a3fbba9da380a8b8a576['h05308] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02985] =  I8a0037ad2845a3fbba9da380a8b8a576['h0530a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02986] =  I8a0037ad2845a3fbba9da380a8b8a576['h0530c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02987] =  I8a0037ad2845a3fbba9da380a8b8a576['h0530e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02988] =  I8a0037ad2845a3fbba9da380a8b8a576['h05310] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02989] =  I8a0037ad2845a3fbba9da380a8b8a576['h05312] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0298a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05314] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0298b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05316] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0298c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05318] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0298d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0531a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0298e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0531c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0298f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0531e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02990] =  I8a0037ad2845a3fbba9da380a8b8a576['h05320] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02991] =  I8a0037ad2845a3fbba9da380a8b8a576['h05322] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02992] =  I8a0037ad2845a3fbba9da380a8b8a576['h05324] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02993] =  I8a0037ad2845a3fbba9da380a8b8a576['h05326] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02994] =  I8a0037ad2845a3fbba9da380a8b8a576['h05328] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02995] =  I8a0037ad2845a3fbba9da380a8b8a576['h0532a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02996] =  I8a0037ad2845a3fbba9da380a8b8a576['h0532c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02997] =  I8a0037ad2845a3fbba9da380a8b8a576['h0532e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02998] =  I8a0037ad2845a3fbba9da380a8b8a576['h05330] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02999] =  I8a0037ad2845a3fbba9da380a8b8a576['h05332] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0299a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05334] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0299b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05336] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0299c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05338] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0299d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0533a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0299e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0533c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0299f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0533e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05340] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05342] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05344] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05346] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05348] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0534a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0534c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0534e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05350] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05352] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h05354] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h05356] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h05358] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0535a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0535c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029af] =  I8a0037ad2845a3fbba9da380a8b8a576['h0535e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05360] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05362] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05364] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05366] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05368] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0536a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0536c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0536e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05370] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05372] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h05374] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h05376] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h05378] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0537a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029be] =  I8a0037ad2845a3fbba9da380a8b8a576['h0537c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0537e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05380] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05382] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05384] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05386] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05388] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0538a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0538c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0538e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05390] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05392] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h05394] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h05396] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h05398] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0539a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0539c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0539e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h053a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h053a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h053a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h053a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h053a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h053aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h053ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h053ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h053b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h053b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029da] =  I8a0037ad2845a3fbba9da380a8b8a576['h053b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029db] =  I8a0037ad2845a3fbba9da380a8b8a576['h053b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h053b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h053ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029de] =  I8a0037ad2845a3fbba9da380a8b8a576['h053bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029df] =  I8a0037ad2845a3fbba9da380a8b8a576['h053be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h053c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h053c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h053c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h053c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h053c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h053ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h053cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h053ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h053d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h053d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h053d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h053d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h053d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h053da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h053dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h053de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h053e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h053e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h053e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h053e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h053e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h053ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h053ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h053ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h053f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h053f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h053f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h053f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h053f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h053fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h053fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h029ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h053fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a00] =  I8a0037ad2845a3fbba9da380a8b8a576['h05400] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a01] =  I8a0037ad2845a3fbba9da380a8b8a576['h05402] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a02] =  I8a0037ad2845a3fbba9da380a8b8a576['h05404] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a03] =  I8a0037ad2845a3fbba9da380a8b8a576['h05406] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a04] =  I8a0037ad2845a3fbba9da380a8b8a576['h05408] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a05] =  I8a0037ad2845a3fbba9da380a8b8a576['h0540a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a06] =  I8a0037ad2845a3fbba9da380a8b8a576['h0540c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a07] =  I8a0037ad2845a3fbba9da380a8b8a576['h0540e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a08] =  I8a0037ad2845a3fbba9da380a8b8a576['h05410] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a09] =  I8a0037ad2845a3fbba9da380a8b8a576['h05412] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a0a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05414] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a0b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05416] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a0c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05418] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a0d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0541a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a0e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0541c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a0f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0541e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a10] =  I8a0037ad2845a3fbba9da380a8b8a576['h05420] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a11] =  I8a0037ad2845a3fbba9da380a8b8a576['h05422] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a12] =  I8a0037ad2845a3fbba9da380a8b8a576['h05424] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a13] =  I8a0037ad2845a3fbba9da380a8b8a576['h05426] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a14] =  I8a0037ad2845a3fbba9da380a8b8a576['h05428] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a15] =  I8a0037ad2845a3fbba9da380a8b8a576['h0542a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a16] =  I8a0037ad2845a3fbba9da380a8b8a576['h0542c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a17] =  I8a0037ad2845a3fbba9da380a8b8a576['h0542e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a18] =  I8a0037ad2845a3fbba9da380a8b8a576['h05430] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a19] =  I8a0037ad2845a3fbba9da380a8b8a576['h05432] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a1a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05434] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a1b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05436] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a1c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05438] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a1d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0543a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a1e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0543c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a1f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0543e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a20] =  I8a0037ad2845a3fbba9da380a8b8a576['h05440] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a21] =  I8a0037ad2845a3fbba9da380a8b8a576['h05442] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a22] =  I8a0037ad2845a3fbba9da380a8b8a576['h05444] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a23] =  I8a0037ad2845a3fbba9da380a8b8a576['h05446] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a24] =  I8a0037ad2845a3fbba9da380a8b8a576['h05448] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a25] =  I8a0037ad2845a3fbba9da380a8b8a576['h0544a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a26] =  I8a0037ad2845a3fbba9da380a8b8a576['h0544c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a27] =  I8a0037ad2845a3fbba9da380a8b8a576['h0544e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a28] =  I8a0037ad2845a3fbba9da380a8b8a576['h05450] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a29] =  I8a0037ad2845a3fbba9da380a8b8a576['h05452] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a2a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05454] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a2b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05456] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a2c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05458] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a2d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0545a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a2e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0545c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a2f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0545e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a30] =  I8a0037ad2845a3fbba9da380a8b8a576['h05460] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a31] =  I8a0037ad2845a3fbba9da380a8b8a576['h05462] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a32] =  I8a0037ad2845a3fbba9da380a8b8a576['h05464] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a33] =  I8a0037ad2845a3fbba9da380a8b8a576['h05466] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a34] =  I8a0037ad2845a3fbba9da380a8b8a576['h05468] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a35] =  I8a0037ad2845a3fbba9da380a8b8a576['h0546a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a36] =  I8a0037ad2845a3fbba9da380a8b8a576['h0546c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a37] =  I8a0037ad2845a3fbba9da380a8b8a576['h0546e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a38] =  I8a0037ad2845a3fbba9da380a8b8a576['h05470] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a39] =  I8a0037ad2845a3fbba9da380a8b8a576['h05472] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a3a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05474] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a3b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05476] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a3c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05478] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a3d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0547a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a3e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0547c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a3f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0547e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a40] =  I8a0037ad2845a3fbba9da380a8b8a576['h05480] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a41] =  I8a0037ad2845a3fbba9da380a8b8a576['h05482] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a42] =  I8a0037ad2845a3fbba9da380a8b8a576['h05484] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a43] =  I8a0037ad2845a3fbba9da380a8b8a576['h05486] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a44] =  I8a0037ad2845a3fbba9da380a8b8a576['h05488] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a45] =  I8a0037ad2845a3fbba9da380a8b8a576['h0548a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a46] =  I8a0037ad2845a3fbba9da380a8b8a576['h0548c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a47] =  I8a0037ad2845a3fbba9da380a8b8a576['h0548e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a48] =  I8a0037ad2845a3fbba9da380a8b8a576['h05490] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a49] =  I8a0037ad2845a3fbba9da380a8b8a576['h05492] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a4a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05494] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a4b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05496] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a4c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05498] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a4d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0549a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a4e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0549c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a4f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0549e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a50] =  I8a0037ad2845a3fbba9da380a8b8a576['h054a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a51] =  I8a0037ad2845a3fbba9da380a8b8a576['h054a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a52] =  I8a0037ad2845a3fbba9da380a8b8a576['h054a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a53] =  I8a0037ad2845a3fbba9da380a8b8a576['h054a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a54] =  I8a0037ad2845a3fbba9da380a8b8a576['h054a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a55] =  I8a0037ad2845a3fbba9da380a8b8a576['h054aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a56] =  I8a0037ad2845a3fbba9da380a8b8a576['h054ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a57] =  I8a0037ad2845a3fbba9da380a8b8a576['h054ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a58] =  I8a0037ad2845a3fbba9da380a8b8a576['h054b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a59] =  I8a0037ad2845a3fbba9da380a8b8a576['h054b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a5a] =  I8a0037ad2845a3fbba9da380a8b8a576['h054b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a5b] =  I8a0037ad2845a3fbba9da380a8b8a576['h054b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a5c] =  I8a0037ad2845a3fbba9da380a8b8a576['h054b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a5d] =  I8a0037ad2845a3fbba9da380a8b8a576['h054ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a5e] =  I8a0037ad2845a3fbba9da380a8b8a576['h054bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a5f] =  I8a0037ad2845a3fbba9da380a8b8a576['h054be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a60] =  I8a0037ad2845a3fbba9da380a8b8a576['h054c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a61] =  I8a0037ad2845a3fbba9da380a8b8a576['h054c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a62] =  I8a0037ad2845a3fbba9da380a8b8a576['h054c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a63] =  I8a0037ad2845a3fbba9da380a8b8a576['h054c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a64] =  I8a0037ad2845a3fbba9da380a8b8a576['h054c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a65] =  I8a0037ad2845a3fbba9da380a8b8a576['h054ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a66] =  I8a0037ad2845a3fbba9da380a8b8a576['h054cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a67] =  I8a0037ad2845a3fbba9da380a8b8a576['h054ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a68] =  I8a0037ad2845a3fbba9da380a8b8a576['h054d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a69] =  I8a0037ad2845a3fbba9da380a8b8a576['h054d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a6a] =  I8a0037ad2845a3fbba9da380a8b8a576['h054d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a6b] =  I8a0037ad2845a3fbba9da380a8b8a576['h054d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a6c] =  I8a0037ad2845a3fbba9da380a8b8a576['h054d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a6d] =  I8a0037ad2845a3fbba9da380a8b8a576['h054da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a6e] =  I8a0037ad2845a3fbba9da380a8b8a576['h054dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a6f] =  I8a0037ad2845a3fbba9da380a8b8a576['h054de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a70] =  I8a0037ad2845a3fbba9da380a8b8a576['h054e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a71] =  I8a0037ad2845a3fbba9da380a8b8a576['h054e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a72] =  I8a0037ad2845a3fbba9da380a8b8a576['h054e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a73] =  I8a0037ad2845a3fbba9da380a8b8a576['h054e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a74] =  I8a0037ad2845a3fbba9da380a8b8a576['h054e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a75] =  I8a0037ad2845a3fbba9da380a8b8a576['h054ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a76] =  I8a0037ad2845a3fbba9da380a8b8a576['h054ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a77] =  I8a0037ad2845a3fbba9da380a8b8a576['h054ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a78] =  I8a0037ad2845a3fbba9da380a8b8a576['h054f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a79] =  I8a0037ad2845a3fbba9da380a8b8a576['h054f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a7a] =  I8a0037ad2845a3fbba9da380a8b8a576['h054f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a7b] =  I8a0037ad2845a3fbba9da380a8b8a576['h054f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a7c] =  I8a0037ad2845a3fbba9da380a8b8a576['h054f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a7d] =  I8a0037ad2845a3fbba9da380a8b8a576['h054fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a7e] =  I8a0037ad2845a3fbba9da380a8b8a576['h054fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a7f] =  I8a0037ad2845a3fbba9da380a8b8a576['h054fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a80] =  I8a0037ad2845a3fbba9da380a8b8a576['h05500] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a81] =  I8a0037ad2845a3fbba9da380a8b8a576['h05502] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a82] =  I8a0037ad2845a3fbba9da380a8b8a576['h05504] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a83] =  I8a0037ad2845a3fbba9da380a8b8a576['h05506] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a84] =  I8a0037ad2845a3fbba9da380a8b8a576['h05508] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a85] =  I8a0037ad2845a3fbba9da380a8b8a576['h0550a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a86] =  I8a0037ad2845a3fbba9da380a8b8a576['h0550c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a87] =  I8a0037ad2845a3fbba9da380a8b8a576['h0550e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a88] =  I8a0037ad2845a3fbba9da380a8b8a576['h05510] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a89] =  I8a0037ad2845a3fbba9da380a8b8a576['h05512] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a8a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05514] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a8b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05516] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a8c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05518] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a8d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0551a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a8e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0551c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a8f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0551e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a90] =  I8a0037ad2845a3fbba9da380a8b8a576['h05520] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a91] =  I8a0037ad2845a3fbba9da380a8b8a576['h05522] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a92] =  I8a0037ad2845a3fbba9da380a8b8a576['h05524] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a93] =  I8a0037ad2845a3fbba9da380a8b8a576['h05526] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a94] =  I8a0037ad2845a3fbba9da380a8b8a576['h05528] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a95] =  I8a0037ad2845a3fbba9da380a8b8a576['h0552a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a96] =  I8a0037ad2845a3fbba9da380a8b8a576['h0552c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a97] =  I8a0037ad2845a3fbba9da380a8b8a576['h0552e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a98] =  I8a0037ad2845a3fbba9da380a8b8a576['h05530] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a99] =  I8a0037ad2845a3fbba9da380a8b8a576['h05532] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a9a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05534] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a9b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05536] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a9c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05538] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a9d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0553a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a9e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0553c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02a9f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0553e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02aa0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05540] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02aa1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05542] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02aa2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05544] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02aa3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05546] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02aa4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05548] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02aa5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0554a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02aa6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0554c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02aa7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0554e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02aa8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05550] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02aa9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05552] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02aaa] =  I8a0037ad2845a3fbba9da380a8b8a576['h05554] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02aab] =  I8a0037ad2845a3fbba9da380a8b8a576['h05556] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02aac] =  I8a0037ad2845a3fbba9da380a8b8a576['h05558] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02aad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0555a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02aae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0555c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02aaf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0555e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ab0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05560] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ab1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05562] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ab2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05564] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ab3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05566] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ab4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05568] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ab5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0556a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ab6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0556c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ab7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0556e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ab8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05570] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ab9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05572] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02aba] =  I8a0037ad2845a3fbba9da380a8b8a576['h05574] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02abb] =  I8a0037ad2845a3fbba9da380a8b8a576['h05576] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02abc] =  I8a0037ad2845a3fbba9da380a8b8a576['h05578] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02abd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0557a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02abe] =  I8a0037ad2845a3fbba9da380a8b8a576['h0557c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02abf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0557e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ac0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05580] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ac1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05582] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ac2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05584] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ac3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05586] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ac4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05588] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ac5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0558a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ac6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0558c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ac7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0558e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ac8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05590] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ac9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05592] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02aca] =  I8a0037ad2845a3fbba9da380a8b8a576['h05594] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02acb] =  I8a0037ad2845a3fbba9da380a8b8a576['h05596] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02acc] =  I8a0037ad2845a3fbba9da380a8b8a576['h05598] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02acd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0559a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ace] =  I8a0037ad2845a3fbba9da380a8b8a576['h0559c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02acf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0559e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ad0] =  I8a0037ad2845a3fbba9da380a8b8a576['h055a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ad1] =  I8a0037ad2845a3fbba9da380a8b8a576['h055a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ad2] =  I8a0037ad2845a3fbba9da380a8b8a576['h055a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ad3] =  I8a0037ad2845a3fbba9da380a8b8a576['h055a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ad4] =  I8a0037ad2845a3fbba9da380a8b8a576['h055a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ad5] =  I8a0037ad2845a3fbba9da380a8b8a576['h055aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ad6] =  I8a0037ad2845a3fbba9da380a8b8a576['h055ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ad7] =  I8a0037ad2845a3fbba9da380a8b8a576['h055ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ad8] =  I8a0037ad2845a3fbba9da380a8b8a576['h055b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ad9] =  I8a0037ad2845a3fbba9da380a8b8a576['h055b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ada] =  I8a0037ad2845a3fbba9da380a8b8a576['h055b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02adb] =  I8a0037ad2845a3fbba9da380a8b8a576['h055b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02adc] =  I8a0037ad2845a3fbba9da380a8b8a576['h055b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02add] =  I8a0037ad2845a3fbba9da380a8b8a576['h055ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ade] =  I8a0037ad2845a3fbba9da380a8b8a576['h055bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02adf] =  I8a0037ad2845a3fbba9da380a8b8a576['h055be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ae0] =  I8a0037ad2845a3fbba9da380a8b8a576['h055c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ae1] =  I8a0037ad2845a3fbba9da380a8b8a576['h055c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ae2] =  I8a0037ad2845a3fbba9da380a8b8a576['h055c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ae3] =  I8a0037ad2845a3fbba9da380a8b8a576['h055c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ae4] =  I8a0037ad2845a3fbba9da380a8b8a576['h055c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ae5] =  I8a0037ad2845a3fbba9da380a8b8a576['h055ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ae6] =  I8a0037ad2845a3fbba9da380a8b8a576['h055cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ae7] =  I8a0037ad2845a3fbba9da380a8b8a576['h055ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ae8] =  I8a0037ad2845a3fbba9da380a8b8a576['h055d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ae9] =  I8a0037ad2845a3fbba9da380a8b8a576['h055d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02aea] =  I8a0037ad2845a3fbba9da380a8b8a576['h055d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02aeb] =  I8a0037ad2845a3fbba9da380a8b8a576['h055d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02aec] =  I8a0037ad2845a3fbba9da380a8b8a576['h055d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02aed] =  I8a0037ad2845a3fbba9da380a8b8a576['h055da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02aee] =  I8a0037ad2845a3fbba9da380a8b8a576['h055dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02aef] =  I8a0037ad2845a3fbba9da380a8b8a576['h055de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02af0] =  I8a0037ad2845a3fbba9da380a8b8a576['h055e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02af1] =  I8a0037ad2845a3fbba9da380a8b8a576['h055e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02af2] =  I8a0037ad2845a3fbba9da380a8b8a576['h055e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02af3] =  I8a0037ad2845a3fbba9da380a8b8a576['h055e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02af4] =  I8a0037ad2845a3fbba9da380a8b8a576['h055e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02af5] =  I8a0037ad2845a3fbba9da380a8b8a576['h055ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02af6] =  I8a0037ad2845a3fbba9da380a8b8a576['h055ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02af7] =  I8a0037ad2845a3fbba9da380a8b8a576['h055ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02af8] =  I8a0037ad2845a3fbba9da380a8b8a576['h055f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02af9] =  I8a0037ad2845a3fbba9da380a8b8a576['h055f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02afa] =  I8a0037ad2845a3fbba9da380a8b8a576['h055f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02afb] =  I8a0037ad2845a3fbba9da380a8b8a576['h055f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02afc] =  I8a0037ad2845a3fbba9da380a8b8a576['h055f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02afd] =  I8a0037ad2845a3fbba9da380a8b8a576['h055fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02afe] =  I8a0037ad2845a3fbba9da380a8b8a576['h055fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02aff] =  I8a0037ad2845a3fbba9da380a8b8a576['h055fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b00] =  I8a0037ad2845a3fbba9da380a8b8a576['h05600] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b01] =  I8a0037ad2845a3fbba9da380a8b8a576['h05602] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b02] =  I8a0037ad2845a3fbba9da380a8b8a576['h05604] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b03] =  I8a0037ad2845a3fbba9da380a8b8a576['h05606] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b04] =  I8a0037ad2845a3fbba9da380a8b8a576['h05608] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b05] =  I8a0037ad2845a3fbba9da380a8b8a576['h0560a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b06] =  I8a0037ad2845a3fbba9da380a8b8a576['h0560c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b07] =  I8a0037ad2845a3fbba9da380a8b8a576['h0560e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b08] =  I8a0037ad2845a3fbba9da380a8b8a576['h05610] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b09] =  I8a0037ad2845a3fbba9da380a8b8a576['h05612] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b0a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05614] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b0b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05616] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b0c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05618] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b0d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0561a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b0e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0561c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b0f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0561e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b10] =  I8a0037ad2845a3fbba9da380a8b8a576['h05620] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b11] =  I8a0037ad2845a3fbba9da380a8b8a576['h05622] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b12] =  I8a0037ad2845a3fbba9da380a8b8a576['h05624] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b13] =  I8a0037ad2845a3fbba9da380a8b8a576['h05626] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b14] =  I8a0037ad2845a3fbba9da380a8b8a576['h05628] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b15] =  I8a0037ad2845a3fbba9da380a8b8a576['h0562a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b16] =  I8a0037ad2845a3fbba9da380a8b8a576['h0562c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b17] =  I8a0037ad2845a3fbba9da380a8b8a576['h0562e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b18] =  I8a0037ad2845a3fbba9da380a8b8a576['h05630] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b19] =  I8a0037ad2845a3fbba9da380a8b8a576['h05632] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b1a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05634] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b1b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05636] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b1c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05638] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b1d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0563a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b1e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0563c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b1f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0563e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b20] =  I8a0037ad2845a3fbba9da380a8b8a576['h05640] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b21] =  I8a0037ad2845a3fbba9da380a8b8a576['h05642] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b22] =  I8a0037ad2845a3fbba9da380a8b8a576['h05644] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b23] =  I8a0037ad2845a3fbba9da380a8b8a576['h05646] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b24] =  I8a0037ad2845a3fbba9da380a8b8a576['h05648] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b25] =  I8a0037ad2845a3fbba9da380a8b8a576['h0564a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b26] =  I8a0037ad2845a3fbba9da380a8b8a576['h0564c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b27] =  I8a0037ad2845a3fbba9da380a8b8a576['h0564e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b28] =  I8a0037ad2845a3fbba9da380a8b8a576['h05650] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b29] =  I8a0037ad2845a3fbba9da380a8b8a576['h05652] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b2a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05654] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b2b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05656] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b2c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05658] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b2d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0565a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b2e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0565c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b2f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0565e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b30] =  I8a0037ad2845a3fbba9da380a8b8a576['h05660] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b31] =  I8a0037ad2845a3fbba9da380a8b8a576['h05662] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b32] =  I8a0037ad2845a3fbba9da380a8b8a576['h05664] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b33] =  I8a0037ad2845a3fbba9da380a8b8a576['h05666] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b34] =  I8a0037ad2845a3fbba9da380a8b8a576['h05668] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b35] =  I8a0037ad2845a3fbba9da380a8b8a576['h0566a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b36] =  I8a0037ad2845a3fbba9da380a8b8a576['h0566c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b37] =  I8a0037ad2845a3fbba9da380a8b8a576['h0566e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b38] =  I8a0037ad2845a3fbba9da380a8b8a576['h05670] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b39] =  I8a0037ad2845a3fbba9da380a8b8a576['h05672] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b3a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05674] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b3b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05676] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b3c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05678] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b3d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0567a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b3e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0567c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b3f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0567e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b40] =  I8a0037ad2845a3fbba9da380a8b8a576['h05680] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b41] =  I8a0037ad2845a3fbba9da380a8b8a576['h05682] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b42] =  I8a0037ad2845a3fbba9da380a8b8a576['h05684] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b43] =  I8a0037ad2845a3fbba9da380a8b8a576['h05686] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b44] =  I8a0037ad2845a3fbba9da380a8b8a576['h05688] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b45] =  I8a0037ad2845a3fbba9da380a8b8a576['h0568a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b46] =  I8a0037ad2845a3fbba9da380a8b8a576['h0568c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b47] =  I8a0037ad2845a3fbba9da380a8b8a576['h0568e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b48] =  I8a0037ad2845a3fbba9da380a8b8a576['h05690] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b49] =  I8a0037ad2845a3fbba9da380a8b8a576['h05692] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b4a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05694] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b4b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05696] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b4c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05698] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b4d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0569a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b4e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0569c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b4f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0569e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b50] =  I8a0037ad2845a3fbba9da380a8b8a576['h056a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b51] =  I8a0037ad2845a3fbba9da380a8b8a576['h056a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b52] =  I8a0037ad2845a3fbba9da380a8b8a576['h056a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b53] =  I8a0037ad2845a3fbba9da380a8b8a576['h056a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b54] =  I8a0037ad2845a3fbba9da380a8b8a576['h056a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b55] =  I8a0037ad2845a3fbba9da380a8b8a576['h056aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b56] =  I8a0037ad2845a3fbba9da380a8b8a576['h056ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b57] =  I8a0037ad2845a3fbba9da380a8b8a576['h056ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b58] =  I8a0037ad2845a3fbba9da380a8b8a576['h056b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b59] =  I8a0037ad2845a3fbba9da380a8b8a576['h056b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b5a] =  I8a0037ad2845a3fbba9da380a8b8a576['h056b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b5b] =  I8a0037ad2845a3fbba9da380a8b8a576['h056b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b5c] =  I8a0037ad2845a3fbba9da380a8b8a576['h056b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b5d] =  I8a0037ad2845a3fbba9da380a8b8a576['h056ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b5e] =  I8a0037ad2845a3fbba9da380a8b8a576['h056bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b5f] =  I8a0037ad2845a3fbba9da380a8b8a576['h056be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b60] =  I8a0037ad2845a3fbba9da380a8b8a576['h056c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b61] =  I8a0037ad2845a3fbba9da380a8b8a576['h056c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b62] =  I8a0037ad2845a3fbba9da380a8b8a576['h056c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b63] =  I8a0037ad2845a3fbba9da380a8b8a576['h056c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b64] =  I8a0037ad2845a3fbba9da380a8b8a576['h056c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b65] =  I8a0037ad2845a3fbba9da380a8b8a576['h056ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b66] =  I8a0037ad2845a3fbba9da380a8b8a576['h056cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b67] =  I8a0037ad2845a3fbba9da380a8b8a576['h056ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b68] =  I8a0037ad2845a3fbba9da380a8b8a576['h056d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b69] =  I8a0037ad2845a3fbba9da380a8b8a576['h056d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b6a] =  I8a0037ad2845a3fbba9da380a8b8a576['h056d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b6b] =  I8a0037ad2845a3fbba9da380a8b8a576['h056d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b6c] =  I8a0037ad2845a3fbba9da380a8b8a576['h056d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b6d] =  I8a0037ad2845a3fbba9da380a8b8a576['h056da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b6e] =  I8a0037ad2845a3fbba9da380a8b8a576['h056dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b6f] =  I8a0037ad2845a3fbba9da380a8b8a576['h056de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b70] =  I8a0037ad2845a3fbba9da380a8b8a576['h056e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b71] =  I8a0037ad2845a3fbba9da380a8b8a576['h056e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b72] =  I8a0037ad2845a3fbba9da380a8b8a576['h056e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b73] =  I8a0037ad2845a3fbba9da380a8b8a576['h056e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b74] =  I8a0037ad2845a3fbba9da380a8b8a576['h056e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b75] =  I8a0037ad2845a3fbba9da380a8b8a576['h056ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b76] =  I8a0037ad2845a3fbba9da380a8b8a576['h056ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b77] =  I8a0037ad2845a3fbba9da380a8b8a576['h056ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b78] =  I8a0037ad2845a3fbba9da380a8b8a576['h056f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b79] =  I8a0037ad2845a3fbba9da380a8b8a576['h056f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b7a] =  I8a0037ad2845a3fbba9da380a8b8a576['h056f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b7b] =  I8a0037ad2845a3fbba9da380a8b8a576['h056f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b7c] =  I8a0037ad2845a3fbba9da380a8b8a576['h056f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b7d] =  I8a0037ad2845a3fbba9da380a8b8a576['h056fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b7e] =  I8a0037ad2845a3fbba9da380a8b8a576['h056fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b7f] =  I8a0037ad2845a3fbba9da380a8b8a576['h056fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b80] =  I8a0037ad2845a3fbba9da380a8b8a576['h05700] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b81] =  I8a0037ad2845a3fbba9da380a8b8a576['h05702] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b82] =  I8a0037ad2845a3fbba9da380a8b8a576['h05704] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b83] =  I8a0037ad2845a3fbba9da380a8b8a576['h05706] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b84] =  I8a0037ad2845a3fbba9da380a8b8a576['h05708] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b85] =  I8a0037ad2845a3fbba9da380a8b8a576['h0570a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b86] =  I8a0037ad2845a3fbba9da380a8b8a576['h0570c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b87] =  I8a0037ad2845a3fbba9da380a8b8a576['h0570e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b88] =  I8a0037ad2845a3fbba9da380a8b8a576['h05710] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b89] =  I8a0037ad2845a3fbba9da380a8b8a576['h05712] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b8a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05714] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b8b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05716] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b8c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05718] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b8d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0571a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b8e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0571c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b8f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0571e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b90] =  I8a0037ad2845a3fbba9da380a8b8a576['h05720] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b91] =  I8a0037ad2845a3fbba9da380a8b8a576['h05722] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b92] =  I8a0037ad2845a3fbba9da380a8b8a576['h05724] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b93] =  I8a0037ad2845a3fbba9da380a8b8a576['h05726] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b94] =  I8a0037ad2845a3fbba9da380a8b8a576['h05728] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b95] =  I8a0037ad2845a3fbba9da380a8b8a576['h0572a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b96] =  I8a0037ad2845a3fbba9da380a8b8a576['h0572c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b97] =  I8a0037ad2845a3fbba9da380a8b8a576['h0572e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b98] =  I8a0037ad2845a3fbba9da380a8b8a576['h05730] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b99] =  I8a0037ad2845a3fbba9da380a8b8a576['h05732] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b9a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05734] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b9b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05736] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b9c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05738] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b9d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0573a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b9e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0573c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02b9f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0573e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ba0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05740] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ba1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05742] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ba2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05744] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ba3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05746] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ba4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05748] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ba5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0574a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ba6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0574c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ba7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0574e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ba8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05750] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ba9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05752] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02baa] =  I8a0037ad2845a3fbba9da380a8b8a576['h05754] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bab] =  I8a0037ad2845a3fbba9da380a8b8a576['h05756] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bac] =  I8a0037ad2845a3fbba9da380a8b8a576['h05758] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0575a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0575c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02baf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0575e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bb0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05760] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bb1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05762] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bb2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05764] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bb3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05766] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bb4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05768] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bb5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0576a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bb6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0576c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bb7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0576e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bb8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05770] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bb9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05772] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bba] =  I8a0037ad2845a3fbba9da380a8b8a576['h05774] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bbb] =  I8a0037ad2845a3fbba9da380a8b8a576['h05776] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bbc] =  I8a0037ad2845a3fbba9da380a8b8a576['h05778] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bbd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0577a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bbe] =  I8a0037ad2845a3fbba9da380a8b8a576['h0577c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bbf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0577e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bc0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05780] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bc1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05782] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bc2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05784] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bc3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05786] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bc4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05788] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bc5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0578a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bc6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0578c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bc7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0578e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bc8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05790] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bc9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05792] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bca] =  I8a0037ad2845a3fbba9da380a8b8a576['h05794] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bcb] =  I8a0037ad2845a3fbba9da380a8b8a576['h05796] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bcc] =  I8a0037ad2845a3fbba9da380a8b8a576['h05798] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bcd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0579a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0579c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bcf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0579e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bd0] =  I8a0037ad2845a3fbba9da380a8b8a576['h057a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bd1] =  I8a0037ad2845a3fbba9da380a8b8a576['h057a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bd2] =  I8a0037ad2845a3fbba9da380a8b8a576['h057a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bd3] =  I8a0037ad2845a3fbba9da380a8b8a576['h057a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bd4] =  I8a0037ad2845a3fbba9da380a8b8a576['h057a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bd5] =  I8a0037ad2845a3fbba9da380a8b8a576['h057aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bd6] =  I8a0037ad2845a3fbba9da380a8b8a576['h057ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bd7] =  I8a0037ad2845a3fbba9da380a8b8a576['h057ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bd8] =  I8a0037ad2845a3fbba9da380a8b8a576['h057b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bd9] =  I8a0037ad2845a3fbba9da380a8b8a576['h057b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bda] =  I8a0037ad2845a3fbba9da380a8b8a576['h057b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bdb] =  I8a0037ad2845a3fbba9da380a8b8a576['h057b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bdc] =  I8a0037ad2845a3fbba9da380a8b8a576['h057b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bdd] =  I8a0037ad2845a3fbba9da380a8b8a576['h057ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bde] =  I8a0037ad2845a3fbba9da380a8b8a576['h057bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bdf] =  I8a0037ad2845a3fbba9da380a8b8a576['h057be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02be0] =  I8a0037ad2845a3fbba9da380a8b8a576['h057c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02be1] =  I8a0037ad2845a3fbba9da380a8b8a576['h057c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02be2] =  I8a0037ad2845a3fbba9da380a8b8a576['h057c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02be3] =  I8a0037ad2845a3fbba9da380a8b8a576['h057c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02be4] =  I8a0037ad2845a3fbba9da380a8b8a576['h057c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02be5] =  I8a0037ad2845a3fbba9da380a8b8a576['h057ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02be6] =  I8a0037ad2845a3fbba9da380a8b8a576['h057cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02be7] =  I8a0037ad2845a3fbba9da380a8b8a576['h057ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02be8] =  I8a0037ad2845a3fbba9da380a8b8a576['h057d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02be9] =  I8a0037ad2845a3fbba9da380a8b8a576['h057d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bea] =  I8a0037ad2845a3fbba9da380a8b8a576['h057d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02beb] =  I8a0037ad2845a3fbba9da380a8b8a576['h057d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bec] =  I8a0037ad2845a3fbba9da380a8b8a576['h057d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bed] =  I8a0037ad2845a3fbba9da380a8b8a576['h057da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bee] =  I8a0037ad2845a3fbba9da380a8b8a576['h057dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bef] =  I8a0037ad2845a3fbba9da380a8b8a576['h057de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bf0] =  I8a0037ad2845a3fbba9da380a8b8a576['h057e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bf1] =  I8a0037ad2845a3fbba9da380a8b8a576['h057e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bf2] =  I8a0037ad2845a3fbba9da380a8b8a576['h057e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bf3] =  I8a0037ad2845a3fbba9da380a8b8a576['h057e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bf4] =  I8a0037ad2845a3fbba9da380a8b8a576['h057e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bf5] =  I8a0037ad2845a3fbba9da380a8b8a576['h057ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bf6] =  I8a0037ad2845a3fbba9da380a8b8a576['h057ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bf7] =  I8a0037ad2845a3fbba9da380a8b8a576['h057ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bf8] =  I8a0037ad2845a3fbba9da380a8b8a576['h057f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bf9] =  I8a0037ad2845a3fbba9da380a8b8a576['h057f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bfa] =  I8a0037ad2845a3fbba9da380a8b8a576['h057f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bfb] =  I8a0037ad2845a3fbba9da380a8b8a576['h057f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bfc] =  I8a0037ad2845a3fbba9da380a8b8a576['h057f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bfd] =  I8a0037ad2845a3fbba9da380a8b8a576['h057fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bfe] =  I8a0037ad2845a3fbba9da380a8b8a576['h057fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02bff] =  I8a0037ad2845a3fbba9da380a8b8a576['h057fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c00] =  I8a0037ad2845a3fbba9da380a8b8a576['h05800] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c01] =  I8a0037ad2845a3fbba9da380a8b8a576['h05802] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c02] =  I8a0037ad2845a3fbba9da380a8b8a576['h05804] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c03] =  I8a0037ad2845a3fbba9da380a8b8a576['h05806] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c04] =  I8a0037ad2845a3fbba9da380a8b8a576['h05808] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c05] =  I8a0037ad2845a3fbba9da380a8b8a576['h0580a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c06] =  I8a0037ad2845a3fbba9da380a8b8a576['h0580c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c07] =  I8a0037ad2845a3fbba9da380a8b8a576['h0580e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c08] =  I8a0037ad2845a3fbba9da380a8b8a576['h05810] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c09] =  I8a0037ad2845a3fbba9da380a8b8a576['h05812] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c0a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05814] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c0b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05816] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c0c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05818] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c0d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0581a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c0e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0581c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c0f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0581e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c10] =  I8a0037ad2845a3fbba9da380a8b8a576['h05820] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c11] =  I8a0037ad2845a3fbba9da380a8b8a576['h05822] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c12] =  I8a0037ad2845a3fbba9da380a8b8a576['h05824] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c13] =  I8a0037ad2845a3fbba9da380a8b8a576['h05826] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c14] =  I8a0037ad2845a3fbba9da380a8b8a576['h05828] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c15] =  I8a0037ad2845a3fbba9da380a8b8a576['h0582a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c16] =  I8a0037ad2845a3fbba9da380a8b8a576['h0582c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c17] =  I8a0037ad2845a3fbba9da380a8b8a576['h0582e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c18] =  I8a0037ad2845a3fbba9da380a8b8a576['h05830] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c19] =  I8a0037ad2845a3fbba9da380a8b8a576['h05832] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c1a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05834] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c1b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05836] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c1c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05838] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c1d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0583a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c1e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0583c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c1f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0583e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c20] =  I8a0037ad2845a3fbba9da380a8b8a576['h05840] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c21] =  I8a0037ad2845a3fbba9da380a8b8a576['h05842] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c22] =  I8a0037ad2845a3fbba9da380a8b8a576['h05844] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c23] =  I8a0037ad2845a3fbba9da380a8b8a576['h05846] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c24] =  I8a0037ad2845a3fbba9da380a8b8a576['h05848] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c25] =  I8a0037ad2845a3fbba9da380a8b8a576['h0584a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c26] =  I8a0037ad2845a3fbba9da380a8b8a576['h0584c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c27] =  I8a0037ad2845a3fbba9da380a8b8a576['h0584e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c28] =  I8a0037ad2845a3fbba9da380a8b8a576['h05850] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c29] =  I8a0037ad2845a3fbba9da380a8b8a576['h05852] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c2a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05854] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c2b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05856] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c2c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05858] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c2d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0585a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c2e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0585c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c2f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0585e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c30] =  I8a0037ad2845a3fbba9da380a8b8a576['h05860] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c31] =  I8a0037ad2845a3fbba9da380a8b8a576['h05862] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c32] =  I8a0037ad2845a3fbba9da380a8b8a576['h05864] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c33] =  I8a0037ad2845a3fbba9da380a8b8a576['h05866] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c34] =  I8a0037ad2845a3fbba9da380a8b8a576['h05868] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c35] =  I8a0037ad2845a3fbba9da380a8b8a576['h0586a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c36] =  I8a0037ad2845a3fbba9da380a8b8a576['h0586c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c37] =  I8a0037ad2845a3fbba9da380a8b8a576['h0586e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c38] =  I8a0037ad2845a3fbba9da380a8b8a576['h05870] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c39] =  I8a0037ad2845a3fbba9da380a8b8a576['h05872] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c3a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05874] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c3b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05876] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c3c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05878] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c3d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0587a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c3e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0587c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c3f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0587e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c40] =  I8a0037ad2845a3fbba9da380a8b8a576['h05880] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c41] =  I8a0037ad2845a3fbba9da380a8b8a576['h05882] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c42] =  I8a0037ad2845a3fbba9da380a8b8a576['h05884] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c43] =  I8a0037ad2845a3fbba9da380a8b8a576['h05886] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c44] =  I8a0037ad2845a3fbba9da380a8b8a576['h05888] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c45] =  I8a0037ad2845a3fbba9da380a8b8a576['h0588a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c46] =  I8a0037ad2845a3fbba9da380a8b8a576['h0588c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c47] =  I8a0037ad2845a3fbba9da380a8b8a576['h0588e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c48] =  I8a0037ad2845a3fbba9da380a8b8a576['h05890] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c49] =  I8a0037ad2845a3fbba9da380a8b8a576['h05892] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c4a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05894] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c4b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05896] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c4c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05898] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c4d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0589a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c4e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0589c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c4f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0589e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c50] =  I8a0037ad2845a3fbba9da380a8b8a576['h058a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c51] =  I8a0037ad2845a3fbba9da380a8b8a576['h058a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c52] =  I8a0037ad2845a3fbba9da380a8b8a576['h058a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c53] =  I8a0037ad2845a3fbba9da380a8b8a576['h058a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c54] =  I8a0037ad2845a3fbba9da380a8b8a576['h058a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c55] =  I8a0037ad2845a3fbba9da380a8b8a576['h058aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c56] =  I8a0037ad2845a3fbba9da380a8b8a576['h058ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c57] =  I8a0037ad2845a3fbba9da380a8b8a576['h058ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c58] =  I8a0037ad2845a3fbba9da380a8b8a576['h058b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c59] =  I8a0037ad2845a3fbba9da380a8b8a576['h058b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c5a] =  I8a0037ad2845a3fbba9da380a8b8a576['h058b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c5b] =  I8a0037ad2845a3fbba9da380a8b8a576['h058b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c5c] =  I8a0037ad2845a3fbba9da380a8b8a576['h058b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c5d] =  I8a0037ad2845a3fbba9da380a8b8a576['h058ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c5e] =  I8a0037ad2845a3fbba9da380a8b8a576['h058bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c5f] =  I8a0037ad2845a3fbba9da380a8b8a576['h058be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c60] =  I8a0037ad2845a3fbba9da380a8b8a576['h058c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c61] =  I8a0037ad2845a3fbba9da380a8b8a576['h058c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c62] =  I8a0037ad2845a3fbba9da380a8b8a576['h058c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c63] =  I8a0037ad2845a3fbba9da380a8b8a576['h058c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c64] =  I8a0037ad2845a3fbba9da380a8b8a576['h058c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c65] =  I8a0037ad2845a3fbba9da380a8b8a576['h058ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c66] =  I8a0037ad2845a3fbba9da380a8b8a576['h058cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c67] =  I8a0037ad2845a3fbba9da380a8b8a576['h058ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c68] =  I8a0037ad2845a3fbba9da380a8b8a576['h058d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c69] =  I8a0037ad2845a3fbba9da380a8b8a576['h058d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c6a] =  I8a0037ad2845a3fbba9da380a8b8a576['h058d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c6b] =  I8a0037ad2845a3fbba9da380a8b8a576['h058d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c6c] =  I8a0037ad2845a3fbba9da380a8b8a576['h058d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c6d] =  I8a0037ad2845a3fbba9da380a8b8a576['h058da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c6e] =  I8a0037ad2845a3fbba9da380a8b8a576['h058dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c6f] =  I8a0037ad2845a3fbba9da380a8b8a576['h058de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c70] =  I8a0037ad2845a3fbba9da380a8b8a576['h058e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c71] =  I8a0037ad2845a3fbba9da380a8b8a576['h058e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c72] =  I8a0037ad2845a3fbba9da380a8b8a576['h058e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c73] =  I8a0037ad2845a3fbba9da380a8b8a576['h058e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c74] =  I8a0037ad2845a3fbba9da380a8b8a576['h058e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c75] =  I8a0037ad2845a3fbba9da380a8b8a576['h058ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c76] =  I8a0037ad2845a3fbba9da380a8b8a576['h058ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c77] =  I8a0037ad2845a3fbba9da380a8b8a576['h058ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c78] =  I8a0037ad2845a3fbba9da380a8b8a576['h058f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c79] =  I8a0037ad2845a3fbba9da380a8b8a576['h058f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c7a] =  I8a0037ad2845a3fbba9da380a8b8a576['h058f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c7b] =  I8a0037ad2845a3fbba9da380a8b8a576['h058f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c7c] =  I8a0037ad2845a3fbba9da380a8b8a576['h058f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c7d] =  I8a0037ad2845a3fbba9da380a8b8a576['h058fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c7e] =  I8a0037ad2845a3fbba9da380a8b8a576['h058fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c7f] =  I8a0037ad2845a3fbba9da380a8b8a576['h058fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c80] =  I8a0037ad2845a3fbba9da380a8b8a576['h05900] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c81] =  I8a0037ad2845a3fbba9da380a8b8a576['h05902] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c82] =  I8a0037ad2845a3fbba9da380a8b8a576['h05904] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c83] =  I8a0037ad2845a3fbba9da380a8b8a576['h05906] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c84] =  I8a0037ad2845a3fbba9da380a8b8a576['h05908] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c85] =  I8a0037ad2845a3fbba9da380a8b8a576['h0590a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c86] =  I8a0037ad2845a3fbba9da380a8b8a576['h0590c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c87] =  I8a0037ad2845a3fbba9da380a8b8a576['h0590e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c88] =  I8a0037ad2845a3fbba9da380a8b8a576['h05910] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c89] =  I8a0037ad2845a3fbba9da380a8b8a576['h05912] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c8a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05914] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c8b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05916] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c8c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05918] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c8d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0591a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c8e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0591c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c8f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0591e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c90] =  I8a0037ad2845a3fbba9da380a8b8a576['h05920] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c91] =  I8a0037ad2845a3fbba9da380a8b8a576['h05922] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c92] =  I8a0037ad2845a3fbba9da380a8b8a576['h05924] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c93] =  I8a0037ad2845a3fbba9da380a8b8a576['h05926] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c94] =  I8a0037ad2845a3fbba9da380a8b8a576['h05928] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c95] =  I8a0037ad2845a3fbba9da380a8b8a576['h0592a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c96] =  I8a0037ad2845a3fbba9da380a8b8a576['h0592c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c97] =  I8a0037ad2845a3fbba9da380a8b8a576['h0592e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c98] =  I8a0037ad2845a3fbba9da380a8b8a576['h05930] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c99] =  I8a0037ad2845a3fbba9da380a8b8a576['h05932] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c9a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05934] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c9b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05936] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c9c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05938] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c9d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0593a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c9e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0593c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02c9f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0593e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ca0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05940] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ca1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05942] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ca2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05944] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ca3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05946] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ca4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05948] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ca5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0594a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ca6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0594c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ca7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0594e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ca8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05950] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ca9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05952] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02caa] =  I8a0037ad2845a3fbba9da380a8b8a576['h05954] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cab] =  I8a0037ad2845a3fbba9da380a8b8a576['h05956] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cac] =  I8a0037ad2845a3fbba9da380a8b8a576['h05958] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0595a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0595c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02caf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0595e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cb0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05960] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cb1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05962] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cb2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05964] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cb3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05966] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cb4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05968] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cb5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0596a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cb6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0596c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cb7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0596e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cb8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05970] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cb9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05972] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cba] =  I8a0037ad2845a3fbba9da380a8b8a576['h05974] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cbb] =  I8a0037ad2845a3fbba9da380a8b8a576['h05976] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cbc] =  I8a0037ad2845a3fbba9da380a8b8a576['h05978] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cbd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0597a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cbe] =  I8a0037ad2845a3fbba9da380a8b8a576['h0597c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cbf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0597e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cc0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05980] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cc1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05982] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cc2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05984] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cc3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05986] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cc4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05988] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cc5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0598a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cc6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0598c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cc7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0598e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cc8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05990] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cc9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05992] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cca] =  I8a0037ad2845a3fbba9da380a8b8a576['h05994] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ccb] =  I8a0037ad2845a3fbba9da380a8b8a576['h05996] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ccc] =  I8a0037ad2845a3fbba9da380a8b8a576['h05998] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ccd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0599a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0599c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ccf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0599e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cd0] =  I8a0037ad2845a3fbba9da380a8b8a576['h059a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cd1] =  I8a0037ad2845a3fbba9da380a8b8a576['h059a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cd2] =  I8a0037ad2845a3fbba9da380a8b8a576['h059a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cd3] =  I8a0037ad2845a3fbba9da380a8b8a576['h059a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cd4] =  I8a0037ad2845a3fbba9da380a8b8a576['h059a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cd5] =  I8a0037ad2845a3fbba9da380a8b8a576['h059aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cd6] =  I8a0037ad2845a3fbba9da380a8b8a576['h059ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cd7] =  I8a0037ad2845a3fbba9da380a8b8a576['h059ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cd8] =  I8a0037ad2845a3fbba9da380a8b8a576['h059b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cd9] =  I8a0037ad2845a3fbba9da380a8b8a576['h059b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cda] =  I8a0037ad2845a3fbba9da380a8b8a576['h059b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cdb] =  I8a0037ad2845a3fbba9da380a8b8a576['h059b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cdc] =  I8a0037ad2845a3fbba9da380a8b8a576['h059b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cdd] =  I8a0037ad2845a3fbba9da380a8b8a576['h059ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cde] =  I8a0037ad2845a3fbba9da380a8b8a576['h059bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cdf] =  I8a0037ad2845a3fbba9da380a8b8a576['h059be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ce0] =  I8a0037ad2845a3fbba9da380a8b8a576['h059c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ce1] =  I8a0037ad2845a3fbba9da380a8b8a576['h059c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ce2] =  I8a0037ad2845a3fbba9da380a8b8a576['h059c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ce3] =  I8a0037ad2845a3fbba9da380a8b8a576['h059c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ce4] =  I8a0037ad2845a3fbba9da380a8b8a576['h059c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ce5] =  I8a0037ad2845a3fbba9da380a8b8a576['h059ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ce6] =  I8a0037ad2845a3fbba9da380a8b8a576['h059cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ce7] =  I8a0037ad2845a3fbba9da380a8b8a576['h059ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ce8] =  I8a0037ad2845a3fbba9da380a8b8a576['h059d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ce9] =  I8a0037ad2845a3fbba9da380a8b8a576['h059d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cea] =  I8a0037ad2845a3fbba9da380a8b8a576['h059d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ceb] =  I8a0037ad2845a3fbba9da380a8b8a576['h059d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cec] =  I8a0037ad2845a3fbba9da380a8b8a576['h059d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ced] =  I8a0037ad2845a3fbba9da380a8b8a576['h059da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cee] =  I8a0037ad2845a3fbba9da380a8b8a576['h059dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cef] =  I8a0037ad2845a3fbba9da380a8b8a576['h059de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cf0] =  I8a0037ad2845a3fbba9da380a8b8a576['h059e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cf1] =  I8a0037ad2845a3fbba9da380a8b8a576['h059e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cf2] =  I8a0037ad2845a3fbba9da380a8b8a576['h059e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cf3] =  I8a0037ad2845a3fbba9da380a8b8a576['h059e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cf4] =  I8a0037ad2845a3fbba9da380a8b8a576['h059e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cf5] =  I8a0037ad2845a3fbba9da380a8b8a576['h059ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cf6] =  I8a0037ad2845a3fbba9da380a8b8a576['h059ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cf7] =  I8a0037ad2845a3fbba9da380a8b8a576['h059ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cf8] =  I8a0037ad2845a3fbba9da380a8b8a576['h059f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cf9] =  I8a0037ad2845a3fbba9da380a8b8a576['h059f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cfa] =  I8a0037ad2845a3fbba9da380a8b8a576['h059f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cfb] =  I8a0037ad2845a3fbba9da380a8b8a576['h059f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cfc] =  I8a0037ad2845a3fbba9da380a8b8a576['h059f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cfd] =  I8a0037ad2845a3fbba9da380a8b8a576['h059fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cfe] =  I8a0037ad2845a3fbba9da380a8b8a576['h059fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02cff] =  I8a0037ad2845a3fbba9da380a8b8a576['h059fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d00] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d01] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d02] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d03] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d04] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d05] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d06] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d07] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d08] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d09] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d0a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d0b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d0c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d0d] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d0e] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d0f] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d10] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d11] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d12] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d13] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d14] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d15] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d16] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d17] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d18] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d19] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d1a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d1b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d1c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d1d] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d1e] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d1f] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d20] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d21] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d22] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d23] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d24] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d25] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d26] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d27] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d28] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d29] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d2a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d2b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d2c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d2d] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d2e] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d2f] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d30] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d31] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d32] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d33] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d34] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d35] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d36] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d37] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d38] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d39] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d3a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d3b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d3c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d3d] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d3e] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d3f] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d40] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d41] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d42] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d43] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d44] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d45] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d46] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d47] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d48] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d49] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d4a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d4b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d4c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d4d] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d4e] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d4f] =  I8a0037ad2845a3fbba9da380a8b8a576['h05a9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d50] =  I8a0037ad2845a3fbba9da380a8b8a576['h05aa0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d51] =  I8a0037ad2845a3fbba9da380a8b8a576['h05aa2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d52] =  I8a0037ad2845a3fbba9da380a8b8a576['h05aa4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d53] =  I8a0037ad2845a3fbba9da380a8b8a576['h05aa6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d54] =  I8a0037ad2845a3fbba9da380a8b8a576['h05aa8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d55] =  I8a0037ad2845a3fbba9da380a8b8a576['h05aaa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d56] =  I8a0037ad2845a3fbba9da380a8b8a576['h05aac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d57] =  I8a0037ad2845a3fbba9da380a8b8a576['h05aae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d58] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ab0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d59] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ab2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d5a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ab4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d5b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ab6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d5c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ab8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d5d] =  I8a0037ad2845a3fbba9da380a8b8a576['h05aba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d5e] =  I8a0037ad2845a3fbba9da380a8b8a576['h05abc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d5f] =  I8a0037ad2845a3fbba9da380a8b8a576['h05abe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d60] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ac0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d61] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ac2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d62] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ac4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d63] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ac6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d64] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ac8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d65] =  I8a0037ad2845a3fbba9da380a8b8a576['h05aca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d66] =  I8a0037ad2845a3fbba9da380a8b8a576['h05acc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d67] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ace] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d68] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ad0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d69] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ad2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d6a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ad4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d6b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ad6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d6c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ad8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d6d] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ada] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d6e] =  I8a0037ad2845a3fbba9da380a8b8a576['h05adc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d6f] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ade] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d70] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ae0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d71] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ae2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d72] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ae4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d73] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ae6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d74] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ae8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d75] =  I8a0037ad2845a3fbba9da380a8b8a576['h05aea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d76] =  I8a0037ad2845a3fbba9da380a8b8a576['h05aec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d77] =  I8a0037ad2845a3fbba9da380a8b8a576['h05aee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d78] =  I8a0037ad2845a3fbba9da380a8b8a576['h05af0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d79] =  I8a0037ad2845a3fbba9da380a8b8a576['h05af2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d7a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05af4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d7b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05af6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d7c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05af8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d7d] =  I8a0037ad2845a3fbba9da380a8b8a576['h05afa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d7e] =  I8a0037ad2845a3fbba9da380a8b8a576['h05afc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d7f] =  I8a0037ad2845a3fbba9da380a8b8a576['h05afe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d80] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d81] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d82] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d83] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d84] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d85] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d86] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d87] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d88] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d89] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d8a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d8b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d8c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d8d] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d8e] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d8f] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d90] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d91] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d92] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d93] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d94] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d95] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d96] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d97] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d98] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d99] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d9a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d9b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d9c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d9d] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d9e] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02d9f] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02da0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02da1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02da2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02da3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02da4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02da5] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02da6] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02da7] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02da8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02da9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02daa] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dab] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dac] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dad] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dae] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02daf] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02db0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02db1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02db2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02db3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02db4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02db5] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02db6] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02db7] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02db8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02db9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dba] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dbb] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dbc] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dbd] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dbe] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dbf] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dc0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dc1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dc2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dc3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dc4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dc5] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dc6] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dc7] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dc8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dc9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dca] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dcb] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dcc] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dcd] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dce] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dcf] =  I8a0037ad2845a3fbba9da380a8b8a576['h05b9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dd0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ba0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dd1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ba2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dd2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ba4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dd3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ba6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dd4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ba8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dd5] =  I8a0037ad2845a3fbba9da380a8b8a576['h05baa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dd6] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dd7] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dd8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dd9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dda] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ddb] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ddc] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ddd] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dde] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ddf] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02de0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02de1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02de2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02de3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02de4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02de5] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02de6] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bcc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02de7] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02de8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02de9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dea] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02deb] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dec] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ded] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dee] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bdc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02def] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02df0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05be0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02df1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05be2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02df2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05be4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02df3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05be6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02df4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05be8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02df5] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02df6] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02df7] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02df8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bf0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02df9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bf2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dfa] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bf4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dfb] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bf6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dfc] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bf8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dfd] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bfa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dfe] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bfc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02dff] =  I8a0037ad2845a3fbba9da380a8b8a576['h05bfe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e00] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e01] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e02] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e03] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e04] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e05] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e06] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e07] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e08] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e09] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e0a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e0b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e0c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e0d] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e0e] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e0f] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e10] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e11] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e12] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e13] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e14] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e15] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e16] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e17] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e18] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e19] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e1a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e1b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e1c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e1d] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e1e] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e1f] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e20] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e21] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e22] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e23] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e24] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e25] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e26] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e27] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e28] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e29] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e2a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e2b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e2c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e2d] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e2e] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e2f] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e30] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e31] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e32] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e33] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e34] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e35] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e36] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e37] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e38] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e39] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e3a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e3b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e3c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e3d] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e3e] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e3f] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e40] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e41] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e42] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e43] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e44] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e45] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e46] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e47] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e48] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e49] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e4a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e4b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e4c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e4d] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e4e] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e4f] =  I8a0037ad2845a3fbba9da380a8b8a576['h05c9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e50] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ca0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e51] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ca2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e52] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ca4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e53] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ca6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e54] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ca8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e55] =  I8a0037ad2845a3fbba9da380a8b8a576['h05caa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e56] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e57] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e58] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e59] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e5a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e5b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e5c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e5d] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e5e] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e5f] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e60] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e61] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e62] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e63] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e64] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e65] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e66] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ccc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e67] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e68] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e69] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e6a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e6b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e6c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e6d] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e6e] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cdc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e6f] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e70] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ce0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e71] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ce2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e72] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ce4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e73] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ce6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e74] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ce8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e75] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e76] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e77] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e78] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cf0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e79] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cf2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e7a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cf4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e7b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cf6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e7c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cf8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e7d] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cfa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e7e] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cfc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e7f] =  I8a0037ad2845a3fbba9da380a8b8a576['h05cfe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e80] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e81] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e82] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e83] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e84] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e85] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e86] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e87] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e88] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e89] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e8a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e8b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e8c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e8d] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e8e] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e8f] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e90] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e91] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e92] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e93] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e94] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e95] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e96] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e97] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e98] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e99] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e9a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e9b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e9c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e9d] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e9e] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02e9f] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ea0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ea1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ea2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ea3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ea4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ea5] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ea6] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ea7] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ea8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ea9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02eaa] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02eab] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02eac] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ead] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02eae] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02eaf] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02eb0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02eb1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02eb2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02eb3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02eb4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02eb5] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02eb6] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02eb7] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02eb8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02eb9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02eba] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ebb] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ebc] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ebd] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ebe] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ebf] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ec0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ec1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ec2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ec3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ec4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ec5] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ec6] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ec7] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ec8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ec9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02eca] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ecb] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ecc] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ecd] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ece] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ecf] =  I8a0037ad2845a3fbba9da380a8b8a576['h05d9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ed0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05da0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ed1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05da2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ed2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05da4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ed3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05da6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ed4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05da8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ed5] =  I8a0037ad2845a3fbba9da380a8b8a576['h05daa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ed6] =  I8a0037ad2845a3fbba9da380a8b8a576['h05dac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ed7] =  I8a0037ad2845a3fbba9da380a8b8a576['h05dae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ed8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05db0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ed9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05db2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02eda] =  I8a0037ad2845a3fbba9da380a8b8a576['h05db4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02edb] =  I8a0037ad2845a3fbba9da380a8b8a576['h05db6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02edc] =  I8a0037ad2845a3fbba9da380a8b8a576['h05db8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02edd] =  I8a0037ad2845a3fbba9da380a8b8a576['h05dba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ede] =  I8a0037ad2845a3fbba9da380a8b8a576['h05dbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02edf] =  I8a0037ad2845a3fbba9da380a8b8a576['h05dbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ee0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05dc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ee1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05dc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ee2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05dc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ee3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05dc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ee4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05dc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ee5] =  I8a0037ad2845a3fbba9da380a8b8a576['h05dca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ee6] =  I8a0037ad2845a3fbba9da380a8b8a576['h05dcc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ee7] =  I8a0037ad2845a3fbba9da380a8b8a576['h05dce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ee8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05dd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ee9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05dd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02eea] =  I8a0037ad2845a3fbba9da380a8b8a576['h05dd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02eeb] =  I8a0037ad2845a3fbba9da380a8b8a576['h05dd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02eec] =  I8a0037ad2845a3fbba9da380a8b8a576['h05dd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02eed] =  I8a0037ad2845a3fbba9da380a8b8a576['h05dda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02eee] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ddc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02eef] =  I8a0037ad2845a3fbba9da380a8b8a576['h05dde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ef0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05de0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ef1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05de2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ef2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05de4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ef3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05de6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ef4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05de8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ef5] =  I8a0037ad2845a3fbba9da380a8b8a576['h05dea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ef6] =  I8a0037ad2845a3fbba9da380a8b8a576['h05dec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ef7] =  I8a0037ad2845a3fbba9da380a8b8a576['h05dee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ef8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05df0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ef9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05df2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02efa] =  I8a0037ad2845a3fbba9da380a8b8a576['h05df4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02efb] =  I8a0037ad2845a3fbba9da380a8b8a576['h05df6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02efc] =  I8a0037ad2845a3fbba9da380a8b8a576['h05df8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02efd] =  I8a0037ad2845a3fbba9da380a8b8a576['h05dfa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02efe] =  I8a0037ad2845a3fbba9da380a8b8a576['h05dfc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02eff] =  I8a0037ad2845a3fbba9da380a8b8a576['h05dfe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f00] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f01] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f02] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f03] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f04] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f05] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f06] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f07] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f08] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f09] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f0a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f0b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f0c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f0d] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f0e] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f0f] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f10] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f11] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f12] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f13] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f14] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f15] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f16] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f17] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f18] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f19] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f1a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f1b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f1c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f1d] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f1e] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f1f] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f20] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f21] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f22] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f23] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f24] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f25] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f26] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f27] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f28] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f29] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f2a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f2b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f2c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f2d] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f2e] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f2f] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f30] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f31] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f32] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f33] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f34] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f35] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f36] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f37] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f38] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f39] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f3a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f3b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f3c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f3d] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f3e] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f3f] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f40] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f41] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f42] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f43] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f44] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f45] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f46] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f47] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f48] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f49] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f4a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f4b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f4c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f4d] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f4e] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f4f] =  I8a0037ad2845a3fbba9da380a8b8a576['h05e9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f50] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ea0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f51] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ea2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f52] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ea4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f53] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ea6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f54] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ea8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f55] =  I8a0037ad2845a3fbba9da380a8b8a576['h05eaa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f56] =  I8a0037ad2845a3fbba9da380a8b8a576['h05eac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f57] =  I8a0037ad2845a3fbba9da380a8b8a576['h05eae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f58] =  I8a0037ad2845a3fbba9da380a8b8a576['h05eb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f59] =  I8a0037ad2845a3fbba9da380a8b8a576['h05eb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f5a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05eb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f5b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05eb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f5c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05eb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f5d] =  I8a0037ad2845a3fbba9da380a8b8a576['h05eba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f5e] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ebc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f5f] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ebe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f60] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ec0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f61] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ec2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f62] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ec4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f63] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ec6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f64] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ec8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f65] =  I8a0037ad2845a3fbba9da380a8b8a576['h05eca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f66] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ecc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f67] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ece] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f68] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ed0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f69] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ed2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f6a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ed4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f6b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ed6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f6c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ed8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f6d] =  I8a0037ad2845a3fbba9da380a8b8a576['h05eda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f6e] =  I8a0037ad2845a3fbba9da380a8b8a576['h05edc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f6f] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ede] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f70] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ee0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f71] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ee2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f72] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ee4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f73] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ee6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f74] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ee8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f75] =  I8a0037ad2845a3fbba9da380a8b8a576['h05eea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f76] =  I8a0037ad2845a3fbba9da380a8b8a576['h05eec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f77] =  I8a0037ad2845a3fbba9da380a8b8a576['h05eee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f78] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ef0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f79] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ef2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f7a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ef4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f7b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ef6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f7c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ef8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f7d] =  I8a0037ad2845a3fbba9da380a8b8a576['h05efa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f7e] =  I8a0037ad2845a3fbba9da380a8b8a576['h05efc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f7f] =  I8a0037ad2845a3fbba9da380a8b8a576['h05efe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f80] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f81] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f82] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f83] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f84] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f85] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f86] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f87] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f88] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f89] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f8a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f8b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f8c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f8d] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f8e] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f8f] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f90] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f91] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f92] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f93] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f94] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f95] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f96] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f97] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f98] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f99] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f9a] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f9b] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f9c] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f9d] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f9e] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02f9f] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fa0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fa1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fa2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fa3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fa4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fa5] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fa6] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fa7] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fa8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fa9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02faa] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fab] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fac] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fad] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fae] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02faf] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fb0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fb1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fb2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fb3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fb4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fb5] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fb6] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fb7] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fb8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fb9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fba] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fbb] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fbc] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fbd] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fbe] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fbf] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fc0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fc1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fc2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fc3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fc4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fc5] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fc6] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fc7] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fc8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fc9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fca] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fcb] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fcc] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fcd] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fce] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fcf] =  I8a0037ad2845a3fbba9da380a8b8a576['h05f9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fd0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fa0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fd1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fa2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fd2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fa4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fd3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fa6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fd4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fa8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fd5] =  I8a0037ad2845a3fbba9da380a8b8a576['h05faa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fd6] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fd7] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fd8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fd9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fda] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fdb] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fdc] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fdd] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fde] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fdf] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fe0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fe1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fe2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fe3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fe4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fe5] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fe6] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fcc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fe7] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fe8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fe9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fea] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02feb] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fec] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fed] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fee] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fdc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fef] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ff0] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fe0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ff1] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fe2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ff2] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fe4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ff3] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fe6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ff4] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fe8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ff5] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ff6] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ff7] =  I8a0037ad2845a3fbba9da380a8b8a576['h05fee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ff8] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ff0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ff9] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ff2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ffa] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ff4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ffb] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ff6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ffc] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ff8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ffd] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ffa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02ffe] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ffc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h02fff] =  I8a0037ad2845a3fbba9da380a8b8a576['h05ffe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03000] =  I8a0037ad2845a3fbba9da380a8b8a576['h06000] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03001] =  I8a0037ad2845a3fbba9da380a8b8a576['h06002] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03002] =  I8a0037ad2845a3fbba9da380a8b8a576['h06004] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03003] =  I8a0037ad2845a3fbba9da380a8b8a576['h06006] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03004] =  I8a0037ad2845a3fbba9da380a8b8a576['h06008] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03005] =  I8a0037ad2845a3fbba9da380a8b8a576['h0600a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03006] =  I8a0037ad2845a3fbba9da380a8b8a576['h0600c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03007] =  I8a0037ad2845a3fbba9da380a8b8a576['h0600e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03008] =  I8a0037ad2845a3fbba9da380a8b8a576['h06010] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03009] =  I8a0037ad2845a3fbba9da380a8b8a576['h06012] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0300a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06014] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0300b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06016] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0300c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06018] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0300d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0601a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0300e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0601c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0300f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0601e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03010] =  I8a0037ad2845a3fbba9da380a8b8a576['h06020] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03011] =  I8a0037ad2845a3fbba9da380a8b8a576['h06022] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03012] =  I8a0037ad2845a3fbba9da380a8b8a576['h06024] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03013] =  I8a0037ad2845a3fbba9da380a8b8a576['h06026] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03014] =  I8a0037ad2845a3fbba9da380a8b8a576['h06028] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03015] =  I8a0037ad2845a3fbba9da380a8b8a576['h0602a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03016] =  I8a0037ad2845a3fbba9da380a8b8a576['h0602c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03017] =  I8a0037ad2845a3fbba9da380a8b8a576['h0602e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03018] =  I8a0037ad2845a3fbba9da380a8b8a576['h06030] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03019] =  I8a0037ad2845a3fbba9da380a8b8a576['h06032] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0301a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06034] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0301b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06036] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0301c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06038] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0301d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0603a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0301e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0603c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0301f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0603e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03020] =  I8a0037ad2845a3fbba9da380a8b8a576['h06040] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03021] =  I8a0037ad2845a3fbba9da380a8b8a576['h06042] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03022] =  I8a0037ad2845a3fbba9da380a8b8a576['h06044] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03023] =  I8a0037ad2845a3fbba9da380a8b8a576['h06046] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03024] =  I8a0037ad2845a3fbba9da380a8b8a576['h06048] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03025] =  I8a0037ad2845a3fbba9da380a8b8a576['h0604a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03026] =  I8a0037ad2845a3fbba9da380a8b8a576['h0604c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03027] =  I8a0037ad2845a3fbba9da380a8b8a576['h0604e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03028] =  I8a0037ad2845a3fbba9da380a8b8a576['h06050] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03029] =  I8a0037ad2845a3fbba9da380a8b8a576['h06052] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0302a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06054] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0302b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06056] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0302c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06058] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0302d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0605a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0302e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0605c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0302f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0605e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03030] =  I8a0037ad2845a3fbba9da380a8b8a576['h06060] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03031] =  I8a0037ad2845a3fbba9da380a8b8a576['h06062] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03032] =  I8a0037ad2845a3fbba9da380a8b8a576['h06064] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03033] =  I8a0037ad2845a3fbba9da380a8b8a576['h06066] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03034] =  I8a0037ad2845a3fbba9da380a8b8a576['h06068] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03035] =  I8a0037ad2845a3fbba9da380a8b8a576['h0606a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03036] =  I8a0037ad2845a3fbba9da380a8b8a576['h0606c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03037] =  I8a0037ad2845a3fbba9da380a8b8a576['h0606e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03038] =  I8a0037ad2845a3fbba9da380a8b8a576['h06070] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03039] =  I8a0037ad2845a3fbba9da380a8b8a576['h06072] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0303a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06074] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0303b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06076] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0303c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06078] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0303d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0607a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0303e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0607c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0303f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0607e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03040] =  I8a0037ad2845a3fbba9da380a8b8a576['h06080] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03041] =  I8a0037ad2845a3fbba9da380a8b8a576['h06082] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03042] =  I8a0037ad2845a3fbba9da380a8b8a576['h06084] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03043] =  I8a0037ad2845a3fbba9da380a8b8a576['h06086] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03044] =  I8a0037ad2845a3fbba9da380a8b8a576['h06088] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03045] =  I8a0037ad2845a3fbba9da380a8b8a576['h0608a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03046] =  I8a0037ad2845a3fbba9da380a8b8a576['h0608c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03047] =  I8a0037ad2845a3fbba9da380a8b8a576['h0608e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03048] =  I8a0037ad2845a3fbba9da380a8b8a576['h06090] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03049] =  I8a0037ad2845a3fbba9da380a8b8a576['h06092] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0304a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06094] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0304b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06096] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0304c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06098] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0304d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0609a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0304e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0609c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0304f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0609e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03050] =  I8a0037ad2845a3fbba9da380a8b8a576['h060a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03051] =  I8a0037ad2845a3fbba9da380a8b8a576['h060a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03052] =  I8a0037ad2845a3fbba9da380a8b8a576['h060a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03053] =  I8a0037ad2845a3fbba9da380a8b8a576['h060a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03054] =  I8a0037ad2845a3fbba9da380a8b8a576['h060a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03055] =  I8a0037ad2845a3fbba9da380a8b8a576['h060aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03056] =  I8a0037ad2845a3fbba9da380a8b8a576['h060ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03057] =  I8a0037ad2845a3fbba9da380a8b8a576['h060ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03058] =  I8a0037ad2845a3fbba9da380a8b8a576['h060b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03059] =  I8a0037ad2845a3fbba9da380a8b8a576['h060b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0305a] =  I8a0037ad2845a3fbba9da380a8b8a576['h060b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0305b] =  I8a0037ad2845a3fbba9da380a8b8a576['h060b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0305c] =  I8a0037ad2845a3fbba9da380a8b8a576['h060b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0305d] =  I8a0037ad2845a3fbba9da380a8b8a576['h060ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0305e] =  I8a0037ad2845a3fbba9da380a8b8a576['h060bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0305f] =  I8a0037ad2845a3fbba9da380a8b8a576['h060be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03060] =  I8a0037ad2845a3fbba9da380a8b8a576['h060c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03061] =  I8a0037ad2845a3fbba9da380a8b8a576['h060c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03062] =  I8a0037ad2845a3fbba9da380a8b8a576['h060c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03063] =  I8a0037ad2845a3fbba9da380a8b8a576['h060c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03064] =  I8a0037ad2845a3fbba9da380a8b8a576['h060c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03065] =  I8a0037ad2845a3fbba9da380a8b8a576['h060ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03066] =  I8a0037ad2845a3fbba9da380a8b8a576['h060cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03067] =  I8a0037ad2845a3fbba9da380a8b8a576['h060ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03068] =  I8a0037ad2845a3fbba9da380a8b8a576['h060d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03069] =  I8a0037ad2845a3fbba9da380a8b8a576['h060d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0306a] =  I8a0037ad2845a3fbba9da380a8b8a576['h060d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0306b] =  I8a0037ad2845a3fbba9da380a8b8a576['h060d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0306c] =  I8a0037ad2845a3fbba9da380a8b8a576['h060d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0306d] =  I8a0037ad2845a3fbba9da380a8b8a576['h060da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0306e] =  I8a0037ad2845a3fbba9da380a8b8a576['h060dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0306f] =  I8a0037ad2845a3fbba9da380a8b8a576['h060de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03070] =  I8a0037ad2845a3fbba9da380a8b8a576['h060e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03071] =  I8a0037ad2845a3fbba9da380a8b8a576['h060e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03072] =  I8a0037ad2845a3fbba9da380a8b8a576['h060e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03073] =  I8a0037ad2845a3fbba9da380a8b8a576['h060e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03074] =  I8a0037ad2845a3fbba9da380a8b8a576['h060e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03075] =  I8a0037ad2845a3fbba9da380a8b8a576['h060ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03076] =  I8a0037ad2845a3fbba9da380a8b8a576['h060ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03077] =  I8a0037ad2845a3fbba9da380a8b8a576['h060ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03078] =  I8a0037ad2845a3fbba9da380a8b8a576['h060f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03079] =  I8a0037ad2845a3fbba9da380a8b8a576['h060f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0307a] =  I8a0037ad2845a3fbba9da380a8b8a576['h060f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0307b] =  I8a0037ad2845a3fbba9da380a8b8a576['h060f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0307c] =  I8a0037ad2845a3fbba9da380a8b8a576['h060f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0307d] =  I8a0037ad2845a3fbba9da380a8b8a576['h060fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0307e] =  I8a0037ad2845a3fbba9da380a8b8a576['h060fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0307f] =  I8a0037ad2845a3fbba9da380a8b8a576['h060fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03080] =  I8a0037ad2845a3fbba9da380a8b8a576['h06100] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03081] =  I8a0037ad2845a3fbba9da380a8b8a576['h06102] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03082] =  I8a0037ad2845a3fbba9da380a8b8a576['h06104] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03083] =  I8a0037ad2845a3fbba9da380a8b8a576['h06106] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03084] =  I8a0037ad2845a3fbba9da380a8b8a576['h06108] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03085] =  I8a0037ad2845a3fbba9da380a8b8a576['h0610a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03086] =  I8a0037ad2845a3fbba9da380a8b8a576['h0610c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03087] =  I8a0037ad2845a3fbba9da380a8b8a576['h0610e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03088] =  I8a0037ad2845a3fbba9da380a8b8a576['h06110] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03089] =  I8a0037ad2845a3fbba9da380a8b8a576['h06112] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0308a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06114] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0308b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06116] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0308c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06118] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0308d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0611a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0308e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0611c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0308f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0611e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03090] =  I8a0037ad2845a3fbba9da380a8b8a576['h06120] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03091] =  I8a0037ad2845a3fbba9da380a8b8a576['h06122] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03092] =  I8a0037ad2845a3fbba9da380a8b8a576['h06124] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03093] =  I8a0037ad2845a3fbba9da380a8b8a576['h06126] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03094] =  I8a0037ad2845a3fbba9da380a8b8a576['h06128] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03095] =  I8a0037ad2845a3fbba9da380a8b8a576['h0612a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03096] =  I8a0037ad2845a3fbba9da380a8b8a576['h0612c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03097] =  I8a0037ad2845a3fbba9da380a8b8a576['h0612e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03098] =  I8a0037ad2845a3fbba9da380a8b8a576['h06130] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03099] =  I8a0037ad2845a3fbba9da380a8b8a576['h06132] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0309a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06134] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0309b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06136] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0309c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06138] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0309d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0613a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0309e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0613c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0309f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0613e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06140] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06142] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06144] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06146] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06148] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0614a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0614c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0614e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06150] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06152] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h06154] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h06156] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h06158] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0615a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0615c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030af] =  I8a0037ad2845a3fbba9da380a8b8a576['h0615e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06160] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06162] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06164] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06166] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06168] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0616a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0616c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0616e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06170] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06172] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h06174] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h06176] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h06178] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0617a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030be] =  I8a0037ad2845a3fbba9da380a8b8a576['h0617c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0617e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06180] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06182] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06184] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06186] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06188] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0618a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0618c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0618e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06190] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06192] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h06194] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h06196] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h06198] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0619a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0619c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0619e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h061a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h061a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h061a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h061a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h061a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h061aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h061ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h061ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h061b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h061b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030da] =  I8a0037ad2845a3fbba9da380a8b8a576['h061b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030db] =  I8a0037ad2845a3fbba9da380a8b8a576['h061b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h061b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h061ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030de] =  I8a0037ad2845a3fbba9da380a8b8a576['h061bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030df] =  I8a0037ad2845a3fbba9da380a8b8a576['h061be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h061c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h061c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h061c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h061c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h061c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h061ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h061cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h061ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h061d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h061d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h061d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h061d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h061d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h061da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h061dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h061de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h061e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h061e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h061e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h061e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h061e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h061ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h061ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h061ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h061f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h061f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h061f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h061f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h061f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h061fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h061fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h030ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h061fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03100] =  I8a0037ad2845a3fbba9da380a8b8a576['h06200] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03101] =  I8a0037ad2845a3fbba9da380a8b8a576['h06202] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03102] =  I8a0037ad2845a3fbba9da380a8b8a576['h06204] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03103] =  I8a0037ad2845a3fbba9da380a8b8a576['h06206] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03104] =  I8a0037ad2845a3fbba9da380a8b8a576['h06208] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03105] =  I8a0037ad2845a3fbba9da380a8b8a576['h0620a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03106] =  I8a0037ad2845a3fbba9da380a8b8a576['h0620c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03107] =  I8a0037ad2845a3fbba9da380a8b8a576['h0620e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03108] =  I8a0037ad2845a3fbba9da380a8b8a576['h06210] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03109] =  I8a0037ad2845a3fbba9da380a8b8a576['h06212] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0310a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06214] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0310b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06216] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0310c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06218] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0310d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0621a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0310e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0621c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0310f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0621e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03110] =  I8a0037ad2845a3fbba9da380a8b8a576['h06220] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03111] =  I8a0037ad2845a3fbba9da380a8b8a576['h06222] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03112] =  I8a0037ad2845a3fbba9da380a8b8a576['h06224] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03113] =  I8a0037ad2845a3fbba9da380a8b8a576['h06226] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03114] =  I8a0037ad2845a3fbba9da380a8b8a576['h06228] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03115] =  I8a0037ad2845a3fbba9da380a8b8a576['h0622a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03116] =  I8a0037ad2845a3fbba9da380a8b8a576['h0622c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03117] =  I8a0037ad2845a3fbba9da380a8b8a576['h0622e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03118] =  I8a0037ad2845a3fbba9da380a8b8a576['h06230] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03119] =  I8a0037ad2845a3fbba9da380a8b8a576['h06232] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0311a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06234] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0311b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06236] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0311c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06238] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0311d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0623a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0311e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0623c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0311f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0623e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03120] =  I8a0037ad2845a3fbba9da380a8b8a576['h06240] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03121] =  I8a0037ad2845a3fbba9da380a8b8a576['h06242] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03122] =  I8a0037ad2845a3fbba9da380a8b8a576['h06244] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03123] =  I8a0037ad2845a3fbba9da380a8b8a576['h06246] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03124] =  I8a0037ad2845a3fbba9da380a8b8a576['h06248] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03125] =  I8a0037ad2845a3fbba9da380a8b8a576['h0624a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03126] =  I8a0037ad2845a3fbba9da380a8b8a576['h0624c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03127] =  I8a0037ad2845a3fbba9da380a8b8a576['h0624e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03128] =  I8a0037ad2845a3fbba9da380a8b8a576['h06250] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03129] =  I8a0037ad2845a3fbba9da380a8b8a576['h06252] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0312a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06254] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0312b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06256] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0312c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06258] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0312d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0625a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0312e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0625c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0312f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0625e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03130] =  I8a0037ad2845a3fbba9da380a8b8a576['h06260] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03131] =  I8a0037ad2845a3fbba9da380a8b8a576['h06262] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03132] =  I8a0037ad2845a3fbba9da380a8b8a576['h06264] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03133] =  I8a0037ad2845a3fbba9da380a8b8a576['h06266] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03134] =  I8a0037ad2845a3fbba9da380a8b8a576['h06268] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03135] =  I8a0037ad2845a3fbba9da380a8b8a576['h0626a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03136] =  I8a0037ad2845a3fbba9da380a8b8a576['h0626c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03137] =  I8a0037ad2845a3fbba9da380a8b8a576['h0626e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03138] =  I8a0037ad2845a3fbba9da380a8b8a576['h06270] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03139] =  I8a0037ad2845a3fbba9da380a8b8a576['h06272] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0313a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06274] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0313b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06276] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0313c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06278] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0313d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0627a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0313e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0627c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0313f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0627e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03140] =  I8a0037ad2845a3fbba9da380a8b8a576['h06280] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03141] =  I8a0037ad2845a3fbba9da380a8b8a576['h06282] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03142] =  I8a0037ad2845a3fbba9da380a8b8a576['h06284] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03143] =  I8a0037ad2845a3fbba9da380a8b8a576['h06286] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03144] =  I8a0037ad2845a3fbba9da380a8b8a576['h06288] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03145] =  I8a0037ad2845a3fbba9da380a8b8a576['h0628a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03146] =  I8a0037ad2845a3fbba9da380a8b8a576['h0628c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03147] =  I8a0037ad2845a3fbba9da380a8b8a576['h0628e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03148] =  I8a0037ad2845a3fbba9da380a8b8a576['h06290] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03149] =  I8a0037ad2845a3fbba9da380a8b8a576['h06292] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0314a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06294] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0314b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06296] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0314c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06298] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0314d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0629a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0314e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0629c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0314f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0629e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03150] =  I8a0037ad2845a3fbba9da380a8b8a576['h062a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03151] =  I8a0037ad2845a3fbba9da380a8b8a576['h062a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03152] =  I8a0037ad2845a3fbba9da380a8b8a576['h062a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03153] =  I8a0037ad2845a3fbba9da380a8b8a576['h062a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03154] =  I8a0037ad2845a3fbba9da380a8b8a576['h062a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03155] =  I8a0037ad2845a3fbba9da380a8b8a576['h062aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03156] =  I8a0037ad2845a3fbba9da380a8b8a576['h062ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03157] =  I8a0037ad2845a3fbba9da380a8b8a576['h062ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03158] =  I8a0037ad2845a3fbba9da380a8b8a576['h062b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03159] =  I8a0037ad2845a3fbba9da380a8b8a576['h062b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0315a] =  I8a0037ad2845a3fbba9da380a8b8a576['h062b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0315b] =  I8a0037ad2845a3fbba9da380a8b8a576['h062b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0315c] =  I8a0037ad2845a3fbba9da380a8b8a576['h062b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0315d] =  I8a0037ad2845a3fbba9da380a8b8a576['h062ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0315e] =  I8a0037ad2845a3fbba9da380a8b8a576['h062bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0315f] =  I8a0037ad2845a3fbba9da380a8b8a576['h062be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03160] =  I8a0037ad2845a3fbba9da380a8b8a576['h062c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03161] =  I8a0037ad2845a3fbba9da380a8b8a576['h062c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03162] =  I8a0037ad2845a3fbba9da380a8b8a576['h062c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03163] =  I8a0037ad2845a3fbba9da380a8b8a576['h062c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03164] =  I8a0037ad2845a3fbba9da380a8b8a576['h062c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03165] =  I8a0037ad2845a3fbba9da380a8b8a576['h062ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03166] =  I8a0037ad2845a3fbba9da380a8b8a576['h062cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03167] =  I8a0037ad2845a3fbba9da380a8b8a576['h062ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03168] =  I8a0037ad2845a3fbba9da380a8b8a576['h062d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03169] =  I8a0037ad2845a3fbba9da380a8b8a576['h062d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0316a] =  I8a0037ad2845a3fbba9da380a8b8a576['h062d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0316b] =  I8a0037ad2845a3fbba9da380a8b8a576['h062d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0316c] =  I8a0037ad2845a3fbba9da380a8b8a576['h062d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0316d] =  I8a0037ad2845a3fbba9da380a8b8a576['h062da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0316e] =  I8a0037ad2845a3fbba9da380a8b8a576['h062dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0316f] =  I8a0037ad2845a3fbba9da380a8b8a576['h062de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03170] =  I8a0037ad2845a3fbba9da380a8b8a576['h062e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03171] =  I8a0037ad2845a3fbba9da380a8b8a576['h062e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03172] =  I8a0037ad2845a3fbba9da380a8b8a576['h062e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03173] =  I8a0037ad2845a3fbba9da380a8b8a576['h062e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03174] =  I8a0037ad2845a3fbba9da380a8b8a576['h062e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03175] =  I8a0037ad2845a3fbba9da380a8b8a576['h062ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03176] =  I8a0037ad2845a3fbba9da380a8b8a576['h062ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03177] =  I8a0037ad2845a3fbba9da380a8b8a576['h062ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03178] =  I8a0037ad2845a3fbba9da380a8b8a576['h062f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03179] =  I8a0037ad2845a3fbba9da380a8b8a576['h062f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0317a] =  I8a0037ad2845a3fbba9da380a8b8a576['h062f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0317b] =  I8a0037ad2845a3fbba9da380a8b8a576['h062f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0317c] =  I8a0037ad2845a3fbba9da380a8b8a576['h062f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0317d] =  I8a0037ad2845a3fbba9da380a8b8a576['h062fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0317e] =  I8a0037ad2845a3fbba9da380a8b8a576['h062fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0317f] =  I8a0037ad2845a3fbba9da380a8b8a576['h062fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03180] =  I8a0037ad2845a3fbba9da380a8b8a576['h06300] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03181] =  I8a0037ad2845a3fbba9da380a8b8a576['h06302] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03182] =  I8a0037ad2845a3fbba9da380a8b8a576['h06304] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03183] =  I8a0037ad2845a3fbba9da380a8b8a576['h06306] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03184] =  I8a0037ad2845a3fbba9da380a8b8a576['h06308] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03185] =  I8a0037ad2845a3fbba9da380a8b8a576['h0630a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03186] =  I8a0037ad2845a3fbba9da380a8b8a576['h0630c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03187] =  I8a0037ad2845a3fbba9da380a8b8a576['h0630e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03188] =  I8a0037ad2845a3fbba9da380a8b8a576['h06310] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03189] =  I8a0037ad2845a3fbba9da380a8b8a576['h06312] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0318a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06314] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0318b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06316] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0318c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06318] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0318d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0631a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0318e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0631c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0318f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0631e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03190] =  I8a0037ad2845a3fbba9da380a8b8a576['h06320] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03191] =  I8a0037ad2845a3fbba9da380a8b8a576['h06322] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03192] =  I8a0037ad2845a3fbba9da380a8b8a576['h06324] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03193] =  I8a0037ad2845a3fbba9da380a8b8a576['h06326] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03194] =  I8a0037ad2845a3fbba9da380a8b8a576['h06328] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03195] =  I8a0037ad2845a3fbba9da380a8b8a576['h0632a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03196] =  I8a0037ad2845a3fbba9da380a8b8a576['h0632c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03197] =  I8a0037ad2845a3fbba9da380a8b8a576['h0632e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03198] =  I8a0037ad2845a3fbba9da380a8b8a576['h06330] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03199] =  I8a0037ad2845a3fbba9da380a8b8a576['h06332] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0319a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06334] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0319b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06336] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0319c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06338] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0319d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0633a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0319e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0633c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0319f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0633e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06340] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06342] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06344] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06346] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06348] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0634a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0634c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0634e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06350] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06352] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h06354] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h06356] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h06358] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0635a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0635c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031af] =  I8a0037ad2845a3fbba9da380a8b8a576['h0635e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06360] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06362] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06364] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06366] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06368] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0636a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0636c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0636e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06370] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06372] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h06374] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h06376] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h06378] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0637a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031be] =  I8a0037ad2845a3fbba9da380a8b8a576['h0637c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0637e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06380] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06382] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06384] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06386] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06388] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0638a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0638c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0638e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06390] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06392] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h06394] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h06396] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h06398] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0639a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0639c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0639e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h063a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h063a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h063a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h063a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h063a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h063aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h063ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h063ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h063b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h063b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031da] =  I8a0037ad2845a3fbba9da380a8b8a576['h063b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031db] =  I8a0037ad2845a3fbba9da380a8b8a576['h063b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h063b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h063ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031de] =  I8a0037ad2845a3fbba9da380a8b8a576['h063bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031df] =  I8a0037ad2845a3fbba9da380a8b8a576['h063be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h063c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h063c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h063c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h063c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h063c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h063ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h063cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h063ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h063d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h063d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h063d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h063d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h063d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h063da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h063dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h063de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h063e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h063e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h063e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h063e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h063e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h063ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h063ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h063ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h063f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h063f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h063f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h063f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h063f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h063fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h063fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h031ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h063fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03200] =  I8a0037ad2845a3fbba9da380a8b8a576['h06400] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03201] =  I8a0037ad2845a3fbba9da380a8b8a576['h06402] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03202] =  I8a0037ad2845a3fbba9da380a8b8a576['h06404] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03203] =  I8a0037ad2845a3fbba9da380a8b8a576['h06406] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03204] =  I8a0037ad2845a3fbba9da380a8b8a576['h06408] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03205] =  I8a0037ad2845a3fbba9da380a8b8a576['h0640a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03206] =  I8a0037ad2845a3fbba9da380a8b8a576['h0640c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03207] =  I8a0037ad2845a3fbba9da380a8b8a576['h0640e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03208] =  I8a0037ad2845a3fbba9da380a8b8a576['h06410] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03209] =  I8a0037ad2845a3fbba9da380a8b8a576['h06412] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0320a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06414] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0320b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06416] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0320c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06418] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0320d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0641a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0320e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0641c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0320f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0641e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03210] =  I8a0037ad2845a3fbba9da380a8b8a576['h06420] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03211] =  I8a0037ad2845a3fbba9da380a8b8a576['h06422] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03212] =  I8a0037ad2845a3fbba9da380a8b8a576['h06424] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03213] =  I8a0037ad2845a3fbba9da380a8b8a576['h06426] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03214] =  I8a0037ad2845a3fbba9da380a8b8a576['h06428] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03215] =  I8a0037ad2845a3fbba9da380a8b8a576['h0642a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03216] =  I8a0037ad2845a3fbba9da380a8b8a576['h0642c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03217] =  I8a0037ad2845a3fbba9da380a8b8a576['h0642e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03218] =  I8a0037ad2845a3fbba9da380a8b8a576['h06430] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03219] =  I8a0037ad2845a3fbba9da380a8b8a576['h06432] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0321a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06434] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0321b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06436] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0321c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06438] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0321d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0643a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0321e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0643c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0321f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0643e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03220] =  I8a0037ad2845a3fbba9da380a8b8a576['h06440] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03221] =  I8a0037ad2845a3fbba9da380a8b8a576['h06442] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03222] =  I8a0037ad2845a3fbba9da380a8b8a576['h06444] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03223] =  I8a0037ad2845a3fbba9da380a8b8a576['h06446] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03224] =  I8a0037ad2845a3fbba9da380a8b8a576['h06448] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03225] =  I8a0037ad2845a3fbba9da380a8b8a576['h0644a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03226] =  I8a0037ad2845a3fbba9da380a8b8a576['h0644c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03227] =  I8a0037ad2845a3fbba9da380a8b8a576['h0644e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03228] =  I8a0037ad2845a3fbba9da380a8b8a576['h06450] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03229] =  I8a0037ad2845a3fbba9da380a8b8a576['h06452] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0322a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06454] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0322b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06456] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0322c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06458] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0322d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0645a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0322e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0645c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0322f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0645e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03230] =  I8a0037ad2845a3fbba9da380a8b8a576['h06460] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03231] =  I8a0037ad2845a3fbba9da380a8b8a576['h06462] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03232] =  I8a0037ad2845a3fbba9da380a8b8a576['h06464] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03233] =  I8a0037ad2845a3fbba9da380a8b8a576['h06466] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03234] =  I8a0037ad2845a3fbba9da380a8b8a576['h06468] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03235] =  I8a0037ad2845a3fbba9da380a8b8a576['h0646a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03236] =  I8a0037ad2845a3fbba9da380a8b8a576['h0646c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03237] =  I8a0037ad2845a3fbba9da380a8b8a576['h0646e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03238] =  I8a0037ad2845a3fbba9da380a8b8a576['h06470] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03239] =  I8a0037ad2845a3fbba9da380a8b8a576['h06472] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0323a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06474] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0323b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06476] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0323c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06478] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0323d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0647a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0323e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0647c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0323f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0647e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03240] =  I8a0037ad2845a3fbba9da380a8b8a576['h06480] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03241] =  I8a0037ad2845a3fbba9da380a8b8a576['h06482] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03242] =  I8a0037ad2845a3fbba9da380a8b8a576['h06484] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03243] =  I8a0037ad2845a3fbba9da380a8b8a576['h06486] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03244] =  I8a0037ad2845a3fbba9da380a8b8a576['h06488] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03245] =  I8a0037ad2845a3fbba9da380a8b8a576['h0648a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03246] =  I8a0037ad2845a3fbba9da380a8b8a576['h0648c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03247] =  I8a0037ad2845a3fbba9da380a8b8a576['h0648e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03248] =  I8a0037ad2845a3fbba9da380a8b8a576['h06490] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03249] =  I8a0037ad2845a3fbba9da380a8b8a576['h06492] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0324a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06494] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0324b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06496] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0324c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06498] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0324d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0649a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0324e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0649c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0324f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0649e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03250] =  I8a0037ad2845a3fbba9da380a8b8a576['h064a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03251] =  I8a0037ad2845a3fbba9da380a8b8a576['h064a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03252] =  I8a0037ad2845a3fbba9da380a8b8a576['h064a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03253] =  I8a0037ad2845a3fbba9da380a8b8a576['h064a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03254] =  I8a0037ad2845a3fbba9da380a8b8a576['h064a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03255] =  I8a0037ad2845a3fbba9da380a8b8a576['h064aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03256] =  I8a0037ad2845a3fbba9da380a8b8a576['h064ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03257] =  I8a0037ad2845a3fbba9da380a8b8a576['h064ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03258] =  I8a0037ad2845a3fbba9da380a8b8a576['h064b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03259] =  I8a0037ad2845a3fbba9da380a8b8a576['h064b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0325a] =  I8a0037ad2845a3fbba9da380a8b8a576['h064b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0325b] =  I8a0037ad2845a3fbba9da380a8b8a576['h064b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0325c] =  I8a0037ad2845a3fbba9da380a8b8a576['h064b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0325d] =  I8a0037ad2845a3fbba9da380a8b8a576['h064ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0325e] =  I8a0037ad2845a3fbba9da380a8b8a576['h064bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0325f] =  I8a0037ad2845a3fbba9da380a8b8a576['h064be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03260] =  I8a0037ad2845a3fbba9da380a8b8a576['h064c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03261] =  I8a0037ad2845a3fbba9da380a8b8a576['h064c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03262] =  I8a0037ad2845a3fbba9da380a8b8a576['h064c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03263] =  I8a0037ad2845a3fbba9da380a8b8a576['h064c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03264] =  I8a0037ad2845a3fbba9da380a8b8a576['h064c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03265] =  I8a0037ad2845a3fbba9da380a8b8a576['h064ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03266] =  I8a0037ad2845a3fbba9da380a8b8a576['h064cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03267] =  I8a0037ad2845a3fbba9da380a8b8a576['h064ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03268] =  I8a0037ad2845a3fbba9da380a8b8a576['h064d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03269] =  I8a0037ad2845a3fbba9da380a8b8a576['h064d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0326a] =  I8a0037ad2845a3fbba9da380a8b8a576['h064d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0326b] =  I8a0037ad2845a3fbba9da380a8b8a576['h064d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0326c] =  I8a0037ad2845a3fbba9da380a8b8a576['h064d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0326d] =  I8a0037ad2845a3fbba9da380a8b8a576['h064da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0326e] =  I8a0037ad2845a3fbba9da380a8b8a576['h064dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0326f] =  I8a0037ad2845a3fbba9da380a8b8a576['h064de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03270] =  I8a0037ad2845a3fbba9da380a8b8a576['h064e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03271] =  I8a0037ad2845a3fbba9da380a8b8a576['h064e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03272] =  I8a0037ad2845a3fbba9da380a8b8a576['h064e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03273] =  I8a0037ad2845a3fbba9da380a8b8a576['h064e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03274] =  I8a0037ad2845a3fbba9da380a8b8a576['h064e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03275] =  I8a0037ad2845a3fbba9da380a8b8a576['h064ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03276] =  I8a0037ad2845a3fbba9da380a8b8a576['h064ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03277] =  I8a0037ad2845a3fbba9da380a8b8a576['h064ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03278] =  I8a0037ad2845a3fbba9da380a8b8a576['h064f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03279] =  I8a0037ad2845a3fbba9da380a8b8a576['h064f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0327a] =  I8a0037ad2845a3fbba9da380a8b8a576['h064f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0327b] =  I8a0037ad2845a3fbba9da380a8b8a576['h064f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0327c] =  I8a0037ad2845a3fbba9da380a8b8a576['h064f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0327d] =  I8a0037ad2845a3fbba9da380a8b8a576['h064fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0327e] =  I8a0037ad2845a3fbba9da380a8b8a576['h064fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0327f] =  I8a0037ad2845a3fbba9da380a8b8a576['h064fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03280] =  I8a0037ad2845a3fbba9da380a8b8a576['h06500] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03281] =  I8a0037ad2845a3fbba9da380a8b8a576['h06502] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03282] =  I8a0037ad2845a3fbba9da380a8b8a576['h06504] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03283] =  I8a0037ad2845a3fbba9da380a8b8a576['h06506] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03284] =  I8a0037ad2845a3fbba9da380a8b8a576['h06508] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03285] =  I8a0037ad2845a3fbba9da380a8b8a576['h0650a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03286] =  I8a0037ad2845a3fbba9da380a8b8a576['h0650c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03287] =  I8a0037ad2845a3fbba9da380a8b8a576['h0650e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03288] =  I8a0037ad2845a3fbba9da380a8b8a576['h06510] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03289] =  I8a0037ad2845a3fbba9da380a8b8a576['h06512] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0328a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06514] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0328b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06516] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0328c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06518] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0328d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0651a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0328e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0651c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0328f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0651e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03290] =  I8a0037ad2845a3fbba9da380a8b8a576['h06520] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03291] =  I8a0037ad2845a3fbba9da380a8b8a576['h06522] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03292] =  I8a0037ad2845a3fbba9da380a8b8a576['h06524] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03293] =  I8a0037ad2845a3fbba9da380a8b8a576['h06526] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03294] =  I8a0037ad2845a3fbba9da380a8b8a576['h06528] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03295] =  I8a0037ad2845a3fbba9da380a8b8a576['h0652a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03296] =  I8a0037ad2845a3fbba9da380a8b8a576['h0652c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03297] =  I8a0037ad2845a3fbba9da380a8b8a576['h0652e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03298] =  I8a0037ad2845a3fbba9da380a8b8a576['h06530] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03299] =  I8a0037ad2845a3fbba9da380a8b8a576['h06532] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0329a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06534] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0329b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06536] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0329c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06538] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0329d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0653a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0329e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0653c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0329f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0653e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06540] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06542] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06544] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06546] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06548] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0654a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0654c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0654e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06550] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06552] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h06554] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h06556] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h06558] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0655a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0655c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032af] =  I8a0037ad2845a3fbba9da380a8b8a576['h0655e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06560] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06562] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06564] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06566] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06568] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0656a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0656c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0656e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06570] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06572] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h06574] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h06576] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h06578] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0657a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032be] =  I8a0037ad2845a3fbba9da380a8b8a576['h0657c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0657e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06580] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06582] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06584] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06586] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06588] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0658a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0658c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0658e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06590] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06592] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h06594] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h06596] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h06598] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0659a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0659c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0659e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h065a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h065a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h065a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h065a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h065a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h065aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h065ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h065ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h065b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h065b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032da] =  I8a0037ad2845a3fbba9da380a8b8a576['h065b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032db] =  I8a0037ad2845a3fbba9da380a8b8a576['h065b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h065b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h065ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032de] =  I8a0037ad2845a3fbba9da380a8b8a576['h065bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032df] =  I8a0037ad2845a3fbba9da380a8b8a576['h065be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h065c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h065c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h065c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h065c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h065c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h065ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h065cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h065ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h065d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h065d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h065d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h065d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h065d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h065da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h065dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h065de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h065e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h065e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h065e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h065e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h065e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h065ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h065ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h065ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h065f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h065f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h065f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h065f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h065f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h065fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h065fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h032ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h065fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03300] =  I8a0037ad2845a3fbba9da380a8b8a576['h06600] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03301] =  I8a0037ad2845a3fbba9da380a8b8a576['h06602] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03302] =  I8a0037ad2845a3fbba9da380a8b8a576['h06604] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03303] =  I8a0037ad2845a3fbba9da380a8b8a576['h06606] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03304] =  I8a0037ad2845a3fbba9da380a8b8a576['h06608] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03305] =  I8a0037ad2845a3fbba9da380a8b8a576['h0660a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03306] =  I8a0037ad2845a3fbba9da380a8b8a576['h0660c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03307] =  I8a0037ad2845a3fbba9da380a8b8a576['h0660e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03308] =  I8a0037ad2845a3fbba9da380a8b8a576['h06610] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03309] =  I8a0037ad2845a3fbba9da380a8b8a576['h06612] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0330a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06614] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0330b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06616] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0330c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06618] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0330d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0661a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0330e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0661c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0330f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0661e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03310] =  I8a0037ad2845a3fbba9da380a8b8a576['h06620] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03311] =  I8a0037ad2845a3fbba9da380a8b8a576['h06622] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03312] =  I8a0037ad2845a3fbba9da380a8b8a576['h06624] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03313] =  I8a0037ad2845a3fbba9da380a8b8a576['h06626] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03314] =  I8a0037ad2845a3fbba9da380a8b8a576['h06628] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03315] =  I8a0037ad2845a3fbba9da380a8b8a576['h0662a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03316] =  I8a0037ad2845a3fbba9da380a8b8a576['h0662c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03317] =  I8a0037ad2845a3fbba9da380a8b8a576['h0662e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03318] =  I8a0037ad2845a3fbba9da380a8b8a576['h06630] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03319] =  I8a0037ad2845a3fbba9da380a8b8a576['h06632] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0331a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06634] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0331b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06636] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0331c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06638] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0331d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0663a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0331e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0663c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0331f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0663e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03320] =  I8a0037ad2845a3fbba9da380a8b8a576['h06640] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03321] =  I8a0037ad2845a3fbba9da380a8b8a576['h06642] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03322] =  I8a0037ad2845a3fbba9da380a8b8a576['h06644] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03323] =  I8a0037ad2845a3fbba9da380a8b8a576['h06646] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03324] =  I8a0037ad2845a3fbba9da380a8b8a576['h06648] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03325] =  I8a0037ad2845a3fbba9da380a8b8a576['h0664a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03326] =  I8a0037ad2845a3fbba9da380a8b8a576['h0664c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03327] =  I8a0037ad2845a3fbba9da380a8b8a576['h0664e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03328] =  I8a0037ad2845a3fbba9da380a8b8a576['h06650] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03329] =  I8a0037ad2845a3fbba9da380a8b8a576['h06652] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0332a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06654] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0332b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06656] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0332c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06658] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0332d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0665a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0332e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0665c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0332f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0665e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03330] =  I8a0037ad2845a3fbba9da380a8b8a576['h06660] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03331] =  I8a0037ad2845a3fbba9da380a8b8a576['h06662] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03332] =  I8a0037ad2845a3fbba9da380a8b8a576['h06664] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03333] =  I8a0037ad2845a3fbba9da380a8b8a576['h06666] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03334] =  I8a0037ad2845a3fbba9da380a8b8a576['h06668] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03335] =  I8a0037ad2845a3fbba9da380a8b8a576['h0666a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03336] =  I8a0037ad2845a3fbba9da380a8b8a576['h0666c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03337] =  I8a0037ad2845a3fbba9da380a8b8a576['h0666e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03338] =  I8a0037ad2845a3fbba9da380a8b8a576['h06670] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03339] =  I8a0037ad2845a3fbba9da380a8b8a576['h06672] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0333a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06674] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0333b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06676] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0333c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06678] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0333d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0667a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0333e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0667c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0333f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0667e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03340] =  I8a0037ad2845a3fbba9da380a8b8a576['h06680] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03341] =  I8a0037ad2845a3fbba9da380a8b8a576['h06682] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03342] =  I8a0037ad2845a3fbba9da380a8b8a576['h06684] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03343] =  I8a0037ad2845a3fbba9da380a8b8a576['h06686] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03344] =  I8a0037ad2845a3fbba9da380a8b8a576['h06688] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03345] =  I8a0037ad2845a3fbba9da380a8b8a576['h0668a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03346] =  I8a0037ad2845a3fbba9da380a8b8a576['h0668c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03347] =  I8a0037ad2845a3fbba9da380a8b8a576['h0668e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03348] =  I8a0037ad2845a3fbba9da380a8b8a576['h06690] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03349] =  I8a0037ad2845a3fbba9da380a8b8a576['h06692] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0334a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06694] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0334b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06696] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0334c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06698] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0334d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0669a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0334e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0669c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0334f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0669e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03350] =  I8a0037ad2845a3fbba9da380a8b8a576['h066a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03351] =  I8a0037ad2845a3fbba9da380a8b8a576['h066a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03352] =  I8a0037ad2845a3fbba9da380a8b8a576['h066a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03353] =  I8a0037ad2845a3fbba9da380a8b8a576['h066a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03354] =  I8a0037ad2845a3fbba9da380a8b8a576['h066a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03355] =  I8a0037ad2845a3fbba9da380a8b8a576['h066aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03356] =  I8a0037ad2845a3fbba9da380a8b8a576['h066ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03357] =  I8a0037ad2845a3fbba9da380a8b8a576['h066ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03358] =  I8a0037ad2845a3fbba9da380a8b8a576['h066b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03359] =  I8a0037ad2845a3fbba9da380a8b8a576['h066b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0335a] =  I8a0037ad2845a3fbba9da380a8b8a576['h066b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0335b] =  I8a0037ad2845a3fbba9da380a8b8a576['h066b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0335c] =  I8a0037ad2845a3fbba9da380a8b8a576['h066b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0335d] =  I8a0037ad2845a3fbba9da380a8b8a576['h066ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0335e] =  I8a0037ad2845a3fbba9da380a8b8a576['h066bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0335f] =  I8a0037ad2845a3fbba9da380a8b8a576['h066be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03360] =  I8a0037ad2845a3fbba9da380a8b8a576['h066c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03361] =  I8a0037ad2845a3fbba9da380a8b8a576['h066c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03362] =  I8a0037ad2845a3fbba9da380a8b8a576['h066c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03363] =  I8a0037ad2845a3fbba9da380a8b8a576['h066c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03364] =  I8a0037ad2845a3fbba9da380a8b8a576['h066c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03365] =  I8a0037ad2845a3fbba9da380a8b8a576['h066ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03366] =  I8a0037ad2845a3fbba9da380a8b8a576['h066cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03367] =  I8a0037ad2845a3fbba9da380a8b8a576['h066ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03368] =  I8a0037ad2845a3fbba9da380a8b8a576['h066d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03369] =  I8a0037ad2845a3fbba9da380a8b8a576['h066d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0336a] =  I8a0037ad2845a3fbba9da380a8b8a576['h066d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0336b] =  I8a0037ad2845a3fbba9da380a8b8a576['h066d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0336c] =  I8a0037ad2845a3fbba9da380a8b8a576['h066d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0336d] =  I8a0037ad2845a3fbba9da380a8b8a576['h066da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0336e] =  I8a0037ad2845a3fbba9da380a8b8a576['h066dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0336f] =  I8a0037ad2845a3fbba9da380a8b8a576['h066de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03370] =  I8a0037ad2845a3fbba9da380a8b8a576['h066e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03371] =  I8a0037ad2845a3fbba9da380a8b8a576['h066e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03372] =  I8a0037ad2845a3fbba9da380a8b8a576['h066e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03373] =  I8a0037ad2845a3fbba9da380a8b8a576['h066e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03374] =  I8a0037ad2845a3fbba9da380a8b8a576['h066e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03375] =  I8a0037ad2845a3fbba9da380a8b8a576['h066ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03376] =  I8a0037ad2845a3fbba9da380a8b8a576['h066ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03377] =  I8a0037ad2845a3fbba9da380a8b8a576['h066ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03378] =  I8a0037ad2845a3fbba9da380a8b8a576['h066f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03379] =  I8a0037ad2845a3fbba9da380a8b8a576['h066f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0337a] =  I8a0037ad2845a3fbba9da380a8b8a576['h066f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0337b] =  I8a0037ad2845a3fbba9da380a8b8a576['h066f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0337c] =  I8a0037ad2845a3fbba9da380a8b8a576['h066f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0337d] =  I8a0037ad2845a3fbba9da380a8b8a576['h066fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0337e] =  I8a0037ad2845a3fbba9da380a8b8a576['h066fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0337f] =  I8a0037ad2845a3fbba9da380a8b8a576['h066fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03380] =  I8a0037ad2845a3fbba9da380a8b8a576['h06700] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03381] =  I8a0037ad2845a3fbba9da380a8b8a576['h06702] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03382] =  I8a0037ad2845a3fbba9da380a8b8a576['h06704] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03383] =  I8a0037ad2845a3fbba9da380a8b8a576['h06706] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03384] =  I8a0037ad2845a3fbba9da380a8b8a576['h06708] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03385] =  I8a0037ad2845a3fbba9da380a8b8a576['h0670a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03386] =  I8a0037ad2845a3fbba9da380a8b8a576['h0670c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03387] =  I8a0037ad2845a3fbba9da380a8b8a576['h0670e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03388] =  I8a0037ad2845a3fbba9da380a8b8a576['h06710] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03389] =  I8a0037ad2845a3fbba9da380a8b8a576['h06712] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0338a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06714] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0338b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06716] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0338c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06718] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0338d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0671a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0338e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0671c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0338f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0671e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03390] =  I8a0037ad2845a3fbba9da380a8b8a576['h06720] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03391] =  I8a0037ad2845a3fbba9da380a8b8a576['h06722] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03392] =  I8a0037ad2845a3fbba9da380a8b8a576['h06724] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03393] =  I8a0037ad2845a3fbba9da380a8b8a576['h06726] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03394] =  I8a0037ad2845a3fbba9da380a8b8a576['h06728] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03395] =  I8a0037ad2845a3fbba9da380a8b8a576['h0672a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03396] =  I8a0037ad2845a3fbba9da380a8b8a576['h0672c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03397] =  I8a0037ad2845a3fbba9da380a8b8a576['h0672e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03398] =  I8a0037ad2845a3fbba9da380a8b8a576['h06730] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03399] =  I8a0037ad2845a3fbba9da380a8b8a576['h06732] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0339a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06734] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0339b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06736] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0339c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06738] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0339d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0673a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0339e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0673c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0339f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0673e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06740] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06742] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06744] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06746] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06748] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0674a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0674c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0674e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06750] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06752] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h06754] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h06756] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h06758] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0675a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0675c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033af] =  I8a0037ad2845a3fbba9da380a8b8a576['h0675e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06760] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06762] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06764] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06766] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06768] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0676a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0676c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0676e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06770] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06772] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h06774] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h06776] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h06778] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0677a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033be] =  I8a0037ad2845a3fbba9da380a8b8a576['h0677c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0677e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06780] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06782] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06784] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06786] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06788] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0678a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0678c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0678e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06790] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06792] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h06794] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h06796] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h06798] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0679a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0679c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0679e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h067a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h067a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h067a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h067a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h067a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h067aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h067ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h067ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h067b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h067b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033da] =  I8a0037ad2845a3fbba9da380a8b8a576['h067b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033db] =  I8a0037ad2845a3fbba9da380a8b8a576['h067b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h067b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h067ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033de] =  I8a0037ad2845a3fbba9da380a8b8a576['h067bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033df] =  I8a0037ad2845a3fbba9da380a8b8a576['h067be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h067c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h067c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h067c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h067c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h067c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h067ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h067cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h067ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h067d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h067d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h067d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h067d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h067d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h067da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h067dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h067de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h067e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h067e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h067e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h067e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h067e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h067ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h067ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h067ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h067f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h067f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h067f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h067f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h067f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h067fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h067fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h033ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h067fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03400] =  I8a0037ad2845a3fbba9da380a8b8a576['h06800] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03401] =  I8a0037ad2845a3fbba9da380a8b8a576['h06802] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03402] =  I8a0037ad2845a3fbba9da380a8b8a576['h06804] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03403] =  I8a0037ad2845a3fbba9da380a8b8a576['h06806] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03404] =  I8a0037ad2845a3fbba9da380a8b8a576['h06808] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03405] =  I8a0037ad2845a3fbba9da380a8b8a576['h0680a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03406] =  I8a0037ad2845a3fbba9da380a8b8a576['h0680c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03407] =  I8a0037ad2845a3fbba9da380a8b8a576['h0680e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03408] =  I8a0037ad2845a3fbba9da380a8b8a576['h06810] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03409] =  I8a0037ad2845a3fbba9da380a8b8a576['h06812] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0340a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06814] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0340b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06816] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0340c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06818] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0340d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0681a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0340e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0681c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0340f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0681e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03410] =  I8a0037ad2845a3fbba9da380a8b8a576['h06820] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03411] =  I8a0037ad2845a3fbba9da380a8b8a576['h06822] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03412] =  I8a0037ad2845a3fbba9da380a8b8a576['h06824] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03413] =  I8a0037ad2845a3fbba9da380a8b8a576['h06826] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03414] =  I8a0037ad2845a3fbba9da380a8b8a576['h06828] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03415] =  I8a0037ad2845a3fbba9da380a8b8a576['h0682a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03416] =  I8a0037ad2845a3fbba9da380a8b8a576['h0682c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03417] =  I8a0037ad2845a3fbba9da380a8b8a576['h0682e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03418] =  I8a0037ad2845a3fbba9da380a8b8a576['h06830] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03419] =  I8a0037ad2845a3fbba9da380a8b8a576['h06832] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0341a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06834] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0341b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06836] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0341c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06838] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0341d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0683a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0341e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0683c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0341f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0683e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03420] =  I8a0037ad2845a3fbba9da380a8b8a576['h06840] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03421] =  I8a0037ad2845a3fbba9da380a8b8a576['h06842] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03422] =  I8a0037ad2845a3fbba9da380a8b8a576['h06844] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03423] =  I8a0037ad2845a3fbba9da380a8b8a576['h06846] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03424] =  I8a0037ad2845a3fbba9da380a8b8a576['h06848] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03425] =  I8a0037ad2845a3fbba9da380a8b8a576['h0684a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03426] =  I8a0037ad2845a3fbba9da380a8b8a576['h0684c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03427] =  I8a0037ad2845a3fbba9da380a8b8a576['h0684e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03428] =  I8a0037ad2845a3fbba9da380a8b8a576['h06850] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03429] =  I8a0037ad2845a3fbba9da380a8b8a576['h06852] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0342a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06854] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0342b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06856] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0342c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06858] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0342d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0685a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0342e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0685c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0342f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0685e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03430] =  I8a0037ad2845a3fbba9da380a8b8a576['h06860] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03431] =  I8a0037ad2845a3fbba9da380a8b8a576['h06862] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03432] =  I8a0037ad2845a3fbba9da380a8b8a576['h06864] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03433] =  I8a0037ad2845a3fbba9da380a8b8a576['h06866] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03434] =  I8a0037ad2845a3fbba9da380a8b8a576['h06868] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03435] =  I8a0037ad2845a3fbba9da380a8b8a576['h0686a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03436] =  I8a0037ad2845a3fbba9da380a8b8a576['h0686c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03437] =  I8a0037ad2845a3fbba9da380a8b8a576['h0686e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03438] =  I8a0037ad2845a3fbba9da380a8b8a576['h06870] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03439] =  I8a0037ad2845a3fbba9da380a8b8a576['h06872] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0343a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06874] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0343b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06876] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0343c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06878] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0343d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0687a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0343e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0687c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0343f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0687e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03440] =  I8a0037ad2845a3fbba9da380a8b8a576['h06880] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03441] =  I8a0037ad2845a3fbba9da380a8b8a576['h06882] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03442] =  I8a0037ad2845a3fbba9da380a8b8a576['h06884] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03443] =  I8a0037ad2845a3fbba9da380a8b8a576['h06886] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03444] =  I8a0037ad2845a3fbba9da380a8b8a576['h06888] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03445] =  I8a0037ad2845a3fbba9da380a8b8a576['h0688a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03446] =  I8a0037ad2845a3fbba9da380a8b8a576['h0688c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03447] =  I8a0037ad2845a3fbba9da380a8b8a576['h0688e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03448] =  I8a0037ad2845a3fbba9da380a8b8a576['h06890] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03449] =  I8a0037ad2845a3fbba9da380a8b8a576['h06892] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0344a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06894] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0344b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06896] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0344c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06898] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0344d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0689a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0344e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0689c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0344f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0689e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03450] =  I8a0037ad2845a3fbba9da380a8b8a576['h068a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03451] =  I8a0037ad2845a3fbba9da380a8b8a576['h068a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03452] =  I8a0037ad2845a3fbba9da380a8b8a576['h068a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03453] =  I8a0037ad2845a3fbba9da380a8b8a576['h068a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03454] =  I8a0037ad2845a3fbba9da380a8b8a576['h068a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03455] =  I8a0037ad2845a3fbba9da380a8b8a576['h068aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03456] =  I8a0037ad2845a3fbba9da380a8b8a576['h068ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03457] =  I8a0037ad2845a3fbba9da380a8b8a576['h068ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03458] =  I8a0037ad2845a3fbba9da380a8b8a576['h068b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03459] =  I8a0037ad2845a3fbba9da380a8b8a576['h068b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0345a] =  I8a0037ad2845a3fbba9da380a8b8a576['h068b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0345b] =  I8a0037ad2845a3fbba9da380a8b8a576['h068b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0345c] =  I8a0037ad2845a3fbba9da380a8b8a576['h068b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0345d] =  I8a0037ad2845a3fbba9da380a8b8a576['h068ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0345e] =  I8a0037ad2845a3fbba9da380a8b8a576['h068bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0345f] =  I8a0037ad2845a3fbba9da380a8b8a576['h068be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03460] =  I8a0037ad2845a3fbba9da380a8b8a576['h068c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03461] =  I8a0037ad2845a3fbba9da380a8b8a576['h068c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03462] =  I8a0037ad2845a3fbba9da380a8b8a576['h068c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03463] =  I8a0037ad2845a3fbba9da380a8b8a576['h068c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03464] =  I8a0037ad2845a3fbba9da380a8b8a576['h068c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03465] =  I8a0037ad2845a3fbba9da380a8b8a576['h068ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03466] =  I8a0037ad2845a3fbba9da380a8b8a576['h068cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03467] =  I8a0037ad2845a3fbba9da380a8b8a576['h068ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03468] =  I8a0037ad2845a3fbba9da380a8b8a576['h068d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03469] =  I8a0037ad2845a3fbba9da380a8b8a576['h068d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0346a] =  I8a0037ad2845a3fbba9da380a8b8a576['h068d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0346b] =  I8a0037ad2845a3fbba9da380a8b8a576['h068d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0346c] =  I8a0037ad2845a3fbba9da380a8b8a576['h068d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0346d] =  I8a0037ad2845a3fbba9da380a8b8a576['h068da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0346e] =  I8a0037ad2845a3fbba9da380a8b8a576['h068dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0346f] =  I8a0037ad2845a3fbba9da380a8b8a576['h068de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03470] =  I8a0037ad2845a3fbba9da380a8b8a576['h068e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03471] =  I8a0037ad2845a3fbba9da380a8b8a576['h068e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03472] =  I8a0037ad2845a3fbba9da380a8b8a576['h068e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03473] =  I8a0037ad2845a3fbba9da380a8b8a576['h068e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03474] =  I8a0037ad2845a3fbba9da380a8b8a576['h068e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03475] =  I8a0037ad2845a3fbba9da380a8b8a576['h068ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03476] =  I8a0037ad2845a3fbba9da380a8b8a576['h068ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03477] =  I8a0037ad2845a3fbba9da380a8b8a576['h068ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03478] =  I8a0037ad2845a3fbba9da380a8b8a576['h068f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03479] =  I8a0037ad2845a3fbba9da380a8b8a576['h068f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0347a] =  I8a0037ad2845a3fbba9da380a8b8a576['h068f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0347b] =  I8a0037ad2845a3fbba9da380a8b8a576['h068f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0347c] =  I8a0037ad2845a3fbba9da380a8b8a576['h068f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0347d] =  I8a0037ad2845a3fbba9da380a8b8a576['h068fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0347e] =  I8a0037ad2845a3fbba9da380a8b8a576['h068fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0347f] =  I8a0037ad2845a3fbba9da380a8b8a576['h068fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03480] =  I8a0037ad2845a3fbba9da380a8b8a576['h06900] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03481] =  I8a0037ad2845a3fbba9da380a8b8a576['h06902] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03482] =  I8a0037ad2845a3fbba9da380a8b8a576['h06904] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03483] =  I8a0037ad2845a3fbba9da380a8b8a576['h06906] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03484] =  I8a0037ad2845a3fbba9da380a8b8a576['h06908] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03485] =  I8a0037ad2845a3fbba9da380a8b8a576['h0690a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03486] =  I8a0037ad2845a3fbba9da380a8b8a576['h0690c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03487] =  I8a0037ad2845a3fbba9da380a8b8a576['h0690e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03488] =  I8a0037ad2845a3fbba9da380a8b8a576['h06910] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03489] =  I8a0037ad2845a3fbba9da380a8b8a576['h06912] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0348a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06914] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0348b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06916] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0348c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06918] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0348d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0691a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0348e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0691c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0348f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0691e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03490] =  I8a0037ad2845a3fbba9da380a8b8a576['h06920] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03491] =  I8a0037ad2845a3fbba9da380a8b8a576['h06922] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03492] =  I8a0037ad2845a3fbba9da380a8b8a576['h06924] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03493] =  I8a0037ad2845a3fbba9da380a8b8a576['h06926] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03494] =  I8a0037ad2845a3fbba9da380a8b8a576['h06928] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03495] =  I8a0037ad2845a3fbba9da380a8b8a576['h0692a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03496] =  I8a0037ad2845a3fbba9da380a8b8a576['h0692c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03497] =  I8a0037ad2845a3fbba9da380a8b8a576['h0692e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03498] =  I8a0037ad2845a3fbba9da380a8b8a576['h06930] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03499] =  I8a0037ad2845a3fbba9da380a8b8a576['h06932] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0349a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06934] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0349b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06936] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0349c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06938] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0349d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0693a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0349e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0693c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0349f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0693e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06940] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06942] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06944] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06946] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06948] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0694a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0694c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0694e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06950] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06952] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h06954] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h06956] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h06958] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0695a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0695c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034af] =  I8a0037ad2845a3fbba9da380a8b8a576['h0695e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06960] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06962] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06964] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06966] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06968] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0696a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0696c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0696e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06970] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06972] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h06974] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h06976] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h06978] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0697a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034be] =  I8a0037ad2845a3fbba9da380a8b8a576['h0697c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0697e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06980] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06982] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06984] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06986] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06988] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0698a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0698c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0698e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06990] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06992] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h06994] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h06996] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h06998] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0699a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0699c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0699e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h069a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h069a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h069a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h069a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h069a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h069aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h069ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h069ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h069b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h069b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034da] =  I8a0037ad2845a3fbba9da380a8b8a576['h069b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034db] =  I8a0037ad2845a3fbba9da380a8b8a576['h069b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h069b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h069ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034de] =  I8a0037ad2845a3fbba9da380a8b8a576['h069bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034df] =  I8a0037ad2845a3fbba9da380a8b8a576['h069be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h069c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h069c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h069c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h069c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h069c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h069ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h069cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h069ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h069d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h069d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h069d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h069d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h069d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h069da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h069dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h069de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h069e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h069e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h069e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h069e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h069e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h069ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h069ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h069ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h069f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h069f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h069f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h069f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h069f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h069fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h069fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h034ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h069fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03500] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03501] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03502] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03503] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03504] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03505] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03506] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03507] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03508] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03509] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0350a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0350b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0350c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0350d] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0350e] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0350f] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03510] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03511] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03512] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03513] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03514] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03515] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03516] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03517] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03518] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03519] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0351a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0351b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0351c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0351d] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0351e] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0351f] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03520] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03521] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03522] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03523] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03524] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03525] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03526] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03527] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03528] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03529] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0352a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0352b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0352c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0352d] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0352e] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0352f] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03530] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03531] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03532] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03533] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03534] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03535] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03536] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03537] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03538] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03539] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0353a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0353b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0353c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0353d] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0353e] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0353f] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03540] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03541] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03542] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03543] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03544] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03545] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03546] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03547] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03548] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03549] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0354a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0354b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0354c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0354d] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0354e] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0354f] =  I8a0037ad2845a3fbba9da380a8b8a576['h06a9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03550] =  I8a0037ad2845a3fbba9da380a8b8a576['h06aa0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03551] =  I8a0037ad2845a3fbba9da380a8b8a576['h06aa2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03552] =  I8a0037ad2845a3fbba9da380a8b8a576['h06aa4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03553] =  I8a0037ad2845a3fbba9da380a8b8a576['h06aa6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03554] =  I8a0037ad2845a3fbba9da380a8b8a576['h06aa8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03555] =  I8a0037ad2845a3fbba9da380a8b8a576['h06aaa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03556] =  I8a0037ad2845a3fbba9da380a8b8a576['h06aac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03557] =  I8a0037ad2845a3fbba9da380a8b8a576['h06aae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03558] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ab0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03559] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ab2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0355a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ab4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0355b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ab6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0355c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ab8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0355d] =  I8a0037ad2845a3fbba9da380a8b8a576['h06aba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0355e] =  I8a0037ad2845a3fbba9da380a8b8a576['h06abc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0355f] =  I8a0037ad2845a3fbba9da380a8b8a576['h06abe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03560] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ac0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03561] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ac2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03562] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ac4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03563] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ac6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03564] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ac8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03565] =  I8a0037ad2845a3fbba9da380a8b8a576['h06aca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03566] =  I8a0037ad2845a3fbba9da380a8b8a576['h06acc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03567] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ace] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03568] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ad0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03569] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ad2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0356a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ad4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0356b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ad6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0356c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ad8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0356d] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ada] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0356e] =  I8a0037ad2845a3fbba9da380a8b8a576['h06adc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0356f] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ade] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03570] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ae0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03571] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ae2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03572] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ae4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03573] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ae6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03574] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ae8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03575] =  I8a0037ad2845a3fbba9da380a8b8a576['h06aea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03576] =  I8a0037ad2845a3fbba9da380a8b8a576['h06aec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03577] =  I8a0037ad2845a3fbba9da380a8b8a576['h06aee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03578] =  I8a0037ad2845a3fbba9da380a8b8a576['h06af0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03579] =  I8a0037ad2845a3fbba9da380a8b8a576['h06af2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0357a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06af4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0357b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06af6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0357c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06af8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0357d] =  I8a0037ad2845a3fbba9da380a8b8a576['h06afa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0357e] =  I8a0037ad2845a3fbba9da380a8b8a576['h06afc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0357f] =  I8a0037ad2845a3fbba9da380a8b8a576['h06afe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03580] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03581] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03582] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03583] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03584] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03585] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03586] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03587] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03588] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03589] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0358a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0358b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0358c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0358d] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0358e] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0358f] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03590] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03591] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03592] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03593] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03594] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03595] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03596] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03597] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03598] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03599] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0359a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0359b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0359c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0359d] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0359e] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0359f] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035af] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035be] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h06b9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ba0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ba2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ba4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ba6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ba8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h06baa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035da] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035db] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035de] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035df] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bcc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bdc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06be0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06be2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06be4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06be6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06be8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bf0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bf2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bf4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bf6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bf8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bfa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bfc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h035ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h06bfe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03600] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03601] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03602] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03603] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03604] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03605] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03606] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03607] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03608] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03609] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0360a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0360b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0360c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0360d] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0360e] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0360f] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03610] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03611] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03612] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03613] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03614] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03615] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03616] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03617] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03618] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03619] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0361a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0361b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0361c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0361d] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0361e] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0361f] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03620] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03621] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03622] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03623] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03624] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03625] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03626] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03627] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03628] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03629] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0362a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0362b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0362c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0362d] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0362e] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0362f] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03630] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03631] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03632] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03633] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03634] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03635] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03636] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03637] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03638] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03639] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0363a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0363b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0363c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0363d] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0363e] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0363f] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03640] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03641] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03642] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03643] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03644] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03645] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03646] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03647] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03648] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03649] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0364a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0364b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0364c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0364d] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0364e] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0364f] =  I8a0037ad2845a3fbba9da380a8b8a576['h06c9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03650] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ca0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03651] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ca2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03652] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ca4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03653] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ca6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03654] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ca8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03655] =  I8a0037ad2845a3fbba9da380a8b8a576['h06caa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03656] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03657] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03658] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03659] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0365a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0365b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0365c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0365d] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0365e] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0365f] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03660] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03661] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03662] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03663] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03664] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03665] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03666] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ccc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03667] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03668] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03669] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0366a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0366b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0366c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0366d] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0366e] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cdc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0366f] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03670] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ce0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03671] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ce2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03672] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ce4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03673] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ce6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03674] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ce8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03675] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03676] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03677] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03678] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cf0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03679] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cf2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0367a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cf4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0367b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cf6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0367c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cf8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0367d] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cfa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0367e] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cfc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0367f] =  I8a0037ad2845a3fbba9da380a8b8a576['h06cfe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03680] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03681] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03682] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03683] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03684] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03685] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03686] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03687] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03688] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03689] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0368a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0368b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0368c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0368d] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0368e] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0368f] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03690] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03691] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03692] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03693] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03694] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03695] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03696] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03697] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03698] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03699] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0369a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0369b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0369c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0369d] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0369e] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0369f] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036af] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036be] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h06d9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06da0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06da2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06da4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06da6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06da8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h06daa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h06dac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h06dae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06db0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06db2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036da] =  I8a0037ad2845a3fbba9da380a8b8a576['h06db4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036db] =  I8a0037ad2845a3fbba9da380a8b8a576['h06db6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h06db8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h06dba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036de] =  I8a0037ad2845a3fbba9da380a8b8a576['h06dbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036df] =  I8a0037ad2845a3fbba9da380a8b8a576['h06dbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06dc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06dc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06dc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06dc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06dc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h06dca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h06dcc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h06dce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06dd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06dd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h06dd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h06dd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h06dd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h06dda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ddc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h06dde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06de0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06de2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06de4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06de6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06de8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h06dea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h06dec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h06dee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06df0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06df2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h06df4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h06df6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h06df8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h06dfa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h06dfc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h036ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h06dfe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03700] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03701] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03702] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03703] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03704] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03705] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03706] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03707] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03708] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03709] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0370a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0370b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0370c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0370d] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0370e] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0370f] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03710] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03711] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03712] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03713] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03714] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03715] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03716] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03717] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03718] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03719] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0371a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0371b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0371c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0371d] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0371e] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0371f] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03720] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03721] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03722] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03723] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03724] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03725] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03726] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03727] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03728] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03729] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0372a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0372b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0372c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0372d] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0372e] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0372f] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03730] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03731] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03732] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03733] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03734] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03735] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03736] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03737] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03738] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03739] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0373a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0373b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0373c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0373d] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0373e] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0373f] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03740] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03741] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03742] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03743] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03744] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03745] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03746] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03747] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03748] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03749] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0374a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0374b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0374c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0374d] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0374e] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0374f] =  I8a0037ad2845a3fbba9da380a8b8a576['h06e9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03750] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ea0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03751] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ea2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03752] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ea4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03753] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ea6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03754] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ea8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03755] =  I8a0037ad2845a3fbba9da380a8b8a576['h06eaa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03756] =  I8a0037ad2845a3fbba9da380a8b8a576['h06eac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03757] =  I8a0037ad2845a3fbba9da380a8b8a576['h06eae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03758] =  I8a0037ad2845a3fbba9da380a8b8a576['h06eb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03759] =  I8a0037ad2845a3fbba9da380a8b8a576['h06eb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0375a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06eb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0375b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06eb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0375c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06eb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0375d] =  I8a0037ad2845a3fbba9da380a8b8a576['h06eba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0375e] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ebc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0375f] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ebe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03760] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ec0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03761] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ec2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03762] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ec4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03763] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ec6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03764] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ec8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03765] =  I8a0037ad2845a3fbba9da380a8b8a576['h06eca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03766] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ecc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03767] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ece] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03768] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ed0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03769] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ed2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0376a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ed4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0376b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ed6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0376c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ed8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0376d] =  I8a0037ad2845a3fbba9da380a8b8a576['h06eda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0376e] =  I8a0037ad2845a3fbba9da380a8b8a576['h06edc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0376f] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ede] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03770] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ee0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03771] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ee2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03772] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ee4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03773] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ee6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03774] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ee8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03775] =  I8a0037ad2845a3fbba9da380a8b8a576['h06eea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03776] =  I8a0037ad2845a3fbba9da380a8b8a576['h06eec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03777] =  I8a0037ad2845a3fbba9da380a8b8a576['h06eee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03778] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ef0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03779] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ef2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0377a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ef4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0377b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ef6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0377c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ef8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0377d] =  I8a0037ad2845a3fbba9da380a8b8a576['h06efa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0377e] =  I8a0037ad2845a3fbba9da380a8b8a576['h06efc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0377f] =  I8a0037ad2845a3fbba9da380a8b8a576['h06efe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03780] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03781] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03782] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03783] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03784] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03785] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03786] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03787] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03788] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03789] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0378a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0378b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0378c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0378d] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0378e] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0378f] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03790] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03791] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03792] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03793] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03794] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03795] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03796] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03797] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03798] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03799] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0379a] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0379b] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0379c] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0379d] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0379e] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0379f] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037af] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037be] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h06f9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fa0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fa2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fa4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fa6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fa8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h06faa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037da] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037db] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037de] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037df] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fcc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fdc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fe0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fe2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fe4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fe6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fe8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h06fee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ff0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ff2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ff4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ff6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ff8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ffa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ffc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h037ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h06ffe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03800] =  I8a0037ad2845a3fbba9da380a8b8a576['h07000] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03801] =  I8a0037ad2845a3fbba9da380a8b8a576['h07002] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03802] =  I8a0037ad2845a3fbba9da380a8b8a576['h07004] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03803] =  I8a0037ad2845a3fbba9da380a8b8a576['h07006] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03804] =  I8a0037ad2845a3fbba9da380a8b8a576['h07008] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03805] =  I8a0037ad2845a3fbba9da380a8b8a576['h0700a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03806] =  I8a0037ad2845a3fbba9da380a8b8a576['h0700c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03807] =  I8a0037ad2845a3fbba9da380a8b8a576['h0700e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03808] =  I8a0037ad2845a3fbba9da380a8b8a576['h07010] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03809] =  I8a0037ad2845a3fbba9da380a8b8a576['h07012] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0380a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07014] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0380b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07016] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0380c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07018] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0380d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0701a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0380e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0701c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0380f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0701e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03810] =  I8a0037ad2845a3fbba9da380a8b8a576['h07020] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03811] =  I8a0037ad2845a3fbba9da380a8b8a576['h07022] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03812] =  I8a0037ad2845a3fbba9da380a8b8a576['h07024] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03813] =  I8a0037ad2845a3fbba9da380a8b8a576['h07026] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03814] =  I8a0037ad2845a3fbba9da380a8b8a576['h07028] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03815] =  I8a0037ad2845a3fbba9da380a8b8a576['h0702a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03816] =  I8a0037ad2845a3fbba9da380a8b8a576['h0702c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03817] =  I8a0037ad2845a3fbba9da380a8b8a576['h0702e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03818] =  I8a0037ad2845a3fbba9da380a8b8a576['h07030] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03819] =  I8a0037ad2845a3fbba9da380a8b8a576['h07032] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0381a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07034] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0381b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07036] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0381c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07038] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0381d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0703a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0381e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0703c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0381f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0703e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03820] =  I8a0037ad2845a3fbba9da380a8b8a576['h07040] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03821] =  I8a0037ad2845a3fbba9da380a8b8a576['h07042] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03822] =  I8a0037ad2845a3fbba9da380a8b8a576['h07044] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03823] =  I8a0037ad2845a3fbba9da380a8b8a576['h07046] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03824] =  I8a0037ad2845a3fbba9da380a8b8a576['h07048] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03825] =  I8a0037ad2845a3fbba9da380a8b8a576['h0704a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03826] =  I8a0037ad2845a3fbba9da380a8b8a576['h0704c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03827] =  I8a0037ad2845a3fbba9da380a8b8a576['h0704e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03828] =  I8a0037ad2845a3fbba9da380a8b8a576['h07050] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03829] =  I8a0037ad2845a3fbba9da380a8b8a576['h07052] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0382a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07054] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0382b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07056] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0382c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07058] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0382d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0705a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0382e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0705c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0382f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0705e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03830] =  I8a0037ad2845a3fbba9da380a8b8a576['h07060] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03831] =  I8a0037ad2845a3fbba9da380a8b8a576['h07062] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03832] =  I8a0037ad2845a3fbba9da380a8b8a576['h07064] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03833] =  I8a0037ad2845a3fbba9da380a8b8a576['h07066] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03834] =  I8a0037ad2845a3fbba9da380a8b8a576['h07068] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03835] =  I8a0037ad2845a3fbba9da380a8b8a576['h0706a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03836] =  I8a0037ad2845a3fbba9da380a8b8a576['h0706c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03837] =  I8a0037ad2845a3fbba9da380a8b8a576['h0706e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03838] =  I8a0037ad2845a3fbba9da380a8b8a576['h07070] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03839] =  I8a0037ad2845a3fbba9da380a8b8a576['h07072] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0383a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07074] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0383b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07076] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0383c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07078] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0383d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0707a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0383e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0707c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0383f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0707e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03840] =  I8a0037ad2845a3fbba9da380a8b8a576['h07080] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03841] =  I8a0037ad2845a3fbba9da380a8b8a576['h07082] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03842] =  I8a0037ad2845a3fbba9da380a8b8a576['h07084] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03843] =  I8a0037ad2845a3fbba9da380a8b8a576['h07086] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03844] =  I8a0037ad2845a3fbba9da380a8b8a576['h07088] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03845] =  I8a0037ad2845a3fbba9da380a8b8a576['h0708a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03846] =  I8a0037ad2845a3fbba9da380a8b8a576['h0708c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03847] =  I8a0037ad2845a3fbba9da380a8b8a576['h0708e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03848] =  I8a0037ad2845a3fbba9da380a8b8a576['h07090] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03849] =  I8a0037ad2845a3fbba9da380a8b8a576['h07092] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0384a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07094] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0384b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07096] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0384c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07098] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0384d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0709a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0384e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0709c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0384f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0709e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03850] =  I8a0037ad2845a3fbba9da380a8b8a576['h070a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03851] =  I8a0037ad2845a3fbba9da380a8b8a576['h070a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03852] =  I8a0037ad2845a3fbba9da380a8b8a576['h070a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03853] =  I8a0037ad2845a3fbba9da380a8b8a576['h070a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03854] =  I8a0037ad2845a3fbba9da380a8b8a576['h070a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03855] =  I8a0037ad2845a3fbba9da380a8b8a576['h070aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03856] =  I8a0037ad2845a3fbba9da380a8b8a576['h070ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03857] =  I8a0037ad2845a3fbba9da380a8b8a576['h070ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03858] =  I8a0037ad2845a3fbba9da380a8b8a576['h070b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03859] =  I8a0037ad2845a3fbba9da380a8b8a576['h070b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0385a] =  I8a0037ad2845a3fbba9da380a8b8a576['h070b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0385b] =  I8a0037ad2845a3fbba9da380a8b8a576['h070b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0385c] =  I8a0037ad2845a3fbba9da380a8b8a576['h070b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0385d] =  I8a0037ad2845a3fbba9da380a8b8a576['h070ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0385e] =  I8a0037ad2845a3fbba9da380a8b8a576['h070bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0385f] =  I8a0037ad2845a3fbba9da380a8b8a576['h070be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03860] =  I8a0037ad2845a3fbba9da380a8b8a576['h070c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03861] =  I8a0037ad2845a3fbba9da380a8b8a576['h070c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03862] =  I8a0037ad2845a3fbba9da380a8b8a576['h070c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03863] =  I8a0037ad2845a3fbba9da380a8b8a576['h070c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03864] =  I8a0037ad2845a3fbba9da380a8b8a576['h070c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03865] =  I8a0037ad2845a3fbba9da380a8b8a576['h070ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03866] =  I8a0037ad2845a3fbba9da380a8b8a576['h070cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03867] =  I8a0037ad2845a3fbba9da380a8b8a576['h070ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03868] =  I8a0037ad2845a3fbba9da380a8b8a576['h070d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03869] =  I8a0037ad2845a3fbba9da380a8b8a576['h070d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0386a] =  I8a0037ad2845a3fbba9da380a8b8a576['h070d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0386b] =  I8a0037ad2845a3fbba9da380a8b8a576['h070d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0386c] =  I8a0037ad2845a3fbba9da380a8b8a576['h070d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0386d] =  I8a0037ad2845a3fbba9da380a8b8a576['h070da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0386e] =  I8a0037ad2845a3fbba9da380a8b8a576['h070dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0386f] =  I8a0037ad2845a3fbba9da380a8b8a576['h070de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03870] =  I8a0037ad2845a3fbba9da380a8b8a576['h070e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03871] =  I8a0037ad2845a3fbba9da380a8b8a576['h070e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03872] =  I8a0037ad2845a3fbba9da380a8b8a576['h070e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03873] =  I8a0037ad2845a3fbba9da380a8b8a576['h070e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03874] =  I8a0037ad2845a3fbba9da380a8b8a576['h070e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03875] =  I8a0037ad2845a3fbba9da380a8b8a576['h070ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03876] =  I8a0037ad2845a3fbba9da380a8b8a576['h070ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03877] =  I8a0037ad2845a3fbba9da380a8b8a576['h070ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03878] =  I8a0037ad2845a3fbba9da380a8b8a576['h070f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03879] =  I8a0037ad2845a3fbba9da380a8b8a576['h070f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0387a] =  I8a0037ad2845a3fbba9da380a8b8a576['h070f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0387b] =  I8a0037ad2845a3fbba9da380a8b8a576['h070f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0387c] =  I8a0037ad2845a3fbba9da380a8b8a576['h070f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0387d] =  I8a0037ad2845a3fbba9da380a8b8a576['h070fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0387e] =  I8a0037ad2845a3fbba9da380a8b8a576['h070fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0387f] =  I8a0037ad2845a3fbba9da380a8b8a576['h070fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03880] =  I8a0037ad2845a3fbba9da380a8b8a576['h07100] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03881] =  I8a0037ad2845a3fbba9da380a8b8a576['h07102] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03882] =  I8a0037ad2845a3fbba9da380a8b8a576['h07104] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03883] =  I8a0037ad2845a3fbba9da380a8b8a576['h07106] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03884] =  I8a0037ad2845a3fbba9da380a8b8a576['h07108] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03885] =  I8a0037ad2845a3fbba9da380a8b8a576['h0710a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03886] =  I8a0037ad2845a3fbba9da380a8b8a576['h0710c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03887] =  I8a0037ad2845a3fbba9da380a8b8a576['h0710e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03888] =  I8a0037ad2845a3fbba9da380a8b8a576['h07110] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03889] =  I8a0037ad2845a3fbba9da380a8b8a576['h07112] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0388a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07114] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0388b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07116] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0388c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07118] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0388d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0711a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0388e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0711c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0388f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0711e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03890] =  I8a0037ad2845a3fbba9da380a8b8a576['h07120] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03891] =  I8a0037ad2845a3fbba9da380a8b8a576['h07122] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03892] =  I8a0037ad2845a3fbba9da380a8b8a576['h07124] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03893] =  I8a0037ad2845a3fbba9da380a8b8a576['h07126] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03894] =  I8a0037ad2845a3fbba9da380a8b8a576['h07128] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03895] =  I8a0037ad2845a3fbba9da380a8b8a576['h0712a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03896] =  I8a0037ad2845a3fbba9da380a8b8a576['h0712c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03897] =  I8a0037ad2845a3fbba9da380a8b8a576['h0712e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03898] =  I8a0037ad2845a3fbba9da380a8b8a576['h07130] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03899] =  I8a0037ad2845a3fbba9da380a8b8a576['h07132] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0389a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07134] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0389b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07136] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0389c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07138] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0389d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0713a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0389e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0713c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0389f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0713e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07140] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07142] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07144] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07146] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07148] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0714a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0714c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0714e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07150] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07152] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h07154] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h07156] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h07158] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0715a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0715c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038af] =  I8a0037ad2845a3fbba9da380a8b8a576['h0715e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07160] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07162] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07164] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07166] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07168] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0716a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0716c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0716e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07170] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07172] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h07174] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h07176] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h07178] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0717a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038be] =  I8a0037ad2845a3fbba9da380a8b8a576['h0717c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0717e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07180] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07182] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07184] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07186] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07188] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0718a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0718c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0718e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07190] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07192] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h07194] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h07196] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h07198] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0719a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0719c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0719e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h071a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h071a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h071a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h071a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h071a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h071aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h071ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h071ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h071b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h071b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038da] =  I8a0037ad2845a3fbba9da380a8b8a576['h071b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038db] =  I8a0037ad2845a3fbba9da380a8b8a576['h071b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h071b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h071ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038de] =  I8a0037ad2845a3fbba9da380a8b8a576['h071bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038df] =  I8a0037ad2845a3fbba9da380a8b8a576['h071be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h071c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h071c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h071c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h071c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h071c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h071ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h071cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h071ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h071d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h071d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h071d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h071d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h071d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h071da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h071dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h071de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h071e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h071e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h071e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h071e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h071e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h071ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h071ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h071ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h071f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h071f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h071f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h071f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h071f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h071fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h071fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h038ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h071fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03900] =  I8a0037ad2845a3fbba9da380a8b8a576['h07200] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03901] =  I8a0037ad2845a3fbba9da380a8b8a576['h07202] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03902] =  I8a0037ad2845a3fbba9da380a8b8a576['h07204] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03903] =  I8a0037ad2845a3fbba9da380a8b8a576['h07206] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03904] =  I8a0037ad2845a3fbba9da380a8b8a576['h07208] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03905] =  I8a0037ad2845a3fbba9da380a8b8a576['h0720a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03906] =  I8a0037ad2845a3fbba9da380a8b8a576['h0720c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03907] =  I8a0037ad2845a3fbba9da380a8b8a576['h0720e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03908] =  I8a0037ad2845a3fbba9da380a8b8a576['h07210] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03909] =  I8a0037ad2845a3fbba9da380a8b8a576['h07212] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0390a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07214] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0390b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07216] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0390c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07218] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0390d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0721a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0390e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0721c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0390f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0721e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03910] =  I8a0037ad2845a3fbba9da380a8b8a576['h07220] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03911] =  I8a0037ad2845a3fbba9da380a8b8a576['h07222] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03912] =  I8a0037ad2845a3fbba9da380a8b8a576['h07224] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03913] =  I8a0037ad2845a3fbba9da380a8b8a576['h07226] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03914] =  I8a0037ad2845a3fbba9da380a8b8a576['h07228] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03915] =  I8a0037ad2845a3fbba9da380a8b8a576['h0722a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03916] =  I8a0037ad2845a3fbba9da380a8b8a576['h0722c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03917] =  I8a0037ad2845a3fbba9da380a8b8a576['h0722e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03918] =  I8a0037ad2845a3fbba9da380a8b8a576['h07230] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03919] =  I8a0037ad2845a3fbba9da380a8b8a576['h07232] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0391a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07234] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0391b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07236] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0391c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07238] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0391d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0723a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0391e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0723c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0391f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0723e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03920] =  I8a0037ad2845a3fbba9da380a8b8a576['h07240] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03921] =  I8a0037ad2845a3fbba9da380a8b8a576['h07242] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03922] =  I8a0037ad2845a3fbba9da380a8b8a576['h07244] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03923] =  I8a0037ad2845a3fbba9da380a8b8a576['h07246] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03924] =  I8a0037ad2845a3fbba9da380a8b8a576['h07248] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03925] =  I8a0037ad2845a3fbba9da380a8b8a576['h0724a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03926] =  I8a0037ad2845a3fbba9da380a8b8a576['h0724c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03927] =  I8a0037ad2845a3fbba9da380a8b8a576['h0724e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03928] =  I8a0037ad2845a3fbba9da380a8b8a576['h07250] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03929] =  I8a0037ad2845a3fbba9da380a8b8a576['h07252] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0392a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07254] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0392b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07256] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0392c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07258] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0392d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0725a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0392e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0725c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0392f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0725e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03930] =  I8a0037ad2845a3fbba9da380a8b8a576['h07260] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03931] =  I8a0037ad2845a3fbba9da380a8b8a576['h07262] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03932] =  I8a0037ad2845a3fbba9da380a8b8a576['h07264] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03933] =  I8a0037ad2845a3fbba9da380a8b8a576['h07266] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03934] =  I8a0037ad2845a3fbba9da380a8b8a576['h07268] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03935] =  I8a0037ad2845a3fbba9da380a8b8a576['h0726a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03936] =  I8a0037ad2845a3fbba9da380a8b8a576['h0726c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03937] =  I8a0037ad2845a3fbba9da380a8b8a576['h0726e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03938] =  I8a0037ad2845a3fbba9da380a8b8a576['h07270] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03939] =  I8a0037ad2845a3fbba9da380a8b8a576['h07272] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0393a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07274] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0393b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07276] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0393c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07278] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0393d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0727a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0393e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0727c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0393f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0727e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03940] =  I8a0037ad2845a3fbba9da380a8b8a576['h07280] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03941] =  I8a0037ad2845a3fbba9da380a8b8a576['h07282] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03942] =  I8a0037ad2845a3fbba9da380a8b8a576['h07284] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03943] =  I8a0037ad2845a3fbba9da380a8b8a576['h07286] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03944] =  I8a0037ad2845a3fbba9da380a8b8a576['h07288] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03945] =  I8a0037ad2845a3fbba9da380a8b8a576['h0728a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03946] =  I8a0037ad2845a3fbba9da380a8b8a576['h0728c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03947] =  I8a0037ad2845a3fbba9da380a8b8a576['h0728e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03948] =  I8a0037ad2845a3fbba9da380a8b8a576['h07290] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03949] =  I8a0037ad2845a3fbba9da380a8b8a576['h07292] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0394a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07294] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0394b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07296] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0394c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07298] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0394d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0729a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0394e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0729c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0394f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0729e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03950] =  I8a0037ad2845a3fbba9da380a8b8a576['h072a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03951] =  I8a0037ad2845a3fbba9da380a8b8a576['h072a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03952] =  I8a0037ad2845a3fbba9da380a8b8a576['h072a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03953] =  I8a0037ad2845a3fbba9da380a8b8a576['h072a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03954] =  I8a0037ad2845a3fbba9da380a8b8a576['h072a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03955] =  I8a0037ad2845a3fbba9da380a8b8a576['h072aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03956] =  I8a0037ad2845a3fbba9da380a8b8a576['h072ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03957] =  I8a0037ad2845a3fbba9da380a8b8a576['h072ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03958] =  I8a0037ad2845a3fbba9da380a8b8a576['h072b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03959] =  I8a0037ad2845a3fbba9da380a8b8a576['h072b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0395a] =  I8a0037ad2845a3fbba9da380a8b8a576['h072b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0395b] =  I8a0037ad2845a3fbba9da380a8b8a576['h072b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0395c] =  I8a0037ad2845a3fbba9da380a8b8a576['h072b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0395d] =  I8a0037ad2845a3fbba9da380a8b8a576['h072ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0395e] =  I8a0037ad2845a3fbba9da380a8b8a576['h072bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0395f] =  I8a0037ad2845a3fbba9da380a8b8a576['h072be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03960] =  I8a0037ad2845a3fbba9da380a8b8a576['h072c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03961] =  I8a0037ad2845a3fbba9da380a8b8a576['h072c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03962] =  I8a0037ad2845a3fbba9da380a8b8a576['h072c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03963] =  I8a0037ad2845a3fbba9da380a8b8a576['h072c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03964] =  I8a0037ad2845a3fbba9da380a8b8a576['h072c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03965] =  I8a0037ad2845a3fbba9da380a8b8a576['h072ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03966] =  I8a0037ad2845a3fbba9da380a8b8a576['h072cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03967] =  I8a0037ad2845a3fbba9da380a8b8a576['h072ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03968] =  I8a0037ad2845a3fbba9da380a8b8a576['h072d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03969] =  I8a0037ad2845a3fbba9da380a8b8a576['h072d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0396a] =  I8a0037ad2845a3fbba9da380a8b8a576['h072d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0396b] =  I8a0037ad2845a3fbba9da380a8b8a576['h072d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0396c] =  I8a0037ad2845a3fbba9da380a8b8a576['h072d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0396d] =  I8a0037ad2845a3fbba9da380a8b8a576['h072da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0396e] =  I8a0037ad2845a3fbba9da380a8b8a576['h072dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0396f] =  I8a0037ad2845a3fbba9da380a8b8a576['h072de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03970] =  I8a0037ad2845a3fbba9da380a8b8a576['h072e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03971] =  I8a0037ad2845a3fbba9da380a8b8a576['h072e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03972] =  I8a0037ad2845a3fbba9da380a8b8a576['h072e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03973] =  I8a0037ad2845a3fbba9da380a8b8a576['h072e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03974] =  I8a0037ad2845a3fbba9da380a8b8a576['h072e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03975] =  I8a0037ad2845a3fbba9da380a8b8a576['h072ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03976] =  I8a0037ad2845a3fbba9da380a8b8a576['h072ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03977] =  I8a0037ad2845a3fbba9da380a8b8a576['h072ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03978] =  I8a0037ad2845a3fbba9da380a8b8a576['h072f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03979] =  I8a0037ad2845a3fbba9da380a8b8a576['h072f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0397a] =  I8a0037ad2845a3fbba9da380a8b8a576['h072f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0397b] =  I8a0037ad2845a3fbba9da380a8b8a576['h072f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0397c] =  I8a0037ad2845a3fbba9da380a8b8a576['h072f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0397d] =  I8a0037ad2845a3fbba9da380a8b8a576['h072fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0397e] =  I8a0037ad2845a3fbba9da380a8b8a576['h072fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0397f] =  I8a0037ad2845a3fbba9da380a8b8a576['h072fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03980] =  I8a0037ad2845a3fbba9da380a8b8a576['h07300] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03981] =  I8a0037ad2845a3fbba9da380a8b8a576['h07302] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03982] =  I8a0037ad2845a3fbba9da380a8b8a576['h07304] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03983] =  I8a0037ad2845a3fbba9da380a8b8a576['h07306] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03984] =  I8a0037ad2845a3fbba9da380a8b8a576['h07308] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03985] =  I8a0037ad2845a3fbba9da380a8b8a576['h0730a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03986] =  I8a0037ad2845a3fbba9da380a8b8a576['h0730c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03987] =  I8a0037ad2845a3fbba9da380a8b8a576['h0730e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03988] =  I8a0037ad2845a3fbba9da380a8b8a576['h07310] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03989] =  I8a0037ad2845a3fbba9da380a8b8a576['h07312] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0398a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07314] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0398b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07316] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0398c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07318] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0398d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0731a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0398e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0731c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0398f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0731e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03990] =  I8a0037ad2845a3fbba9da380a8b8a576['h07320] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03991] =  I8a0037ad2845a3fbba9da380a8b8a576['h07322] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03992] =  I8a0037ad2845a3fbba9da380a8b8a576['h07324] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03993] =  I8a0037ad2845a3fbba9da380a8b8a576['h07326] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03994] =  I8a0037ad2845a3fbba9da380a8b8a576['h07328] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03995] =  I8a0037ad2845a3fbba9da380a8b8a576['h0732a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03996] =  I8a0037ad2845a3fbba9da380a8b8a576['h0732c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03997] =  I8a0037ad2845a3fbba9da380a8b8a576['h0732e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03998] =  I8a0037ad2845a3fbba9da380a8b8a576['h07330] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03999] =  I8a0037ad2845a3fbba9da380a8b8a576['h07332] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0399a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07334] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0399b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07336] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0399c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07338] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0399d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0733a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0399e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0733c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h0399f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0733e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039a0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07340] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039a1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07342] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039a2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07344] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039a3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07346] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039a4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07348] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039a5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0734a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039a6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0734c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039a7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0734e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039a8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07350] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039a9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07352] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039aa] =  I8a0037ad2845a3fbba9da380a8b8a576['h07354] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039ab] =  I8a0037ad2845a3fbba9da380a8b8a576['h07356] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039ac] =  I8a0037ad2845a3fbba9da380a8b8a576['h07358] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039ad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0735a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039ae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0735c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039af] =  I8a0037ad2845a3fbba9da380a8b8a576['h0735e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039b0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07360] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039b1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07362] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039b2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07364] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039b3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07366] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039b4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07368] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039b5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0736a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039b6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0736c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039b7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0736e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039b8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07370] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039b9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07372] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039ba] =  I8a0037ad2845a3fbba9da380a8b8a576['h07374] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039bb] =  I8a0037ad2845a3fbba9da380a8b8a576['h07376] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039bc] =  I8a0037ad2845a3fbba9da380a8b8a576['h07378] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039bd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0737a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039be] =  I8a0037ad2845a3fbba9da380a8b8a576['h0737c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039bf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0737e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039c0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07380] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039c1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07382] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039c2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07384] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039c3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07386] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039c4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07388] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039c5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0738a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039c6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0738c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039c7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0738e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039c8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07390] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039c9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07392] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039ca] =  I8a0037ad2845a3fbba9da380a8b8a576['h07394] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039cb] =  I8a0037ad2845a3fbba9da380a8b8a576['h07396] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039cc] =  I8a0037ad2845a3fbba9da380a8b8a576['h07398] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039cd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0739a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039ce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0739c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039cf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0739e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039d0] =  I8a0037ad2845a3fbba9da380a8b8a576['h073a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039d1] =  I8a0037ad2845a3fbba9da380a8b8a576['h073a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039d2] =  I8a0037ad2845a3fbba9da380a8b8a576['h073a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039d3] =  I8a0037ad2845a3fbba9da380a8b8a576['h073a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039d4] =  I8a0037ad2845a3fbba9da380a8b8a576['h073a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039d5] =  I8a0037ad2845a3fbba9da380a8b8a576['h073aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039d6] =  I8a0037ad2845a3fbba9da380a8b8a576['h073ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039d7] =  I8a0037ad2845a3fbba9da380a8b8a576['h073ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039d8] =  I8a0037ad2845a3fbba9da380a8b8a576['h073b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039d9] =  I8a0037ad2845a3fbba9da380a8b8a576['h073b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039da] =  I8a0037ad2845a3fbba9da380a8b8a576['h073b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039db] =  I8a0037ad2845a3fbba9da380a8b8a576['h073b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039dc] =  I8a0037ad2845a3fbba9da380a8b8a576['h073b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039dd] =  I8a0037ad2845a3fbba9da380a8b8a576['h073ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039de] =  I8a0037ad2845a3fbba9da380a8b8a576['h073bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039df] =  I8a0037ad2845a3fbba9da380a8b8a576['h073be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039e0] =  I8a0037ad2845a3fbba9da380a8b8a576['h073c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039e1] =  I8a0037ad2845a3fbba9da380a8b8a576['h073c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039e2] =  I8a0037ad2845a3fbba9da380a8b8a576['h073c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039e3] =  I8a0037ad2845a3fbba9da380a8b8a576['h073c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039e4] =  I8a0037ad2845a3fbba9da380a8b8a576['h073c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039e5] =  I8a0037ad2845a3fbba9da380a8b8a576['h073ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039e6] =  I8a0037ad2845a3fbba9da380a8b8a576['h073cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039e7] =  I8a0037ad2845a3fbba9da380a8b8a576['h073ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039e8] =  I8a0037ad2845a3fbba9da380a8b8a576['h073d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039e9] =  I8a0037ad2845a3fbba9da380a8b8a576['h073d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039ea] =  I8a0037ad2845a3fbba9da380a8b8a576['h073d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039eb] =  I8a0037ad2845a3fbba9da380a8b8a576['h073d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039ec] =  I8a0037ad2845a3fbba9da380a8b8a576['h073d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039ed] =  I8a0037ad2845a3fbba9da380a8b8a576['h073da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039ee] =  I8a0037ad2845a3fbba9da380a8b8a576['h073dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039ef] =  I8a0037ad2845a3fbba9da380a8b8a576['h073de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039f0] =  I8a0037ad2845a3fbba9da380a8b8a576['h073e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039f1] =  I8a0037ad2845a3fbba9da380a8b8a576['h073e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039f2] =  I8a0037ad2845a3fbba9da380a8b8a576['h073e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039f3] =  I8a0037ad2845a3fbba9da380a8b8a576['h073e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039f4] =  I8a0037ad2845a3fbba9da380a8b8a576['h073e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039f5] =  I8a0037ad2845a3fbba9da380a8b8a576['h073ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039f6] =  I8a0037ad2845a3fbba9da380a8b8a576['h073ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039f7] =  I8a0037ad2845a3fbba9da380a8b8a576['h073ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039f8] =  I8a0037ad2845a3fbba9da380a8b8a576['h073f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039f9] =  I8a0037ad2845a3fbba9da380a8b8a576['h073f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039fa] =  I8a0037ad2845a3fbba9da380a8b8a576['h073f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039fb] =  I8a0037ad2845a3fbba9da380a8b8a576['h073f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039fc] =  I8a0037ad2845a3fbba9da380a8b8a576['h073f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039fd] =  I8a0037ad2845a3fbba9da380a8b8a576['h073fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039fe] =  I8a0037ad2845a3fbba9da380a8b8a576['h073fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h039ff] =  I8a0037ad2845a3fbba9da380a8b8a576['h073fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a00] =  I8a0037ad2845a3fbba9da380a8b8a576['h07400] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a01] =  I8a0037ad2845a3fbba9da380a8b8a576['h07402] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a02] =  I8a0037ad2845a3fbba9da380a8b8a576['h07404] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a03] =  I8a0037ad2845a3fbba9da380a8b8a576['h07406] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a04] =  I8a0037ad2845a3fbba9da380a8b8a576['h07408] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a05] =  I8a0037ad2845a3fbba9da380a8b8a576['h0740a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a06] =  I8a0037ad2845a3fbba9da380a8b8a576['h0740c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a07] =  I8a0037ad2845a3fbba9da380a8b8a576['h0740e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a08] =  I8a0037ad2845a3fbba9da380a8b8a576['h07410] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a09] =  I8a0037ad2845a3fbba9da380a8b8a576['h07412] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a0a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07414] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a0b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07416] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a0c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07418] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a0d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0741a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a0e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0741c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a0f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0741e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a10] =  I8a0037ad2845a3fbba9da380a8b8a576['h07420] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a11] =  I8a0037ad2845a3fbba9da380a8b8a576['h07422] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a12] =  I8a0037ad2845a3fbba9da380a8b8a576['h07424] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a13] =  I8a0037ad2845a3fbba9da380a8b8a576['h07426] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a14] =  I8a0037ad2845a3fbba9da380a8b8a576['h07428] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a15] =  I8a0037ad2845a3fbba9da380a8b8a576['h0742a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a16] =  I8a0037ad2845a3fbba9da380a8b8a576['h0742c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a17] =  I8a0037ad2845a3fbba9da380a8b8a576['h0742e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a18] =  I8a0037ad2845a3fbba9da380a8b8a576['h07430] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a19] =  I8a0037ad2845a3fbba9da380a8b8a576['h07432] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a1a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07434] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a1b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07436] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a1c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07438] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a1d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0743a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a1e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0743c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a1f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0743e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a20] =  I8a0037ad2845a3fbba9da380a8b8a576['h07440] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a21] =  I8a0037ad2845a3fbba9da380a8b8a576['h07442] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a22] =  I8a0037ad2845a3fbba9da380a8b8a576['h07444] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a23] =  I8a0037ad2845a3fbba9da380a8b8a576['h07446] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a24] =  I8a0037ad2845a3fbba9da380a8b8a576['h07448] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a25] =  I8a0037ad2845a3fbba9da380a8b8a576['h0744a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a26] =  I8a0037ad2845a3fbba9da380a8b8a576['h0744c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a27] =  I8a0037ad2845a3fbba9da380a8b8a576['h0744e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a28] =  I8a0037ad2845a3fbba9da380a8b8a576['h07450] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a29] =  I8a0037ad2845a3fbba9da380a8b8a576['h07452] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a2a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07454] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a2b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07456] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a2c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07458] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a2d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0745a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a2e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0745c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a2f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0745e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a30] =  I8a0037ad2845a3fbba9da380a8b8a576['h07460] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a31] =  I8a0037ad2845a3fbba9da380a8b8a576['h07462] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a32] =  I8a0037ad2845a3fbba9da380a8b8a576['h07464] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a33] =  I8a0037ad2845a3fbba9da380a8b8a576['h07466] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a34] =  I8a0037ad2845a3fbba9da380a8b8a576['h07468] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a35] =  I8a0037ad2845a3fbba9da380a8b8a576['h0746a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a36] =  I8a0037ad2845a3fbba9da380a8b8a576['h0746c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a37] =  I8a0037ad2845a3fbba9da380a8b8a576['h0746e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a38] =  I8a0037ad2845a3fbba9da380a8b8a576['h07470] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a39] =  I8a0037ad2845a3fbba9da380a8b8a576['h07472] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a3a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07474] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a3b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07476] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a3c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07478] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a3d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0747a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a3e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0747c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a3f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0747e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a40] =  I8a0037ad2845a3fbba9da380a8b8a576['h07480] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a41] =  I8a0037ad2845a3fbba9da380a8b8a576['h07482] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a42] =  I8a0037ad2845a3fbba9da380a8b8a576['h07484] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a43] =  I8a0037ad2845a3fbba9da380a8b8a576['h07486] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a44] =  I8a0037ad2845a3fbba9da380a8b8a576['h07488] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a45] =  I8a0037ad2845a3fbba9da380a8b8a576['h0748a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a46] =  I8a0037ad2845a3fbba9da380a8b8a576['h0748c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a47] =  I8a0037ad2845a3fbba9da380a8b8a576['h0748e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a48] =  I8a0037ad2845a3fbba9da380a8b8a576['h07490] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a49] =  I8a0037ad2845a3fbba9da380a8b8a576['h07492] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a4a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07494] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a4b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07496] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a4c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07498] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a4d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0749a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a4e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0749c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a4f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0749e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a50] =  I8a0037ad2845a3fbba9da380a8b8a576['h074a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a51] =  I8a0037ad2845a3fbba9da380a8b8a576['h074a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a52] =  I8a0037ad2845a3fbba9da380a8b8a576['h074a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a53] =  I8a0037ad2845a3fbba9da380a8b8a576['h074a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a54] =  I8a0037ad2845a3fbba9da380a8b8a576['h074a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a55] =  I8a0037ad2845a3fbba9da380a8b8a576['h074aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a56] =  I8a0037ad2845a3fbba9da380a8b8a576['h074ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a57] =  I8a0037ad2845a3fbba9da380a8b8a576['h074ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a58] =  I8a0037ad2845a3fbba9da380a8b8a576['h074b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a59] =  I8a0037ad2845a3fbba9da380a8b8a576['h074b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a5a] =  I8a0037ad2845a3fbba9da380a8b8a576['h074b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a5b] =  I8a0037ad2845a3fbba9da380a8b8a576['h074b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a5c] =  I8a0037ad2845a3fbba9da380a8b8a576['h074b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a5d] =  I8a0037ad2845a3fbba9da380a8b8a576['h074ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a5e] =  I8a0037ad2845a3fbba9da380a8b8a576['h074bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a5f] =  I8a0037ad2845a3fbba9da380a8b8a576['h074be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a60] =  I8a0037ad2845a3fbba9da380a8b8a576['h074c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a61] =  I8a0037ad2845a3fbba9da380a8b8a576['h074c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a62] =  I8a0037ad2845a3fbba9da380a8b8a576['h074c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a63] =  I8a0037ad2845a3fbba9da380a8b8a576['h074c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a64] =  I8a0037ad2845a3fbba9da380a8b8a576['h074c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a65] =  I8a0037ad2845a3fbba9da380a8b8a576['h074ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a66] =  I8a0037ad2845a3fbba9da380a8b8a576['h074cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a67] =  I8a0037ad2845a3fbba9da380a8b8a576['h074ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a68] =  I8a0037ad2845a3fbba9da380a8b8a576['h074d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a69] =  I8a0037ad2845a3fbba9da380a8b8a576['h074d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a6a] =  I8a0037ad2845a3fbba9da380a8b8a576['h074d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a6b] =  I8a0037ad2845a3fbba9da380a8b8a576['h074d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a6c] =  I8a0037ad2845a3fbba9da380a8b8a576['h074d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a6d] =  I8a0037ad2845a3fbba9da380a8b8a576['h074da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a6e] =  I8a0037ad2845a3fbba9da380a8b8a576['h074dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a6f] =  I8a0037ad2845a3fbba9da380a8b8a576['h074de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a70] =  I8a0037ad2845a3fbba9da380a8b8a576['h074e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a71] =  I8a0037ad2845a3fbba9da380a8b8a576['h074e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a72] =  I8a0037ad2845a3fbba9da380a8b8a576['h074e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a73] =  I8a0037ad2845a3fbba9da380a8b8a576['h074e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a74] =  I8a0037ad2845a3fbba9da380a8b8a576['h074e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a75] =  I8a0037ad2845a3fbba9da380a8b8a576['h074ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a76] =  I8a0037ad2845a3fbba9da380a8b8a576['h074ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a77] =  I8a0037ad2845a3fbba9da380a8b8a576['h074ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a78] =  I8a0037ad2845a3fbba9da380a8b8a576['h074f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a79] =  I8a0037ad2845a3fbba9da380a8b8a576['h074f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a7a] =  I8a0037ad2845a3fbba9da380a8b8a576['h074f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a7b] =  I8a0037ad2845a3fbba9da380a8b8a576['h074f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a7c] =  I8a0037ad2845a3fbba9da380a8b8a576['h074f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a7d] =  I8a0037ad2845a3fbba9da380a8b8a576['h074fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a7e] =  I8a0037ad2845a3fbba9da380a8b8a576['h074fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a7f] =  I8a0037ad2845a3fbba9da380a8b8a576['h074fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a80] =  I8a0037ad2845a3fbba9da380a8b8a576['h07500] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a81] =  I8a0037ad2845a3fbba9da380a8b8a576['h07502] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a82] =  I8a0037ad2845a3fbba9da380a8b8a576['h07504] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a83] =  I8a0037ad2845a3fbba9da380a8b8a576['h07506] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a84] =  I8a0037ad2845a3fbba9da380a8b8a576['h07508] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a85] =  I8a0037ad2845a3fbba9da380a8b8a576['h0750a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a86] =  I8a0037ad2845a3fbba9da380a8b8a576['h0750c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a87] =  I8a0037ad2845a3fbba9da380a8b8a576['h0750e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a88] =  I8a0037ad2845a3fbba9da380a8b8a576['h07510] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a89] =  I8a0037ad2845a3fbba9da380a8b8a576['h07512] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a8a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07514] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a8b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07516] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a8c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07518] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a8d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0751a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a8e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0751c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a8f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0751e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a90] =  I8a0037ad2845a3fbba9da380a8b8a576['h07520] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a91] =  I8a0037ad2845a3fbba9da380a8b8a576['h07522] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a92] =  I8a0037ad2845a3fbba9da380a8b8a576['h07524] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a93] =  I8a0037ad2845a3fbba9da380a8b8a576['h07526] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a94] =  I8a0037ad2845a3fbba9da380a8b8a576['h07528] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a95] =  I8a0037ad2845a3fbba9da380a8b8a576['h0752a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a96] =  I8a0037ad2845a3fbba9da380a8b8a576['h0752c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a97] =  I8a0037ad2845a3fbba9da380a8b8a576['h0752e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a98] =  I8a0037ad2845a3fbba9da380a8b8a576['h07530] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a99] =  I8a0037ad2845a3fbba9da380a8b8a576['h07532] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a9a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07534] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a9b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07536] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a9c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07538] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a9d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0753a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a9e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0753c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03a9f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0753e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03aa0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07540] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03aa1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07542] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03aa2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07544] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03aa3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07546] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03aa4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07548] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03aa5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0754a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03aa6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0754c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03aa7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0754e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03aa8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07550] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03aa9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07552] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03aaa] =  I8a0037ad2845a3fbba9da380a8b8a576['h07554] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03aab] =  I8a0037ad2845a3fbba9da380a8b8a576['h07556] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03aac] =  I8a0037ad2845a3fbba9da380a8b8a576['h07558] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03aad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0755a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03aae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0755c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03aaf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0755e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ab0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07560] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ab1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07562] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ab2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07564] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ab3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07566] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ab4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07568] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ab5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0756a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ab6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0756c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ab7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0756e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ab8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07570] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ab9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07572] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03aba] =  I8a0037ad2845a3fbba9da380a8b8a576['h07574] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03abb] =  I8a0037ad2845a3fbba9da380a8b8a576['h07576] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03abc] =  I8a0037ad2845a3fbba9da380a8b8a576['h07578] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03abd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0757a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03abe] =  I8a0037ad2845a3fbba9da380a8b8a576['h0757c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03abf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0757e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ac0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07580] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ac1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07582] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ac2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07584] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ac3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07586] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ac4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07588] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ac5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0758a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ac6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0758c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ac7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0758e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ac8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07590] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ac9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07592] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03aca] =  I8a0037ad2845a3fbba9da380a8b8a576['h07594] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03acb] =  I8a0037ad2845a3fbba9da380a8b8a576['h07596] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03acc] =  I8a0037ad2845a3fbba9da380a8b8a576['h07598] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03acd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0759a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ace] =  I8a0037ad2845a3fbba9da380a8b8a576['h0759c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03acf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0759e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ad0] =  I8a0037ad2845a3fbba9da380a8b8a576['h075a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ad1] =  I8a0037ad2845a3fbba9da380a8b8a576['h075a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ad2] =  I8a0037ad2845a3fbba9da380a8b8a576['h075a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ad3] =  I8a0037ad2845a3fbba9da380a8b8a576['h075a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ad4] =  I8a0037ad2845a3fbba9da380a8b8a576['h075a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ad5] =  I8a0037ad2845a3fbba9da380a8b8a576['h075aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ad6] =  I8a0037ad2845a3fbba9da380a8b8a576['h075ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ad7] =  I8a0037ad2845a3fbba9da380a8b8a576['h075ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ad8] =  I8a0037ad2845a3fbba9da380a8b8a576['h075b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ad9] =  I8a0037ad2845a3fbba9da380a8b8a576['h075b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ada] =  I8a0037ad2845a3fbba9da380a8b8a576['h075b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03adb] =  I8a0037ad2845a3fbba9da380a8b8a576['h075b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03adc] =  I8a0037ad2845a3fbba9da380a8b8a576['h075b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03add] =  I8a0037ad2845a3fbba9da380a8b8a576['h075ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ade] =  I8a0037ad2845a3fbba9da380a8b8a576['h075bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03adf] =  I8a0037ad2845a3fbba9da380a8b8a576['h075be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ae0] =  I8a0037ad2845a3fbba9da380a8b8a576['h075c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ae1] =  I8a0037ad2845a3fbba9da380a8b8a576['h075c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ae2] =  I8a0037ad2845a3fbba9da380a8b8a576['h075c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ae3] =  I8a0037ad2845a3fbba9da380a8b8a576['h075c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ae4] =  I8a0037ad2845a3fbba9da380a8b8a576['h075c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ae5] =  I8a0037ad2845a3fbba9da380a8b8a576['h075ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ae6] =  I8a0037ad2845a3fbba9da380a8b8a576['h075cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ae7] =  I8a0037ad2845a3fbba9da380a8b8a576['h075ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ae8] =  I8a0037ad2845a3fbba9da380a8b8a576['h075d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ae9] =  I8a0037ad2845a3fbba9da380a8b8a576['h075d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03aea] =  I8a0037ad2845a3fbba9da380a8b8a576['h075d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03aeb] =  I8a0037ad2845a3fbba9da380a8b8a576['h075d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03aec] =  I8a0037ad2845a3fbba9da380a8b8a576['h075d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03aed] =  I8a0037ad2845a3fbba9da380a8b8a576['h075da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03aee] =  I8a0037ad2845a3fbba9da380a8b8a576['h075dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03aef] =  I8a0037ad2845a3fbba9da380a8b8a576['h075de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03af0] =  I8a0037ad2845a3fbba9da380a8b8a576['h075e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03af1] =  I8a0037ad2845a3fbba9da380a8b8a576['h075e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03af2] =  I8a0037ad2845a3fbba9da380a8b8a576['h075e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03af3] =  I8a0037ad2845a3fbba9da380a8b8a576['h075e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03af4] =  I8a0037ad2845a3fbba9da380a8b8a576['h075e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03af5] =  I8a0037ad2845a3fbba9da380a8b8a576['h075ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03af6] =  I8a0037ad2845a3fbba9da380a8b8a576['h075ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03af7] =  I8a0037ad2845a3fbba9da380a8b8a576['h075ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03af8] =  I8a0037ad2845a3fbba9da380a8b8a576['h075f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03af9] =  I8a0037ad2845a3fbba9da380a8b8a576['h075f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03afa] =  I8a0037ad2845a3fbba9da380a8b8a576['h075f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03afb] =  I8a0037ad2845a3fbba9da380a8b8a576['h075f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03afc] =  I8a0037ad2845a3fbba9da380a8b8a576['h075f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03afd] =  I8a0037ad2845a3fbba9da380a8b8a576['h075fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03afe] =  I8a0037ad2845a3fbba9da380a8b8a576['h075fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03aff] =  I8a0037ad2845a3fbba9da380a8b8a576['h075fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b00] =  I8a0037ad2845a3fbba9da380a8b8a576['h07600] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b01] =  I8a0037ad2845a3fbba9da380a8b8a576['h07602] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b02] =  I8a0037ad2845a3fbba9da380a8b8a576['h07604] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b03] =  I8a0037ad2845a3fbba9da380a8b8a576['h07606] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b04] =  I8a0037ad2845a3fbba9da380a8b8a576['h07608] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b05] =  I8a0037ad2845a3fbba9da380a8b8a576['h0760a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b06] =  I8a0037ad2845a3fbba9da380a8b8a576['h0760c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b07] =  I8a0037ad2845a3fbba9da380a8b8a576['h0760e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b08] =  I8a0037ad2845a3fbba9da380a8b8a576['h07610] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b09] =  I8a0037ad2845a3fbba9da380a8b8a576['h07612] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b0a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07614] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b0b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07616] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b0c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07618] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b0d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0761a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b0e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0761c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b0f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0761e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b10] =  I8a0037ad2845a3fbba9da380a8b8a576['h07620] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b11] =  I8a0037ad2845a3fbba9da380a8b8a576['h07622] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b12] =  I8a0037ad2845a3fbba9da380a8b8a576['h07624] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b13] =  I8a0037ad2845a3fbba9da380a8b8a576['h07626] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b14] =  I8a0037ad2845a3fbba9da380a8b8a576['h07628] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b15] =  I8a0037ad2845a3fbba9da380a8b8a576['h0762a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b16] =  I8a0037ad2845a3fbba9da380a8b8a576['h0762c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b17] =  I8a0037ad2845a3fbba9da380a8b8a576['h0762e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b18] =  I8a0037ad2845a3fbba9da380a8b8a576['h07630] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b19] =  I8a0037ad2845a3fbba9da380a8b8a576['h07632] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b1a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07634] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b1b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07636] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b1c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07638] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b1d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0763a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b1e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0763c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b1f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0763e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b20] =  I8a0037ad2845a3fbba9da380a8b8a576['h07640] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b21] =  I8a0037ad2845a3fbba9da380a8b8a576['h07642] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b22] =  I8a0037ad2845a3fbba9da380a8b8a576['h07644] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b23] =  I8a0037ad2845a3fbba9da380a8b8a576['h07646] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b24] =  I8a0037ad2845a3fbba9da380a8b8a576['h07648] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b25] =  I8a0037ad2845a3fbba9da380a8b8a576['h0764a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b26] =  I8a0037ad2845a3fbba9da380a8b8a576['h0764c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b27] =  I8a0037ad2845a3fbba9da380a8b8a576['h0764e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b28] =  I8a0037ad2845a3fbba9da380a8b8a576['h07650] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b29] =  I8a0037ad2845a3fbba9da380a8b8a576['h07652] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b2a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07654] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b2b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07656] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b2c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07658] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b2d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0765a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b2e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0765c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b2f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0765e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b30] =  I8a0037ad2845a3fbba9da380a8b8a576['h07660] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b31] =  I8a0037ad2845a3fbba9da380a8b8a576['h07662] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b32] =  I8a0037ad2845a3fbba9da380a8b8a576['h07664] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b33] =  I8a0037ad2845a3fbba9da380a8b8a576['h07666] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b34] =  I8a0037ad2845a3fbba9da380a8b8a576['h07668] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b35] =  I8a0037ad2845a3fbba9da380a8b8a576['h0766a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b36] =  I8a0037ad2845a3fbba9da380a8b8a576['h0766c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b37] =  I8a0037ad2845a3fbba9da380a8b8a576['h0766e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b38] =  I8a0037ad2845a3fbba9da380a8b8a576['h07670] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b39] =  I8a0037ad2845a3fbba9da380a8b8a576['h07672] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b3a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07674] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b3b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07676] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b3c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07678] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b3d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0767a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b3e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0767c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b3f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0767e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b40] =  I8a0037ad2845a3fbba9da380a8b8a576['h07680] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b41] =  I8a0037ad2845a3fbba9da380a8b8a576['h07682] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b42] =  I8a0037ad2845a3fbba9da380a8b8a576['h07684] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b43] =  I8a0037ad2845a3fbba9da380a8b8a576['h07686] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b44] =  I8a0037ad2845a3fbba9da380a8b8a576['h07688] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b45] =  I8a0037ad2845a3fbba9da380a8b8a576['h0768a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b46] =  I8a0037ad2845a3fbba9da380a8b8a576['h0768c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b47] =  I8a0037ad2845a3fbba9da380a8b8a576['h0768e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b48] =  I8a0037ad2845a3fbba9da380a8b8a576['h07690] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b49] =  I8a0037ad2845a3fbba9da380a8b8a576['h07692] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b4a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07694] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b4b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07696] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b4c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07698] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b4d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0769a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b4e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0769c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b4f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0769e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b50] =  I8a0037ad2845a3fbba9da380a8b8a576['h076a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b51] =  I8a0037ad2845a3fbba9da380a8b8a576['h076a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b52] =  I8a0037ad2845a3fbba9da380a8b8a576['h076a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b53] =  I8a0037ad2845a3fbba9da380a8b8a576['h076a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b54] =  I8a0037ad2845a3fbba9da380a8b8a576['h076a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b55] =  I8a0037ad2845a3fbba9da380a8b8a576['h076aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b56] =  I8a0037ad2845a3fbba9da380a8b8a576['h076ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b57] =  I8a0037ad2845a3fbba9da380a8b8a576['h076ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b58] =  I8a0037ad2845a3fbba9da380a8b8a576['h076b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b59] =  I8a0037ad2845a3fbba9da380a8b8a576['h076b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b5a] =  I8a0037ad2845a3fbba9da380a8b8a576['h076b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b5b] =  I8a0037ad2845a3fbba9da380a8b8a576['h076b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b5c] =  I8a0037ad2845a3fbba9da380a8b8a576['h076b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b5d] =  I8a0037ad2845a3fbba9da380a8b8a576['h076ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b5e] =  I8a0037ad2845a3fbba9da380a8b8a576['h076bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b5f] =  I8a0037ad2845a3fbba9da380a8b8a576['h076be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b60] =  I8a0037ad2845a3fbba9da380a8b8a576['h076c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b61] =  I8a0037ad2845a3fbba9da380a8b8a576['h076c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b62] =  I8a0037ad2845a3fbba9da380a8b8a576['h076c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b63] =  I8a0037ad2845a3fbba9da380a8b8a576['h076c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b64] =  I8a0037ad2845a3fbba9da380a8b8a576['h076c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b65] =  I8a0037ad2845a3fbba9da380a8b8a576['h076ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b66] =  I8a0037ad2845a3fbba9da380a8b8a576['h076cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b67] =  I8a0037ad2845a3fbba9da380a8b8a576['h076ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b68] =  I8a0037ad2845a3fbba9da380a8b8a576['h076d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b69] =  I8a0037ad2845a3fbba9da380a8b8a576['h076d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b6a] =  I8a0037ad2845a3fbba9da380a8b8a576['h076d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b6b] =  I8a0037ad2845a3fbba9da380a8b8a576['h076d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b6c] =  I8a0037ad2845a3fbba9da380a8b8a576['h076d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b6d] =  I8a0037ad2845a3fbba9da380a8b8a576['h076da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b6e] =  I8a0037ad2845a3fbba9da380a8b8a576['h076dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b6f] =  I8a0037ad2845a3fbba9da380a8b8a576['h076de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b70] =  I8a0037ad2845a3fbba9da380a8b8a576['h076e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b71] =  I8a0037ad2845a3fbba9da380a8b8a576['h076e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b72] =  I8a0037ad2845a3fbba9da380a8b8a576['h076e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b73] =  I8a0037ad2845a3fbba9da380a8b8a576['h076e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b74] =  I8a0037ad2845a3fbba9da380a8b8a576['h076e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b75] =  I8a0037ad2845a3fbba9da380a8b8a576['h076ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b76] =  I8a0037ad2845a3fbba9da380a8b8a576['h076ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b77] =  I8a0037ad2845a3fbba9da380a8b8a576['h076ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b78] =  I8a0037ad2845a3fbba9da380a8b8a576['h076f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b79] =  I8a0037ad2845a3fbba9da380a8b8a576['h076f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b7a] =  I8a0037ad2845a3fbba9da380a8b8a576['h076f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b7b] =  I8a0037ad2845a3fbba9da380a8b8a576['h076f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b7c] =  I8a0037ad2845a3fbba9da380a8b8a576['h076f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b7d] =  I8a0037ad2845a3fbba9da380a8b8a576['h076fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b7e] =  I8a0037ad2845a3fbba9da380a8b8a576['h076fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b7f] =  I8a0037ad2845a3fbba9da380a8b8a576['h076fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b80] =  I8a0037ad2845a3fbba9da380a8b8a576['h07700] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b81] =  I8a0037ad2845a3fbba9da380a8b8a576['h07702] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b82] =  I8a0037ad2845a3fbba9da380a8b8a576['h07704] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b83] =  I8a0037ad2845a3fbba9da380a8b8a576['h07706] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b84] =  I8a0037ad2845a3fbba9da380a8b8a576['h07708] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b85] =  I8a0037ad2845a3fbba9da380a8b8a576['h0770a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b86] =  I8a0037ad2845a3fbba9da380a8b8a576['h0770c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b87] =  I8a0037ad2845a3fbba9da380a8b8a576['h0770e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b88] =  I8a0037ad2845a3fbba9da380a8b8a576['h07710] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b89] =  I8a0037ad2845a3fbba9da380a8b8a576['h07712] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b8a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07714] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b8b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07716] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b8c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07718] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b8d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0771a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b8e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0771c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b8f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0771e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b90] =  I8a0037ad2845a3fbba9da380a8b8a576['h07720] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b91] =  I8a0037ad2845a3fbba9da380a8b8a576['h07722] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b92] =  I8a0037ad2845a3fbba9da380a8b8a576['h07724] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b93] =  I8a0037ad2845a3fbba9da380a8b8a576['h07726] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b94] =  I8a0037ad2845a3fbba9da380a8b8a576['h07728] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b95] =  I8a0037ad2845a3fbba9da380a8b8a576['h0772a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b96] =  I8a0037ad2845a3fbba9da380a8b8a576['h0772c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b97] =  I8a0037ad2845a3fbba9da380a8b8a576['h0772e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b98] =  I8a0037ad2845a3fbba9da380a8b8a576['h07730] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b99] =  I8a0037ad2845a3fbba9da380a8b8a576['h07732] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b9a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07734] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b9b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07736] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b9c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07738] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b9d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0773a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b9e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0773c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03b9f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0773e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ba0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07740] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ba1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07742] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ba2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07744] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ba3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07746] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ba4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07748] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ba5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0774a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ba6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0774c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ba7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0774e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ba8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07750] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ba9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07752] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03baa] =  I8a0037ad2845a3fbba9da380a8b8a576['h07754] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bab] =  I8a0037ad2845a3fbba9da380a8b8a576['h07756] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bac] =  I8a0037ad2845a3fbba9da380a8b8a576['h07758] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0775a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0775c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03baf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0775e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bb0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07760] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bb1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07762] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bb2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07764] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bb3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07766] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bb4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07768] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bb5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0776a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bb6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0776c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bb7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0776e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bb8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07770] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bb9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07772] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bba] =  I8a0037ad2845a3fbba9da380a8b8a576['h07774] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bbb] =  I8a0037ad2845a3fbba9da380a8b8a576['h07776] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bbc] =  I8a0037ad2845a3fbba9da380a8b8a576['h07778] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bbd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0777a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bbe] =  I8a0037ad2845a3fbba9da380a8b8a576['h0777c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bbf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0777e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bc0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07780] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bc1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07782] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bc2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07784] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bc3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07786] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bc4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07788] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bc5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0778a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bc6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0778c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bc7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0778e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bc8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07790] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bc9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07792] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bca] =  I8a0037ad2845a3fbba9da380a8b8a576['h07794] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bcb] =  I8a0037ad2845a3fbba9da380a8b8a576['h07796] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bcc] =  I8a0037ad2845a3fbba9da380a8b8a576['h07798] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bcd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0779a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0779c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bcf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0779e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bd0] =  I8a0037ad2845a3fbba9da380a8b8a576['h077a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bd1] =  I8a0037ad2845a3fbba9da380a8b8a576['h077a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bd2] =  I8a0037ad2845a3fbba9da380a8b8a576['h077a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bd3] =  I8a0037ad2845a3fbba9da380a8b8a576['h077a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bd4] =  I8a0037ad2845a3fbba9da380a8b8a576['h077a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bd5] =  I8a0037ad2845a3fbba9da380a8b8a576['h077aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bd6] =  I8a0037ad2845a3fbba9da380a8b8a576['h077ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bd7] =  I8a0037ad2845a3fbba9da380a8b8a576['h077ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bd8] =  I8a0037ad2845a3fbba9da380a8b8a576['h077b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bd9] =  I8a0037ad2845a3fbba9da380a8b8a576['h077b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bda] =  I8a0037ad2845a3fbba9da380a8b8a576['h077b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bdb] =  I8a0037ad2845a3fbba9da380a8b8a576['h077b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bdc] =  I8a0037ad2845a3fbba9da380a8b8a576['h077b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bdd] =  I8a0037ad2845a3fbba9da380a8b8a576['h077ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bde] =  I8a0037ad2845a3fbba9da380a8b8a576['h077bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bdf] =  I8a0037ad2845a3fbba9da380a8b8a576['h077be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03be0] =  I8a0037ad2845a3fbba9da380a8b8a576['h077c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03be1] =  I8a0037ad2845a3fbba9da380a8b8a576['h077c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03be2] =  I8a0037ad2845a3fbba9da380a8b8a576['h077c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03be3] =  I8a0037ad2845a3fbba9da380a8b8a576['h077c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03be4] =  I8a0037ad2845a3fbba9da380a8b8a576['h077c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03be5] =  I8a0037ad2845a3fbba9da380a8b8a576['h077ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03be6] =  I8a0037ad2845a3fbba9da380a8b8a576['h077cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03be7] =  I8a0037ad2845a3fbba9da380a8b8a576['h077ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03be8] =  I8a0037ad2845a3fbba9da380a8b8a576['h077d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03be9] =  I8a0037ad2845a3fbba9da380a8b8a576['h077d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bea] =  I8a0037ad2845a3fbba9da380a8b8a576['h077d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03beb] =  I8a0037ad2845a3fbba9da380a8b8a576['h077d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bec] =  I8a0037ad2845a3fbba9da380a8b8a576['h077d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bed] =  I8a0037ad2845a3fbba9da380a8b8a576['h077da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bee] =  I8a0037ad2845a3fbba9da380a8b8a576['h077dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bef] =  I8a0037ad2845a3fbba9da380a8b8a576['h077de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bf0] =  I8a0037ad2845a3fbba9da380a8b8a576['h077e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bf1] =  I8a0037ad2845a3fbba9da380a8b8a576['h077e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bf2] =  I8a0037ad2845a3fbba9da380a8b8a576['h077e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bf3] =  I8a0037ad2845a3fbba9da380a8b8a576['h077e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bf4] =  I8a0037ad2845a3fbba9da380a8b8a576['h077e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bf5] =  I8a0037ad2845a3fbba9da380a8b8a576['h077ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bf6] =  I8a0037ad2845a3fbba9da380a8b8a576['h077ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bf7] =  I8a0037ad2845a3fbba9da380a8b8a576['h077ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bf8] =  I8a0037ad2845a3fbba9da380a8b8a576['h077f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bf9] =  I8a0037ad2845a3fbba9da380a8b8a576['h077f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bfa] =  I8a0037ad2845a3fbba9da380a8b8a576['h077f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bfb] =  I8a0037ad2845a3fbba9da380a8b8a576['h077f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bfc] =  I8a0037ad2845a3fbba9da380a8b8a576['h077f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bfd] =  I8a0037ad2845a3fbba9da380a8b8a576['h077fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bfe] =  I8a0037ad2845a3fbba9da380a8b8a576['h077fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03bff] =  I8a0037ad2845a3fbba9da380a8b8a576['h077fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c00] =  I8a0037ad2845a3fbba9da380a8b8a576['h07800] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c01] =  I8a0037ad2845a3fbba9da380a8b8a576['h07802] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c02] =  I8a0037ad2845a3fbba9da380a8b8a576['h07804] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c03] =  I8a0037ad2845a3fbba9da380a8b8a576['h07806] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c04] =  I8a0037ad2845a3fbba9da380a8b8a576['h07808] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c05] =  I8a0037ad2845a3fbba9da380a8b8a576['h0780a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c06] =  I8a0037ad2845a3fbba9da380a8b8a576['h0780c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c07] =  I8a0037ad2845a3fbba9da380a8b8a576['h0780e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c08] =  I8a0037ad2845a3fbba9da380a8b8a576['h07810] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c09] =  I8a0037ad2845a3fbba9da380a8b8a576['h07812] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c0a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07814] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c0b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07816] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c0c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07818] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c0d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0781a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c0e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0781c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c0f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0781e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c10] =  I8a0037ad2845a3fbba9da380a8b8a576['h07820] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c11] =  I8a0037ad2845a3fbba9da380a8b8a576['h07822] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c12] =  I8a0037ad2845a3fbba9da380a8b8a576['h07824] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c13] =  I8a0037ad2845a3fbba9da380a8b8a576['h07826] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c14] =  I8a0037ad2845a3fbba9da380a8b8a576['h07828] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c15] =  I8a0037ad2845a3fbba9da380a8b8a576['h0782a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c16] =  I8a0037ad2845a3fbba9da380a8b8a576['h0782c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c17] =  I8a0037ad2845a3fbba9da380a8b8a576['h0782e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c18] =  I8a0037ad2845a3fbba9da380a8b8a576['h07830] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c19] =  I8a0037ad2845a3fbba9da380a8b8a576['h07832] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c1a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07834] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c1b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07836] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c1c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07838] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c1d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0783a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c1e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0783c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c1f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0783e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c20] =  I8a0037ad2845a3fbba9da380a8b8a576['h07840] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c21] =  I8a0037ad2845a3fbba9da380a8b8a576['h07842] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c22] =  I8a0037ad2845a3fbba9da380a8b8a576['h07844] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c23] =  I8a0037ad2845a3fbba9da380a8b8a576['h07846] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c24] =  I8a0037ad2845a3fbba9da380a8b8a576['h07848] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c25] =  I8a0037ad2845a3fbba9da380a8b8a576['h0784a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c26] =  I8a0037ad2845a3fbba9da380a8b8a576['h0784c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c27] =  I8a0037ad2845a3fbba9da380a8b8a576['h0784e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c28] =  I8a0037ad2845a3fbba9da380a8b8a576['h07850] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c29] =  I8a0037ad2845a3fbba9da380a8b8a576['h07852] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c2a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07854] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c2b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07856] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c2c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07858] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c2d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0785a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c2e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0785c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c2f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0785e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c30] =  I8a0037ad2845a3fbba9da380a8b8a576['h07860] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c31] =  I8a0037ad2845a3fbba9da380a8b8a576['h07862] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c32] =  I8a0037ad2845a3fbba9da380a8b8a576['h07864] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c33] =  I8a0037ad2845a3fbba9da380a8b8a576['h07866] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c34] =  I8a0037ad2845a3fbba9da380a8b8a576['h07868] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c35] =  I8a0037ad2845a3fbba9da380a8b8a576['h0786a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c36] =  I8a0037ad2845a3fbba9da380a8b8a576['h0786c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c37] =  I8a0037ad2845a3fbba9da380a8b8a576['h0786e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c38] =  I8a0037ad2845a3fbba9da380a8b8a576['h07870] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c39] =  I8a0037ad2845a3fbba9da380a8b8a576['h07872] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c3a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07874] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c3b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07876] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c3c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07878] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c3d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0787a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c3e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0787c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c3f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0787e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c40] =  I8a0037ad2845a3fbba9da380a8b8a576['h07880] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c41] =  I8a0037ad2845a3fbba9da380a8b8a576['h07882] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c42] =  I8a0037ad2845a3fbba9da380a8b8a576['h07884] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c43] =  I8a0037ad2845a3fbba9da380a8b8a576['h07886] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c44] =  I8a0037ad2845a3fbba9da380a8b8a576['h07888] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c45] =  I8a0037ad2845a3fbba9da380a8b8a576['h0788a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c46] =  I8a0037ad2845a3fbba9da380a8b8a576['h0788c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c47] =  I8a0037ad2845a3fbba9da380a8b8a576['h0788e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c48] =  I8a0037ad2845a3fbba9da380a8b8a576['h07890] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c49] =  I8a0037ad2845a3fbba9da380a8b8a576['h07892] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c4a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07894] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c4b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07896] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c4c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07898] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c4d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0789a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c4e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0789c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c4f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0789e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c50] =  I8a0037ad2845a3fbba9da380a8b8a576['h078a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c51] =  I8a0037ad2845a3fbba9da380a8b8a576['h078a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c52] =  I8a0037ad2845a3fbba9da380a8b8a576['h078a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c53] =  I8a0037ad2845a3fbba9da380a8b8a576['h078a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c54] =  I8a0037ad2845a3fbba9da380a8b8a576['h078a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c55] =  I8a0037ad2845a3fbba9da380a8b8a576['h078aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c56] =  I8a0037ad2845a3fbba9da380a8b8a576['h078ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c57] =  I8a0037ad2845a3fbba9da380a8b8a576['h078ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c58] =  I8a0037ad2845a3fbba9da380a8b8a576['h078b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c59] =  I8a0037ad2845a3fbba9da380a8b8a576['h078b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c5a] =  I8a0037ad2845a3fbba9da380a8b8a576['h078b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c5b] =  I8a0037ad2845a3fbba9da380a8b8a576['h078b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c5c] =  I8a0037ad2845a3fbba9da380a8b8a576['h078b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c5d] =  I8a0037ad2845a3fbba9da380a8b8a576['h078ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c5e] =  I8a0037ad2845a3fbba9da380a8b8a576['h078bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c5f] =  I8a0037ad2845a3fbba9da380a8b8a576['h078be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c60] =  I8a0037ad2845a3fbba9da380a8b8a576['h078c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c61] =  I8a0037ad2845a3fbba9da380a8b8a576['h078c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c62] =  I8a0037ad2845a3fbba9da380a8b8a576['h078c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c63] =  I8a0037ad2845a3fbba9da380a8b8a576['h078c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c64] =  I8a0037ad2845a3fbba9da380a8b8a576['h078c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c65] =  I8a0037ad2845a3fbba9da380a8b8a576['h078ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c66] =  I8a0037ad2845a3fbba9da380a8b8a576['h078cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c67] =  I8a0037ad2845a3fbba9da380a8b8a576['h078ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c68] =  I8a0037ad2845a3fbba9da380a8b8a576['h078d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c69] =  I8a0037ad2845a3fbba9da380a8b8a576['h078d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c6a] =  I8a0037ad2845a3fbba9da380a8b8a576['h078d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c6b] =  I8a0037ad2845a3fbba9da380a8b8a576['h078d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c6c] =  I8a0037ad2845a3fbba9da380a8b8a576['h078d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c6d] =  I8a0037ad2845a3fbba9da380a8b8a576['h078da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c6e] =  I8a0037ad2845a3fbba9da380a8b8a576['h078dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c6f] =  I8a0037ad2845a3fbba9da380a8b8a576['h078de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c70] =  I8a0037ad2845a3fbba9da380a8b8a576['h078e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c71] =  I8a0037ad2845a3fbba9da380a8b8a576['h078e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c72] =  I8a0037ad2845a3fbba9da380a8b8a576['h078e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c73] =  I8a0037ad2845a3fbba9da380a8b8a576['h078e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c74] =  I8a0037ad2845a3fbba9da380a8b8a576['h078e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c75] =  I8a0037ad2845a3fbba9da380a8b8a576['h078ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c76] =  I8a0037ad2845a3fbba9da380a8b8a576['h078ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c77] =  I8a0037ad2845a3fbba9da380a8b8a576['h078ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c78] =  I8a0037ad2845a3fbba9da380a8b8a576['h078f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c79] =  I8a0037ad2845a3fbba9da380a8b8a576['h078f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c7a] =  I8a0037ad2845a3fbba9da380a8b8a576['h078f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c7b] =  I8a0037ad2845a3fbba9da380a8b8a576['h078f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c7c] =  I8a0037ad2845a3fbba9da380a8b8a576['h078f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c7d] =  I8a0037ad2845a3fbba9da380a8b8a576['h078fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c7e] =  I8a0037ad2845a3fbba9da380a8b8a576['h078fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c7f] =  I8a0037ad2845a3fbba9da380a8b8a576['h078fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c80] =  I8a0037ad2845a3fbba9da380a8b8a576['h07900] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c81] =  I8a0037ad2845a3fbba9da380a8b8a576['h07902] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c82] =  I8a0037ad2845a3fbba9da380a8b8a576['h07904] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c83] =  I8a0037ad2845a3fbba9da380a8b8a576['h07906] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c84] =  I8a0037ad2845a3fbba9da380a8b8a576['h07908] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c85] =  I8a0037ad2845a3fbba9da380a8b8a576['h0790a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c86] =  I8a0037ad2845a3fbba9da380a8b8a576['h0790c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c87] =  I8a0037ad2845a3fbba9da380a8b8a576['h0790e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c88] =  I8a0037ad2845a3fbba9da380a8b8a576['h07910] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c89] =  I8a0037ad2845a3fbba9da380a8b8a576['h07912] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c8a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07914] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c8b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07916] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c8c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07918] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c8d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0791a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c8e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0791c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c8f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0791e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c90] =  I8a0037ad2845a3fbba9da380a8b8a576['h07920] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c91] =  I8a0037ad2845a3fbba9da380a8b8a576['h07922] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c92] =  I8a0037ad2845a3fbba9da380a8b8a576['h07924] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c93] =  I8a0037ad2845a3fbba9da380a8b8a576['h07926] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c94] =  I8a0037ad2845a3fbba9da380a8b8a576['h07928] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c95] =  I8a0037ad2845a3fbba9da380a8b8a576['h0792a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c96] =  I8a0037ad2845a3fbba9da380a8b8a576['h0792c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c97] =  I8a0037ad2845a3fbba9da380a8b8a576['h0792e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c98] =  I8a0037ad2845a3fbba9da380a8b8a576['h07930] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c99] =  I8a0037ad2845a3fbba9da380a8b8a576['h07932] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c9a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07934] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c9b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07936] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c9c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07938] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c9d] =  I8a0037ad2845a3fbba9da380a8b8a576['h0793a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c9e] =  I8a0037ad2845a3fbba9da380a8b8a576['h0793c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03c9f] =  I8a0037ad2845a3fbba9da380a8b8a576['h0793e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ca0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07940] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ca1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07942] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ca2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07944] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ca3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07946] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ca4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07948] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ca5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0794a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ca6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0794c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ca7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0794e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ca8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07950] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ca9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07952] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03caa] =  I8a0037ad2845a3fbba9da380a8b8a576['h07954] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cab] =  I8a0037ad2845a3fbba9da380a8b8a576['h07956] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cac] =  I8a0037ad2845a3fbba9da380a8b8a576['h07958] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cad] =  I8a0037ad2845a3fbba9da380a8b8a576['h0795a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cae] =  I8a0037ad2845a3fbba9da380a8b8a576['h0795c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03caf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0795e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cb0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07960] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cb1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07962] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cb2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07964] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cb3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07966] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cb4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07968] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cb5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0796a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cb6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0796c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cb7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0796e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cb8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07970] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cb9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07972] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cba] =  I8a0037ad2845a3fbba9da380a8b8a576['h07974] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cbb] =  I8a0037ad2845a3fbba9da380a8b8a576['h07976] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cbc] =  I8a0037ad2845a3fbba9da380a8b8a576['h07978] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cbd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0797a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cbe] =  I8a0037ad2845a3fbba9da380a8b8a576['h0797c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cbf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0797e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cc0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07980] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cc1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07982] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cc2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07984] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cc3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07986] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cc4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07988] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cc5] =  I8a0037ad2845a3fbba9da380a8b8a576['h0798a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cc6] =  I8a0037ad2845a3fbba9da380a8b8a576['h0798c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cc7] =  I8a0037ad2845a3fbba9da380a8b8a576['h0798e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cc8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07990] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cc9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07992] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cca] =  I8a0037ad2845a3fbba9da380a8b8a576['h07994] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ccb] =  I8a0037ad2845a3fbba9da380a8b8a576['h07996] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ccc] =  I8a0037ad2845a3fbba9da380a8b8a576['h07998] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ccd] =  I8a0037ad2845a3fbba9da380a8b8a576['h0799a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cce] =  I8a0037ad2845a3fbba9da380a8b8a576['h0799c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ccf] =  I8a0037ad2845a3fbba9da380a8b8a576['h0799e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cd0] =  I8a0037ad2845a3fbba9da380a8b8a576['h079a0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cd1] =  I8a0037ad2845a3fbba9da380a8b8a576['h079a2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cd2] =  I8a0037ad2845a3fbba9da380a8b8a576['h079a4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cd3] =  I8a0037ad2845a3fbba9da380a8b8a576['h079a6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cd4] =  I8a0037ad2845a3fbba9da380a8b8a576['h079a8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cd5] =  I8a0037ad2845a3fbba9da380a8b8a576['h079aa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cd6] =  I8a0037ad2845a3fbba9da380a8b8a576['h079ac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cd7] =  I8a0037ad2845a3fbba9da380a8b8a576['h079ae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cd8] =  I8a0037ad2845a3fbba9da380a8b8a576['h079b0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cd9] =  I8a0037ad2845a3fbba9da380a8b8a576['h079b2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cda] =  I8a0037ad2845a3fbba9da380a8b8a576['h079b4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cdb] =  I8a0037ad2845a3fbba9da380a8b8a576['h079b6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cdc] =  I8a0037ad2845a3fbba9da380a8b8a576['h079b8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cdd] =  I8a0037ad2845a3fbba9da380a8b8a576['h079ba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cde] =  I8a0037ad2845a3fbba9da380a8b8a576['h079bc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cdf] =  I8a0037ad2845a3fbba9da380a8b8a576['h079be] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ce0] =  I8a0037ad2845a3fbba9da380a8b8a576['h079c0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ce1] =  I8a0037ad2845a3fbba9da380a8b8a576['h079c2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ce2] =  I8a0037ad2845a3fbba9da380a8b8a576['h079c4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ce3] =  I8a0037ad2845a3fbba9da380a8b8a576['h079c6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ce4] =  I8a0037ad2845a3fbba9da380a8b8a576['h079c8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ce5] =  I8a0037ad2845a3fbba9da380a8b8a576['h079ca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ce6] =  I8a0037ad2845a3fbba9da380a8b8a576['h079cc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ce7] =  I8a0037ad2845a3fbba9da380a8b8a576['h079ce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ce8] =  I8a0037ad2845a3fbba9da380a8b8a576['h079d0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ce9] =  I8a0037ad2845a3fbba9da380a8b8a576['h079d2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cea] =  I8a0037ad2845a3fbba9da380a8b8a576['h079d4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ceb] =  I8a0037ad2845a3fbba9da380a8b8a576['h079d6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cec] =  I8a0037ad2845a3fbba9da380a8b8a576['h079d8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ced] =  I8a0037ad2845a3fbba9da380a8b8a576['h079da] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cee] =  I8a0037ad2845a3fbba9da380a8b8a576['h079dc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cef] =  I8a0037ad2845a3fbba9da380a8b8a576['h079de] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cf0] =  I8a0037ad2845a3fbba9da380a8b8a576['h079e0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cf1] =  I8a0037ad2845a3fbba9da380a8b8a576['h079e2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cf2] =  I8a0037ad2845a3fbba9da380a8b8a576['h079e4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cf3] =  I8a0037ad2845a3fbba9da380a8b8a576['h079e6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cf4] =  I8a0037ad2845a3fbba9da380a8b8a576['h079e8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cf5] =  I8a0037ad2845a3fbba9da380a8b8a576['h079ea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cf6] =  I8a0037ad2845a3fbba9da380a8b8a576['h079ec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cf7] =  I8a0037ad2845a3fbba9da380a8b8a576['h079ee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cf8] =  I8a0037ad2845a3fbba9da380a8b8a576['h079f0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cf9] =  I8a0037ad2845a3fbba9da380a8b8a576['h079f2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cfa] =  I8a0037ad2845a3fbba9da380a8b8a576['h079f4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cfb] =  I8a0037ad2845a3fbba9da380a8b8a576['h079f6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cfc] =  I8a0037ad2845a3fbba9da380a8b8a576['h079f8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cfd] =  I8a0037ad2845a3fbba9da380a8b8a576['h079fa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cfe] =  I8a0037ad2845a3fbba9da380a8b8a576['h079fc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03cff] =  I8a0037ad2845a3fbba9da380a8b8a576['h079fe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d00] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d01] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d02] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d03] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d04] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d05] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d06] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d07] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d08] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d09] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d0a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d0b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d0c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d0d] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d0e] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d0f] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d10] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d11] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d12] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d13] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d14] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d15] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d16] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d17] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d18] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d19] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d1a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d1b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d1c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d1d] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d1e] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d1f] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d20] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d21] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d22] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d23] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d24] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d25] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d26] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d27] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d28] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d29] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d2a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d2b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d2c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d2d] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d2e] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d2f] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d30] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d31] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d32] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d33] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d34] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d35] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d36] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d37] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d38] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d39] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d3a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d3b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d3c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d3d] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d3e] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d3f] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d40] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d41] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d42] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d43] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d44] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d45] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d46] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d47] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d48] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d49] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d4a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d4b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d4c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d4d] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d4e] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d4f] =  I8a0037ad2845a3fbba9da380a8b8a576['h07a9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d50] =  I8a0037ad2845a3fbba9da380a8b8a576['h07aa0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d51] =  I8a0037ad2845a3fbba9da380a8b8a576['h07aa2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d52] =  I8a0037ad2845a3fbba9da380a8b8a576['h07aa4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d53] =  I8a0037ad2845a3fbba9da380a8b8a576['h07aa6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d54] =  I8a0037ad2845a3fbba9da380a8b8a576['h07aa8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d55] =  I8a0037ad2845a3fbba9da380a8b8a576['h07aaa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d56] =  I8a0037ad2845a3fbba9da380a8b8a576['h07aac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d57] =  I8a0037ad2845a3fbba9da380a8b8a576['h07aae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d58] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ab0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d59] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ab2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d5a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ab4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d5b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ab6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d5c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ab8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d5d] =  I8a0037ad2845a3fbba9da380a8b8a576['h07aba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d5e] =  I8a0037ad2845a3fbba9da380a8b8a576['h07abc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d5f] =  I8a0037ad2845a3fbba9da380a8b8a576['h07abe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d60] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ac0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d61] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ac2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d62] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ac4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d63] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ac6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d64] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ac8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d65] =  I8a0037ad2845a3fbba9da380a8b8a576['h07aca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d66] =  I8a0037ad2845a3fbba9da380a8b8a576['h07acc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d67] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ace] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d68] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ad0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d69] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ad2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d6a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ad4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d6b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ad6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d6c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ad8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d6d] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ada] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d6e] =  I8a0037ad2845a3fbba9da380a8b8a576['h07adc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d6f] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ade] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d70] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ae0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d71] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ae2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d72] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ae4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d73] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ae6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d74] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ae8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d75] =  I8a0037ad2845a3fbba9da380a8b8a576['h07aea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d76] =  I8a0037ad2845a3fbba9da380a8b8a576['h07aec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d77] =  I8a0037ad2845a3fbba9da380a8b8a576['h07aee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d78] =  I8a0037ad2845a3fbba9da380a8b8a576['h07af0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d79] =  I8a0037ad2845a3fbba9da380a8b8a576['h07af2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d7a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07af4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d7b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07af6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d7c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07af8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d7d] =  I8a0037ad2845a3fbba9da380a8b8a576['h07afa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d7e] =  I8a0037ad2845a3fbba9da380a8b8a576['h07afc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d7f] =  I8a0037ad2845a3fbba9da380a8b8a576['h07afe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d80] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d81] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d82] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d83] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d84] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d85] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d86] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d87] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d88] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d89] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d8a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d8b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d8c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d8d] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d8e] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d8f] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d90] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d91] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d92] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d93] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d94] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d95] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d96] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d97] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d98] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d99] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d9a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d9b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d9c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d9d] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d9e] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03d9f] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03da0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03da1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03da2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03da3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03da4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03da5] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03da6] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03da7] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03da8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03da9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03daa] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dab] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dac] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dad] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dae] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03daf] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03db0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03db1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03db2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03db3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03db4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03db5] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03db6] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03db7] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03db8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03db9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dba] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dbb] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dbc] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dbd] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dbe] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dbf] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dc0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dc1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dc2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dc3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dc4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dc5] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dc6] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dc7] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dc8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dc9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dca] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dcb] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dcc] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dcd] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dce] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dcf] =  I8a0037ad2845a3fbba9da380a8b8a576['h07b9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dd0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ba0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dd1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ba2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dd2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ba4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dd3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ba6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dd4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ba8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dd5] =  I8a0037ad2845a3fbba9da380a8b8a576['h07baa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dd6] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dd7] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dd8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dd9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dda] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ddb] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ddc] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ddd] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dde] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ddf] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03de0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03de1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03de2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03de3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03de4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03de5] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03de6] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bcc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03de7] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03de8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03de9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dea] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03deb] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dec] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ded] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dee] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bdc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03def] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03df0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07be0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03df1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07be2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03df2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07be4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03df3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07be6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03df4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07be8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03df5] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03df6] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03df7] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03df8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bf0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03df9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bf2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dfa] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bf4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dfb] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bf6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dfc] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bf8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dfd] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bfa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dfe] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bfc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03dff] =  I8a0037ad2845a3fbba9da380a8b8a576['h07bfe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e00] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e01] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e02] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e03] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e04] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e05] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e06] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e07] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e08] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e09] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e0a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e0b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e0c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e0d] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e0e] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e0f] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e10] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e11] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e12] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e13] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e14] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e15] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e16] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e17] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e18] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e19] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e1a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e1b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e1c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e1d] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e1e] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e1f] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e20] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e21] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e22] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e23] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e24] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e25] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e26] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e27] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e28] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e29] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e2a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e2b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e2c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e2d] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e2e] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e2f] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e30] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e31] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e32] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e33] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e34] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e35] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e36] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e37] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e38] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e39] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e3a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e3b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e3c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e3d] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e3e] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e3f] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e40] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e41] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e42] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e43] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e44] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e45] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e46] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e47] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e48] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e49] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e4a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e4b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e4c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e4d] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e4e] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e4f] =  I8a0037ad2845a3fbba9da380a8b8a576['h07c9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e50] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ca0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e51] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ca2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e52] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ca4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e53] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ca6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e54] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ca8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e55] =  I8a0037ad2845a3fbba9da380a8b8a576['h07caa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e56] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e57] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e58] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e59] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e5a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e5b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e5c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e5d] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e5e] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e5f] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e60] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e61] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e62] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e63] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e64] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e65] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e66] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ccc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e67] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e68] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e69] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e6a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e6b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e6c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e6d] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e6e] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cdc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e6f] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e70] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ce0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e71] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ce2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e72] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ce4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e73] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ce6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e74] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ce8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e75] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e76] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e77] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e78] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cf0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e79] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cf2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e7a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cf4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e7b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cf6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e7c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cf8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e7d] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cfa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e7e] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cfc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e7f] =  I8a0037ad2845a3fbba9da380a8b8a576['h07cfe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e80] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e81] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e82] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e83] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e84] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e85] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e86] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e87] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e88] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e89] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e8a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e8b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e8c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e8d] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e8e] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e8f] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e90] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e91] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e92] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e93] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e94] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e95] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e96] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e97] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e98] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e99] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e9a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e9b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e9c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e9d] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e9e] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03e9f] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ea0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ea1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ea2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ea3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ea4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ea5] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ea6] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ea7] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ea8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ea9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03eaa] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03eab] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03eac] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ead] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03eae] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03eaf] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03eb0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03eb1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03eb2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03eb3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03eb4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03eb5] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03eb6] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03eb7] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03eb8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03eb9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03eba] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ebb] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ebc] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ebd] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ebe] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ebf] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ec0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ec1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ec2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ec3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ec4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ec5] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ec6] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ec7] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ec8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ec9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03eca] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ecb] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ecc] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ecd] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ece] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ecf] =  I8a0037ad2845a3fbba9da380a8b8a576['h07d9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ed0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07da0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ed1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07da2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ed2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07da4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ed3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07da6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ed4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07da8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ed5] =  I8a0037ad2845a3fbba9da380a8b8a576['h07daa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ed6] =  I8a0037ad2845a3fbba9da380a8b8a576['h07dac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ed7] =  I8a0037ad2845a3fbba9da380a8b8a576['h07dae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ed8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07db0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ed9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07db2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03eda] =  I8a0037ad2845a3fbba9da380a8b8a576['h07db4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03edb] =  I8a0037ad2845a3fbba9da380a8b8a576['h07db6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03edc] =  I8a0037ad2845a3fbba9da380a8b8a576['h07db8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03edd] =  I8a0037ad2845a3fbba9da380a8b8a576['h07dba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ede] =  I8a0037ad2845a3fbba9da380a8b8a576['h07dbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03edf] =  I8a0037ad2845a3fbba9da380a8b8a576['h07dbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ee0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07dc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ee1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07dc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ee2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07dc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ee3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07dc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ee4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07dc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ee5] =  I8a0037ad2845a3fbba9da380a8b8a576['h07dca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ee6] =  I8a0037ad2845a3fbba9da380a8b8a576['h07dcc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ee7] =  I8a0037ad2845a3fbba9da380a8b8a576['h07dce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ee8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07dd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ee9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07dd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03eea] =  I8a0037ad2845a3fbba9da380a8b8a576['h07dd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03eeb] =  I8a0037ad2845a3fbba9da380a8b8a576['h07dd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03eec] =  I8a0037ad2845a3fbba9da380a8b8a576['h07dd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03eed] =  I8a0037ad2845a3fbba9da380a8b8a576['h07dda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03eee] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ddc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03eef] =  I8a0037ad2845a3fbba9da380a8b8a576['h07dde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ef0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07de0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ef1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07de2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ef2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07de4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ef3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07de6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ef4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07de8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ef5] =  I8a0037ad2845a3fbba9da380a8b8a576['h07dea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ef6] =  I8a0037ad2845a3fbba9da380a8b8a576['h07dec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ef7] =  I8a0037ad2845a3fbba9da380a8b8a576['h07dee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ef8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07df0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ef9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07df2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03efa] =  I8a0037ad2845a3fbba9da380a8b8a576['h07df4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03efb] =  I8a0037ad2845a3fbba9da380a8b8a576['h07df6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03efc] =  I8a0037ad2845a3fbba9da380a8b8a576['h07df8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03efd] =  I8a0037ad2845a3fbba9da380a8b8a576['h07dfa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03efe] =  I8a0037ad2845a3fbba9da380a8b8a576['h07dfc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03eff] =  I8a0037ad2845a3fbba9da380a8b8a576['h07dfe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f00] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f01] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f02] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f03] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f04] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f05] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f06] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f07] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f08] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f09] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f0a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f0b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f0c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f0d] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f0e] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f0f] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f10] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f11] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f12] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f13] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f14] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f15] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f16] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f17] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f18] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f19] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f1a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f1b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f1c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f1d] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f1e] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f1f] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f20] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f21] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f22] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f23] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f24] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f25] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f26] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f27] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f28] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f29] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f2a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f2b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f2c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f2d] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f2e] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f2f] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f30] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f31] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f32] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f33] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f34] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f35] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f36] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f37] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f38] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f39] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f3a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f3b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f3c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f3d] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f3e] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f3f] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f40] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f41] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f42] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f43] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f44] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f45] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f46] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f47] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f48] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f49] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f4a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f4b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f4c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f4d] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f4e] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f4f] =  I8a0037ad2845a3fbba9da380a8b8a576['h07e9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f50] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ea0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f51] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ea2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f52] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ea4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f53] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ea6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f54] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ea8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f55] =  I8a0037ad2845a3fbba9da380a8b8a576['h07eaa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f56] =  I8a0037ad2845a3fbba9da380a8b8a576['h07eac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f57] =  I8a0037ad2845a3fbba9da380a8b8a576['h07eae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f58] =  I8a0037ad2845a3fbba9da380a8b8a576['h07eb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f59] =  I8a0037ad2845a3fbba9da380a8b8a576['h07eb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f5a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07eb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f5b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07eb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f5c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07eb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f5d] =  I8a0037ad2845a3fbba9da380a8b8a576['h07eba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f5e] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ebc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f5f] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ebe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f60] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ec0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f61] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ec2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f62] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ec4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f63] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ec6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f64] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ec8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f65] =  I8a0037ad2845a3fbba9da380a8b8a576['h07eca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f66] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ecc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f67] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ece] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f68] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ed0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f69] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ed2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f6a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ed4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f6b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ed6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f6c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ed8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f6d] =  I8a0037ad2845a3fbba9da380a8b8a576['h07eda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f6e] =  I8a0037ad2845a3fbba9da380a8b8a576['h07edc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f6f] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ede] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f70] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ee0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f71] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ee2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f72] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ee4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f73] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ee6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f74] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ee8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f75] =  I8a0037ad2845a3fbba9da380a8b8a576['h07eea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f76] =  I8a0037ad2845a3fbba9da380a8b8a576['h07eec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f77] =  I8a0037ad2845a3fbba9da380a8b8a576['h07eee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f78] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ef0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f79] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ef2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f7a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ef4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f7b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ef6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f7c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ef8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f7d] =  I8a0037ad2845a3fbba9da380a8b8a576['h07efa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f7e] =  I8a0037ad2845a3fbba9da380a8b8a576['h07efc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f7f] =  I8a0037ad2845a3fbba9da380a8b8a576['h07efe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f80] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f00] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f81] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f02] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f82] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f04] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f83] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f06] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f84] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f08] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f85] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f0a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f86] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f0c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f87] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f0e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f88] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f10] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f89] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f12] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f8a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f14] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f8b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f16] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f8c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f18] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f8d] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f1a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f8e] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f1c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f8f] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f1e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f90] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f20] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f91] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f22] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f92] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f24] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f93] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f26] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f94] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f28] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f95] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f2a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f96] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f2c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f97] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f2e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f98] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f30] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f99] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f32] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f9a] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f34] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f9b] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f36] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f9c] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f38] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f9d] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f3a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f9e] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f3c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03f9f] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f3e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fa0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f40] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fa1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f42] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fa2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f44] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fa3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f46] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fa4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f48] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fa5] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f4a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fa6] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f4c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fa7] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f4e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fa8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f50] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fa9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f52] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03faa] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f54] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fab] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f56] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fac] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f58] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fad] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f5a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fae] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f5c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03faf] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f5e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fb0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f60] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fb1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f62] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fb2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f64] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fb3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f66] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fb4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f68] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fb5] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f6a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fb6] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f6c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fb7] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f6e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fb8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f70] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fb9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f72] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fba] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f74] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fbb] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f76] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fbc] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f78] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fbd] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f7a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fbe] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f7c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fbf] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f7e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fc0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f80] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fc1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f82] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fc2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f84] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fc3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f86] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fc4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f88] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fc5] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f8a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fc6] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f8c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fc7] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f8e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fc8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f90] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fc9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f92] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fca] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f94] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fcb] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f96] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fcc] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f98] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fcd] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f9a] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fce] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f9c] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fcf] =  I8a0037ad2845a3fbba9da380a8b8a576['h07f9e] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fd0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fa0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fd1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fa2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fd2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fa4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fd3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fa6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fd4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fa8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fd5] =  I8a0037ad2845a3fbba9da380a8b8a576['h07faa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fd6] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fac] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fd7] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fae] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fd8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fb0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fd9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fb2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fda] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fb4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fdb] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fb6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fdc] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fb8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fdd] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fba] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fde] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fbc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fdf] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fbe] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fe0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fc0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fe1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fc2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fe2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fc4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fe3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fc6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fe4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fc8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fe5] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fca] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fe6] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fcc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fe7] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fce] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fe8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fd0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fe9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fd2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fea] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fd4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03feb] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fd6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fec] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fd8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fed] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fda] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fee] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fdc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fef] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fde] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ff0] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fe0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ff1] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fe2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ff2] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fe4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ff3] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fe6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ff4] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fe8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ff5] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fea] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ff6] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fec] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ff7] =  I8a0037ad2845a3fbba9da380a8b8a576['h07fee] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ff8] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ff0] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ff9] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ff2] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ffa] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ff4] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ffb] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ff6] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ffc] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ff8] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ffd] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ffa] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03ffe] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ffc] ;
//end
//always_comb begin // 
               I0310077d53ae4ed9904df42e3f81c634['h03fff] =  I8a0037ad2845a3fbba9da380a8b8a576['h07ffe] ;
//end
