 parameter fgallag_WDTH =  20 ;
 reg  [fgallag_WDTH -1 :0] fgallag_sel ;
 reg  [$clog2('h7000+1)-1:0] I7ffcaba1b7d64b619b19a68a22aa495d ;
