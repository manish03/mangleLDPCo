//`include "GF2_LDPC_fgallag_0x00005_assign_inc.sv"
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00000] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00000] : //%
                       Ifd35529b44c957737bf422127283c08e['h00001] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00001] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00002] : //%
                       Ifd35529b44c957737bf422127283c08e['h00003] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00002] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00004] : //%
                       Ifd35529b44c957737bf422127283c08e['h00005] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00003] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00006] : //%
                       Ifd35529b44c957737bf422127283c08e['h00007] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00004] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00008] : //%
                       Ifd35529b44c957737bf422127283c08e['h00009] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00005] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0000a] : //%
                       Ifd35529b44c957737bf422127283c08e['h0000b] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00006] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0000c] : //%
                       Ifd35529b44c957737bf422127283c08e['h0000d] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00007] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0000e] : //%
                       Ifd35529b44c957737bf422127283c08e['h0000f] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00008] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00010] : //%
                       Ifd35529b44c957737bf422127283c08e['h00011] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00009] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00012] : //%
                       Ifd35529b44c957737bf422127283c08e['h00013] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0000a] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00014] : //%
                       Ifd35529b44c957737bf422127283c08e['h00015] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0000b] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00016] : //%
                       Ifd35529b44c957737bf422127283c08e['h00017] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0000c] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00018] : //%
                       Ifd35529b44c957737bf422127283c08e['h00019] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0000d] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0001a] : //%
                       Ifd35529b44c957737bf422127283c08e['h0001b] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0000e] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0001c] : //%
                       Ifd35529b44c957737bf422127283c08e['h0001d] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0000f] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0001e] : //%
                       Ifd35529b44c957737bf422127283c08e['h0001f] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00010] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00020] : //%
                       Ifd35529b44c957737bf422127283c08e['h00021] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00011] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00022] : //%
                       Ifd35529b44c957737bf422127283c08e['h00023] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00012] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00024] : //%
                       Ifd35529b44c957737bf422127283c08e['h00025] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00013] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00026] : //%
                       Ifd35529b44c957737bf422127283c08e['h00027] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00014] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00028] : //%
                       Ifd35529b44c957737bf422127283c08e['h00029] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00015] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0002a] : //%
                       Ifd35529b44c957737bf422127283c08e['h0002b] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00016] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0002c] : //%
                       Ifd35529b44c957737bf422127283c08e['h0002d] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00017] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0002e] : //%
                       Ifd35529b44c957737bf422127283c08e['h0002f] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00018] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00030] : //%
                       Ifd35529b44c957737bf422127283c08e['h00031] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00019] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00032] : //%
                       Ifd35529b44c957737bf422127283c08e['h00033] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0001a] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00034] : //%
                       Ifd35529b44c957737bf422127283c08e['h00035] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0001b] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00036] : //%
                       Ifd35529b44c957737bf422127283c08e['h00037] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0001c] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00038] : //%
                       Ifd35529b44c957737bf422127283c08e['h00039] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0001d] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0003a] : //%
                       Ifd35529b44c957737bf422127283c08e['h0003b] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0001e] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0003c] : //%
                       Ifd35529b44c957737bf422127283c08e['h0003d] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0001f] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0003e] : //%
                       Ifd35529b44c957737bf422127283c08e['h0003f] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00020] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00040] : //%
                       Ifd35529b44c957737bf422127283c08e['h00041] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00021] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00042] : //%
                       Ifd35529b44c957737bf422127283c08e['h00043] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00022] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00044] : //%
                       Ifd35529b44c957737bf422127283c08e['h00045] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00023] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00046] : //%
                       Ifd35529b44c957737bf422127283c08e['h00047] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00024] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00048] : //%
                       Ifd35529b44c957737bf422127283c08e['h00049] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00025] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0004a] : //%
                       Ifd35529b44c957737bf422127283c08e['h0004b] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00026] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0004c] : //%
                       Ifd35529b44c957737bf422127283c08e['h0004d] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00027] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0004e] : //%
                       Ifd35529b44c957737bf422127283c08e['h0004f] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00028] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00050] : //%
                       Ifd35529b44c957737bf422127283c08e['h00051] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00029] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00052] : //%
                       Ifd35529b44c957737bf422127283c08e['h00053] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0002a] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00054] : //%
                       Ifd35529b44c957737bf422127283c08e['h00055] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0002b] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00056] : //%
                       Ifd35529b44c957737bf422127283c08e['h00057] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0002c] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00058] : //%
                       Ifd35529b44c957737bf422127283c08e['h00059] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0002d] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0005a] : //%
                       Ifd35529b44c957737bf422127283c08e['h0005b] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0002e] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0005c] : //%
                       Ifd35529b44c957737bf422127283c08e['h0005d] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0002f] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0005e] : //%
                       Ifd35529b44c957737bf422127283c08e['h0005f] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00030] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00060] : //%
                       Ifd35529b44c957737bf422127283c08e['h00061] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00031] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00062] : //%
                       Ifd35529b44c957737bf422127283c08e['h00063] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00032] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00064] : //%
                       Ifd35529b44c957737bf422127283c08e['h00065] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00033] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00066] : //%
                       Ifd35529b44c957737bf422127283c08e['h00067] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00034] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00068] : //%
                       Ifd35529b44c957737bf422127283c08e['h00069] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00035] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0006a] : //%
                       Ifd35529b44c957737bf422127283c08e['h0006b] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00036] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0006c] : //%
                       Ifd35529b44c957737bf422127283c08e['h0006d] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00037] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0006e] : //%
                       Ifd35529b44c957737bf422127283c08e['h0006f] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00038] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00070] : //%
                       Ifd35529b44c957737bf422127283c08e['h00071] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00039] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00072] : //%
                       Ifd35529b44c957737bf422127283c08e['h00073] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0003a] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00074] : //%
                       Ifd35529b44c957737bf422127283c08e['h00075] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0003b] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00076] : //%
                       Ifd35529b44c957737bf422127283c08e['h00077] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0003c] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00078] : //%
                       Ifd35529b44c957737bf422127283c08e['h00079] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0003d] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0007a] : //%
                       Ifd35529b44c957737bf422127283c08e['h0007b] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0003e] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0007c] : //%
                       Ifd35529b44c957737bf422127283c08e['h0007d] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0003f] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0007e] : //%
                       Ifd35529b44c957737bf422127283c08e['h0007f] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00040] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00080] : //%
                       Ifd35529b44c957737bf422127283c08e['h00081] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00041] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00082] : //%
                       Ifd35529b44c957737bf422127283c08e['h00083] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00042] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00084] : //%
                       Ifd35529b44c957737bf422127283c08e['h00085] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00043] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00086] : //%
                       Ifd35529b44c957737bf422127283c08e['h00087] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00044] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00088] : //%
                       Ifd35529b44c957737bf422127283c08e['h00089] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00045] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0008a] : //%
                       Ifd35529b44c957737bf422127283c08e['h0008b] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00046] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0008c] : //%
                       Ifd35529b44c957737bf422127283c08e['h0008d] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00047] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0008e] : //%
                       Ifd35529b44c957737bf422127283c08e['h0008f] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00048] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00090] : //%
                       Ifd35529b44c957737bf422127283c08e['h00091] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00049] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00092] : //%
                       Ifd35529b44c957737bf422127283c08e['h00093] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0004a] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00094] : //%
                       Ifd35529b44c957737bf422127283c08e['h00095] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0004b] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00096] : //%
                       Ifd35529b44c957737bf422127283c08e['h00097] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0004c] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00098] : //%
                       Ifd35529b44c957737bf422127283c08e['h00099] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0004d] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0009a] : //%
                       Ifd35529b44c957737bf422127283c08e['h0009b] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0004e] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0009c] : //%
                       Ifd35529b44c957737bf422127283c08e['h0009d] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0004f] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0009e] : //%
                       Ifd35529b44c957737bf422127283c08e['h0009f] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00050] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000a0] : //%
                       Ifd35529b44c957737bf422127283c08e['h000a1] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00051] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000a2] : //%
                       Ifd35529b44c957737bf422127283c08e['h000a3] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00052] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000a4] : //%
                       Ifd35529b44c957737bf422127283c08e['h000a5] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00053] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000a6] : //%
                       Ifd35529b44c957737bf422127283c08e['h000a7] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00054] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000a8] : //%
                       Ifd35529b44c957737bf422127283c08e['h000a9] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00055] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000aa] : //%
                       Ifd35529b44c957737bf422127283c08e['h000ab] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00056] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000ac] : //%
                       Ifd35529b44c957737bf422127283c08e['h000ad] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00057] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000ae] : //%
                       Ifd35529b44c957737bf422127283c08e['h000af] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00058] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000b0] : //%
                       Ifd35529b44c957737bf422127283c08e['h000b1] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00059] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000b2] : //%
                       Ifd35529b44c957737bf422127283c08e['h000b3] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0005a] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000b4] : //%
                       Ifd35529b44c957737bf422127283c08e['h000b5] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0005b] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000b6] : //%
                       Ifd35529b44c957737bf422127283c08e['h000b7] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0005c] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000b8] : //%
                       Ifd35529b44c957737bf422127283c08e['h000b9] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0005d] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000ba] : //%
                       Ifd35529b44c957737bf422127283c08e['h000bb] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0005e] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000bc] : //%
                       Ifd35529b44c957737bf422127283c08e['h000bd] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0005f] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000be] : //%
                       Ifd35529b44c957737bf422127283c08e['h000bf] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00060] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000c0] : //%
                       Ifd35529b44c957737bf422127283c08e['h000c1] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00061] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000c2] : //%
                       Ifd35529b44c957737bf422127283c08e['h000c3] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00062] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000c4] : //%
                       Ifd35529b44c957737bf422127283c08e['h000c5] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00063] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000c6] : //%
                       Ifd35529b44c957737bf422127283c08e['h000c7] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00064] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000c8] : //%
                       Ifd35529b44c957737bf422127283c08e['h000c9] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00065] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000ca] : //%
                       Ifd35529b44c957737bf422127283c08e['h000cb] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00066] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000cc] : //%
                       Ifd35529b44c957737bf422127283c08e['h000cd] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00067] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000ce] : //%
                       Ifd35529b44c957737bf422127283c08e['h000cf] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00068] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000d0] : //%
                       Ifd35529b44c957737bf422127283c08e['h000d1] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00069] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000d2] : //%
                       Ifd35529b44c957737bf422127283c08e['h000d3] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0006a] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000d4] : //%
                       Ifd35529b44c957737bf422127283c08e['h000d5] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0006b] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000d6] : //%
                       Ifd35529b44c957737bf422127283c08e['h000d7] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0006c] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000d8] : //%
                       Ifd35529b44c957737bf422127283c08e['h000d9] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0006d] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000da] : //%
                       Ifd35529b44c957737bf422127283c08e['h000db] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0006e] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000dc] : //%
                       Ifd35529b44c957737bf422127283c08e['h000dd] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0006f] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000de] : //%
                       Ifd35529b44c957737bf422127283c08e['h000df] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00070] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000e0] : //%
                       Ifd35529b44c957737bf422127283c08e['h000e1] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00071] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000e2] : //%
                       Ifd35529b44c957737bf422127283c08e['h000e3] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00072] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000e4] : //%
                       Ifd35529b44c957737bf422127283c08e['h000e5] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00073] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000e6] : //%
                       Ifd35529b44c957737bf422127283c08e['h000e7] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00074] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000e8] : //%
                       Ifd35529b44c957737bf422127283c08e['h000e9] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00075] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000ea] : //%
                       Ifd35529b44c957737bf422127283c08e['h000eb] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00076] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000ec] : //%
                       Ifd35529b44c957737bf422127283c08e['h000ed] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00077] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000ee] : //%
                       Ifd35529b44c957737bf422127283c08e['h000ef] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00078] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000f0] : //%
                       Ifd35529b44c957737bf422127283c08e['h000f1] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00079] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000f2] : //%
                       Ifd35529b44c957737bf422127283c08e['h000f3] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0007a] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000f4] : //%
                       Ifd35529b44c957737bf422127283c08e['h000f5] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0007b] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000f6] : //%
                       Ifd35529b44c957737bf422127283c08e['h000f7] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0007c] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000f8] : //%
                       Ifd35529b44c957737bf422127283c08e['h000f9] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0007d] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000fa] : //%
                       Ifd35529b44c957737bf422127283c08e['h000fb] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0007e] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000fc] : //%
                       Ifd35529b44c957737bf422127283c08e['h000fd] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0007f] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h000fe] : //%
                       Ifd35529b44c957737bf422127283c08e['h000ff] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00080] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00100] : //%
                       Ifd35529b44c957737bf422127283c08e['h00101] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00081] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00102] : //%
                       Ifd35529b44c957737bf422127283c08e['h00103] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00082] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00104] : //%
                       Ifd35529b44c957737bf422127283c08e['h00105] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00083] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00106] : //%
                       Ifd35529b44c957737bf422127283c08e['h00107] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00084] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00108] : //%
                       Ifd35529b44c957737bf422127283c08e['h00109] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00085] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0010a] : //%
                       Ifd35529b44c957737bf422127283c08e['h0010b] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00086] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0010c] : //%
                       Ifd35529b44c957737bf422127283c08e['h0010d] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00087] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0010e] : //%
                       Ifd35529b44c957737bf422127283c08e['h0010f] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00088] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00110] : //%
                       Ifd35529b44c957737bf422127283c08e['h00111] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00089] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00112] : //%
                       Ifd35529b44c957737bf422127283c08e['h00113] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0008a] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00114] : //%
                       Ifd35529b44c957737bf422127283c08e['h00115] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0008b] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00116] : //%
                       Ifd35529b44c957737bf422127283c08e['h00117] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0008c] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00118] : //%
                       Ifd35529b44c957737bf422127283c08e['h00119] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0008d] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0011a] : //%
                       Ifd35529b44c957737bf422127283c08e['h0011b] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0008e] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0011c] : //%
                       Ifd35529b44c957737bf422127283c08e['h0011d] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0008f] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0011e] : //%
                       Ifd35529b44c957737bf422127283c08e['h0011f] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00090] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00120] : //%
                       Ifd35529b44c957737bf422127283c08e['h00121] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00091] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00122] : //%
                       Ifd35529b44c957737bf422127283c08e['h00123] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00092] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00124] : //%
                       Ifd35529b44c957737bf422127283c08e['h00125] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00093] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00126] : //%
                       Ifd35529b44c957737bf422127283c08e['h00127] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00094] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00128] : //%
                       Ifd35529b44c957737bf422127283c08e['h00129] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00095] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0012a] : //%
                       Ifd35529b44c957737bf422127283c08e['h0012b] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00096] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0012c] : //%
                       Ifd35529b44c957737bf422127283c08e['h0012d] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00097] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0012e] : //%
                       Ifd35529b44c957737bf422127283c08e['h0012f] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00098] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00130] : //%
                       Ifd35529b44c957737bf422127283c08e['h00131] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00099] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00132] : //%
                       Ifd35529b44c957737bf422127283c08e['h00133] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0009a] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00134] : //%
                       Ifd35529b44c957737bf422127283c08e['h00135] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0009b] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00136] : //%
                       Ifd35529b44c957737bf422127283c08e['h00137] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0009c] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00138] : //%
                       Ifd35529b44c957737bf422127283c08e['h00139] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0009d] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0013a] : //%
                       Ifd35529b44c957737bf422127283c08e['h0013b] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h0009e] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0013c] : //%
                       Ifd35529b44c957737bf422127283c08e['h0013d] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0009f] =  Ifd35529b44c957737bf422127283c08e['h0013e] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h000a0] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00140] : //%
                       Ifd35529b44c957737bf422127283c08e['h00141] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h000a1] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00142] : //%
                       Ifd35529b44c957737bf422127283c08e['h00143] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h000a2] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00144] : //%
                       Ifd35529b44c957737bf422127283c08e['h00145] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h000a3] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00146] : //%
                       Ifd35529b44c957737bf422127283c08e['h00147] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000a4] =  Ifd35529b44c957737bf422127283c08e['h00148] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h000a5] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0014a] : //%
                       Ifd35529b44c957737bf422127283c08e['h0014b] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h000a6] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0014c] : //%
                       Ifd35529b44c957737bf422127283c08e['h0014d] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000a7] =  Ifd35529b44c957737bf422127283c08e['h0014e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000a8] =  Ifd35529b44c957737bf422127283c08e['h00150] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h000a9] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00152] : //%
                       Ifd35529b44c957737bf422127283c08e['h00153] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000aa] =  Ifd35529b44c957737bf422127283c08e['h00154] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h000ab] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00156] : //%
                       Ifd35529b44c957737bf422127283c08e['h00157] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h000ac] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00158] : //%
                       Ifd35529b44c957737bf422127283c08e['h00159] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000ad] =  Ifd35529b44c957737bf422127283c08e['h0015a] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h000ae] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0015c] : //%
                       Ifd35529b44c957737bf422127283c08e['h0015d] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000af] =  Ifd35529b44c957737bf422127283c08e['h0015e] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h000b0] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00160] : //%
                       Ifd35529b44c957737bf422127283c08e['h00161] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000b1] =  Ifd35529b44c957737bf422127283c08e['h00162] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h000b2] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00164] : //%
                       Ifd35529b44c957737bf422127283c08e['h00165] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000b3] =  Ifd35529b44c957737bf422127283c08e['h00166] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h000b4] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00168] : //%
                       Ifd35529b44c957737bf422127283c08e['h00169] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000b5] =  Ifd35529b44c957737bf422127283c08e['h0016a] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h000b6] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0016c] : //%
                       Ifd35529b44c957737bf422127283c08e['h0016d] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000b7] =  Ifd35529b44c957737bf422127283c08e['h0016e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000b8] =  Ifd35529b44c957737bf422127283c08e['h00170] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h000b9] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00172] : //%
                       Ifd35529b44c957737bf422127283c08e['h00173] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000ba] =  Ifd35529b44c957737bf422127283c08e['h00174] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000bb] =  Ifd35529b44c957737bf422127283c08e['h00176] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h000bc] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00178] : //%
                       Ifd35529b44c957737bf422127283c08e['h00179] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000bd] =  Ifd35529b44c957737bf422127283c08e['h0017a] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h000be] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0017c] : //%
                       Ifd35529b44c957737bf422127283c08e['h0017d] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000bf] =  Ifd35529b44c957737bf422127283c08e['h0017e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000c0] =  Ifd35529b44c957737bf422127283c08e['h00180] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000c1] =  Ifd35529b44c957737bf422127283c08e['h00182] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h000c2] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00184] : //%
                       Ifd35529b44c957737bf422127283c08e['h00185] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000c3] =  Ifd35529b44c957737bf422127283c08e['h00186] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000c4] =  Ifd35529b44c957737bf422127283c08e['h00188] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h000c5] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0018a] : //%
                       Ifd35529b44c957737bf422127283c08e['h0018b] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000c6] =  Ifd35529b44c957737bf422127283c08e['h0018c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000c7] =  Ifd35529b44c957737bf422127283c08e['h0018e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000c8] =  Ifd35529b44c957737bf422127283c08e['h00190] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h000c9] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00192] : //%
                       Ifd35529b44c957737bf422127283c08e['h00193] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000ca] =  Ifd35529b44c957737bf422127283c08e['h00194] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000cb] =  Ifd35529b44c957737bf422127283c08e['h00196] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000cc] =  Ifd35529b44c957737bf422127283c08e['h00198] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000cd] =  Ifd35529b44c957737bf422127283c08e['h0019a] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h000ce] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h0019c] : //%
                       Ifd35529b44c957737bf422127283c08e['h0019d] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000cf] =  Ifd35529b44c957737bf422127283c08e['h0019e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000d0] =  Ifd35529b44c957737bf422127283c08e['h001a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000d1] =  Ifd35529b44c957737bf422127283c08e['h001a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000d2] =  Ifd35529b44c957737bf422127283c08e['h001a4] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h000d3] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h001a6] : //%
                       Ifd35529b44c957737bf422127283c08e['h001a7] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000d4] =  Ifd35529b44c957737bf422127283c08e['h001a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000d5] =  Ifd35529b44c957737bf422127283c08e['h001aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000d6] =  Ifd35529b44c957737bf422127283c08e['h001ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000d7] =  Ifd35529b44c957737bf422127283c08e['h001ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000d8] =  Ifd35529b44c957737bf422127283c08e['h001b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000d9] =  Ifd35529b44c957737bf422127283c08e['h001b2] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h000da] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h001b4] : //%
                       Ifd35529b44c957737bf422127283c08e['h001b5] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000db] =  Ifd35529b44c957737bf422127283c08e['h001b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000dc] =  Ifd35529b44c957737bf422127283c08e['h001b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000dd] =  Ifd35529b44c957737bf422127283c08e['h001ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000de] =  Ifd35529b44c957737bf422127283c08e['h001bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000df] =  Ifd35529b44c957737bf422127283c08e['h001be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000e0] =  Ifd35529b44c957737bf422127283c08e['h001c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000e1] =  Ifd35529b44c957737bf422127283c08e['h001c2] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h000e2] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h001c4] : //%
                       Ifd35529b44c957737bf422127283c08e['h001c5] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000e3] =  Ifd35529b44c957737bf422127283c08e['h001c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000e4] =  Ifd35529b44c957737bf422127283c08e['h001c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000e5] =  Ifd35529b44c957737bf422127283c08e['h001ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000e6] =  Ifd35529b44c957737bf422127283c08e['h001cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000e7] =  Ifd35529b44c957737bf422127283c08e['h001ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000e8] =  Ifd35529b44c957737bf422127283c08e['h001d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000e9] =  Ifd35529b44c957737bf422127283c08e['h001d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000ea] =  Ifd35529b44c957737bf422127283c08e['h001d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000eb] =  Ifd35529b44c957737bf422127283c08e['h001d6] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h000ec] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h001d8] : //%
                       Ifd35529b44c957737bf422127283c08e['h001d9] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000ed] =  Ifd35529b44c957737bf422127283c08e['h001da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000ee] =  Ifd35529b44c957737bf422127283c08e['h001dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000ef] =  Ifd35529b44c957737bf422127283c08e['h001de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000f0] =  Ifd35529b44c957737bf422127283c08e['h001e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000f1] =  Ifd35529b44c957737bf422127283c08e['h001e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000f2] =  Ifd35529b44c957737bf422127283c08e['h001e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000f3] =  Ifd35529b44c957737bf422127283c08e['h001e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000f4] =  Ifd35529b44c957737bf422127283c08e['h001e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000f5] =  Ifd35529b44c957737bf422127283c08e['h001ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000f6] =  Ifd35529b44c957737bf422127283c08e['h001ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000f7] =  Ifd35529b44c957737bf422127283c08e['h001ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000f8] =  Ifd35529b44c957737bf422127283c08e['h001f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000f9] =  Ifd35529b44c957737bf422127283c08e['h001f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000fa] =  Ifd35529b44c957737bf422127283c08e['h001f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000fb] =  Ifd35529b44c957737bf422127283c08e['h001f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000fc] =  Ifd35529b44c957737bf422127283c08e['h001f8] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h000fd] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h001fa] : //%
                       Ifd35529b44c957737bf422127283c08e['h001fb] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000fe] =  Ifd35529b44c957737bf422127283c08e['h001fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h000ff] =  Ifd35529b44c957737bf422127283c08e['h001fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00100] =  Ifd35529b44c957737bf422127283c08e['h00200] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00101] =  Ifd35529b44c957737bf422127283c08e['h00202] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00102] =  Ifd35529b44c957737bf422127283c08e['h00204] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00103] =  Ifd35529b44c957737bf422127283c08e['h00206] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00104] =  Ifd35529b44c957737bf422127283c08e['h00208] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00105] =  Ifd35529b44c957737bf422127283c08e['h0020a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00106] =  Ifd35529b44c957737bf422127283c08e['h0020c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00107] =  Ifd35529b44c957737bf422127283c08e['h0020e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00108] =  Ifd35529b44c957737bf422127283c08e['h00210] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00109] =  Ifd35529b44c957737bf422127283c08e['h00212] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0010a] =  Ifd35529b44c957737bf422127283c08e['h00214] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0010b] =  Ifd35529b44c957737bf422127283c08e['h00216] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0010c] =  Ifd35529b44c957737bf422127283c08e['h00218] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0010d] =  Ifd35529b44c957737bf422127283c08e['h0021a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0010e] =  Ifd35529b44c957737bf422127283c08e['h0021c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0010f] =  Ifd35529b44c957737bf422127283c08e['h0021e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00110] =  Ifd35529b44c957737bf422127283c08e['h00220] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00111] =  Ifd35529b44c957737bf422127283c08e['h00222] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00112] =  Ifd35529b44c957737bf422127283c08e['h00224] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00113] =  Ifd35529b44c957737bf422127283c08e['h00226] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00114] =  Ifd35529b44c957737bf422127283c08e['h00228] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00115] =  Ifd35529b44c957737bf422127283c08e['h0022a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00116] =  Ifd35529b44c957737bf422127283c08e['h0022c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00117] =  Ifd35529b44c957737bf422127283c08e['h0022e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00118] =  Ifd35529b44c957737bf422127283c08e['h00230] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00119] =  Ifd35529b44c957737bf422127283c08e['h00232] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0011a] =  Ifd35529b44c957737bf422127283c08e['h00234] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0011b] =  Ifd35529b44c957737bf422127283c08e['h00236] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0011c] =  Ifd35529b44c957737bf422127283c08e['h00238] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0011d] =  Ifd35529b44c957737bf422127283c08e['h0023a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0011e] =  Ifd35529b44c957737bf422127283c08e['h0023c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0011f] =  Ifd35529b44c957737bf422127283c08e['h0023e] ;
//end
//always_comb begin
              If409768b648a33a7ed878a070d4f6251['h00120] = 
          (!fgallag_sel['h00005]) ? 
                       Ifd35529b44c957737bf422127283c08e['h00240] : //%
                       Ifd35529b44c957737bf422127283c08e['h00241] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00121] =  Ifd35529b44c957737bf422127283c08e['h00242] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00122] =  Ifd35529b44c957737bf422127283c08e['h00244] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00123] =  Ifd35529b44c957737bf422127283c08e['h00246] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00124] =  Ifd35529b44c957737bf422127283c08e['h00248] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00125] =  Ifd35529b44c957737bf422127283c08e['h0024a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00126] =  Ifd35529b44c957737bf422127283c08e['h0024c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00127] =  Ifd35529b44c957737bf422127283c08e['h0024e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00128] =  Ifd35529b44c957737bf422127283c08e['h00250] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00129] =  Ifd35529b44c957737bf422127283c08e['h00252] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0012a] =  Ifd35529b44c957737bf422127283c08e['h00254] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0012b] =  Ifd35529b44c957737bf422127283c08e['h00256] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0012c] =  Ifd35529b44c957737bf422127283c08e['h00258] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0012d] =  Ifd35529b44c957737bf422127283c08e['h0025a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0012e] =  Ifd35529b44c957737bf422127283c08e['h0025c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0012f] =  Ifd35529b44c957737bf422127283c08e['h0025e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00130] =  Ifd35529b44c957737bf422127283c08e['h00260] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00131] =  Ifd35529b44c957737bf422127283c08e['h00262] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00132] =  Ifd35529b44c957737bf422127283c08e['h00264] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00133] =  Ifd35529b44c957737bf422127283c08e['h00266] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00134] =  Ifd35529b44c957737bf422127283c08e['h00268] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00135] =  Ifd35529b44c957737bf422127283c08e['h0026a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00136] =  Ifd35529b44c957737bf422127283c08e['h0026c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00137] =  Ifd35529b44c957737bf422127283c08e['h0026e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00138] =  Ifd35529b44c957737bf422127283c08e['h00270] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00139] =  Ifd35529b44c957737bf422127283c08e['h00272] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0013a] =  Ifd35529b44c957737bf422127283c08e['h00274] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0013b] =  Ifd35529b44c957737bf422127283c08e['h00276] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0013c] =  Ifd35529b44c957737bf422127283c08e['h00278] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0013d] =  Ifd35529b44c957737bf422127283c08e['h0027a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0013e] =  Ifd35529b44c957737bf422127283c08e['h0027c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0013f] =  Ifd35529b44c957737bf422127283c08e['h0027e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00140] =  Ifd35529b44c957737bf422127283c08e['h00280] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00141] =  Ifd35529b44c957737bf422127283c08e['h00282] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00142] =  Ifd35529b44c957737bf422127283c08e['h00284] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00143] =  Ifd35529b44c957737bf422127283c08e['h00286] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00144] =  Ifd35529b44c957737bf422127283c08e['h00288] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00145] =  Ifd35529b44c957737bf422127283c08e['h0028a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00146] =  Ifd35529b44c957737bf422127283c08e['h0028c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00147] =  Ifd35529b44c957737bf422127283c08e['h0028e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00148] =  Ifd35529b44c957737bf422127283c08e['h00290] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00149] =  Ifd35529b44c957737bf422127283c08e['h00292] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0014a] =  Ifd35529b44c957737bf422127283c08e['h00294] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0014b] =  Ifd35529b44c957737bf422127283c08e['h00296] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0014c] =  Ifd35529b44c957737bf422127283c08e['h00298] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0014d] =  Ifd35529b44c957737bf422127283c08e['h0029a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0014e] =  Ifd35529b44c957737bf422127283c08e['h0029c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0014f] =  Ifd35529b44c957737bf422127283c08e['h0029e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00150] =  Ifd35529b44c957737bf422127283c08e['h002a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00151] =  Ifd35529b44c957737bf422127283c08e['h002a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00152] =  Ifd35529b44c957737bf422127283c08e['h002a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00153] =  Ifd35529b44c957737bf422127283c08e['h002a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00154] =  Ifd35529b44c957737bf422127283c08e['h002a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00155] =  Ifd35529b44c957737bf422127283c08e['h002aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00156] =  Ifd35529b44c957737bf422127283c08e['h002ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00157] =  Ifd35529b44c957737bf422127283c08e['h002ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00158] =  Ifd35529b44c957737bf422127283c08e['h002b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00159] =  Ifd35529b44c957737bf422127283c08e['h002b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0015a] =  Ifd35529b44c957737bf422127283c08e['h002b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0015b] =  Ifd35529b44c957737bf422127283c08e['h002b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0015c] =  Ifd35529b44c957737bf422127283c08e['h002b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0015d] =  Ifd35529b44c957737bf422127283c08e['h002ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0015e] =  Ifd35529b44c957737bf422127283c08e['h002bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0015f] =  Ifd35529b44c957737bf422127283c08e['h002be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00160] =  Ifd35529b44c957737bf422127283c08e['h002c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00161] =  Ifd35529b44c957737bf422127283c08e['h002c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00162] =  Ifd35529b44c957737bf422127283c08e['h002c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00163] =  Ifd35529b44c957737bf422127283c08e['h002c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00164] =  Ifd35529b44c957737bf422127283c08e['h002c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00165] =  Ifd35529b44c957737bf422127283c08e['h002ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00166] =  Ifd35529b44c957737bf422127283c08e['h002cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00167] =  Ifd35529b44c957737bf422127283c08e['h002ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00168] =  Ifd35529b44c957737bf422127283c08e['h002d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00169] =  Ifd35529b44c957737bf422127283c08e['h002d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0016a] =  Ifd35529b44c957737bf422127283c08e['h002d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0016b] =  Ifd35529b44c957737bf422127283c08e['h002d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0016c] =  Ifd35529b44c957737bf422127283c08e['h002d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0016d] =  Ifd35529b44c957737bf422127283c08e['h002da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0016e] =  Ifd35529b44c957737bf422127283c08e['h002dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0016f] =  Ifd35529b44c957737bf422127283c08e['h002de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00170] =  Ifd35529b44c957737bf422127283c08e['h002e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00171] =  Ifd35529b44c957737bf422127283c08e['h002e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00172] =  Ifd35529b44c957737bf422127283c08e['h002e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00173] =  Ifd35529b44c957737bf422127283c08e['h002e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00174] =  Ifd35529b44c957737bf422127283c08e['h002e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00175] =  Ifd35529b44c957737bf422127283c08e['h002ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00176] =  Ifd35529b44c957737bf422127283c08e['h002ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00177] =  Ifd35529b44c957737bf422127283c08e['h002ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00178] =  Ifd35529b44c957737bf422127283c08e['h002f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00179] =  Ifd35529b44c957737bf422127283c08e['h002f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0017a] =  Ifd35529b44c957737bf422127283c08e['h002f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0017b] =  Ifd35529b44c957737bf422127283c08e['h002f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0017c] =  Ifd35529b44c957737bf422127283c08e['h002f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0017d] =  Ifd35529b44c957737bf422127283c08e['h002fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0017e] =  Ifd35529b44c957737bf422127283c08e['h002fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0017f] =  Ifd35529b44c957737bf422127283c08e['h002fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00180] =  Ifd35529b44c957737bf422127283c08e['h00300] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00181] =  Ifd35529b44c957737bf422127283c08e['h00302] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00182] =  Ifd35529b44c957737bf422127283c08e['h00304] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00183] =  Ifd35529b44c957737bf422127283c08e['h00306] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00184] =  Ifd35529b44c957737bf422127283c08e['h00308] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00185] =  Ifd35529b44c957737bf422127283c08e['h0030a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00186] =  Ifd35529b44c957737bf422127283c08e['h0030c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00187] =  Ifd35529b44c957737bf422127283c08e['h0030e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00188] =  Ifd35529b44c957737bf422127283c08e['h00310] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00189] =  Ifd35529b44c957737bf422127283c08e['h00312] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0018a] =  Ifd35529b44c957737bf422127283c08e['h00314] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0018b] =  Ifd35529b44c957737bf422127283c08e['h00316] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0018c] =  Ifd35529b44c957737bf422127283c08e['h00318] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0018d] =  Ifd35529b44c957737bf422127283c08e['h0031a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0018e] =  Ifd35529b44c957737bf422127283c08e['h0031c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0018f] =  Ifd35529b44c957737bf422127283c08e['h0031e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00190] =  Ifd35529b44c957737bf422127283c08e['h00320] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00191] =  Ifd35529b44c957737bf422127283c08e['h00322] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00192] =  Ifd35529b44c957737bf422127283c08e['h00324] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00193] =  Ifd35529b44c957737bf422127283c08e['h00326] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00194] =  Ifd35529b44c957737bf422127283c08e['h00328] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00195] =  Ifd35529b44c957737bf422127283c08e['h0032a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00196] =  Ifd35529b44c957737bf422127283c08e['h0032c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00197] =  Ifd35529b44c957737bf422127283c08e['h0032e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00198] =  Ifd35529b44c957737bf422127283c08e['h00330] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00199] =  Ifd35529b44c957737bf422127283c08e['h00332] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0019a] =  Ifd35529b44c957737bf422127283c08e['h00334] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0019b] =  Ifd35529b44c957737bf422127283c08e['h00336] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0019c] =  Ifd35529b44c957737bf422127283c08e['h00338] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0019d] =  Ifd35529b44c957737bf422127283c08e['h0033a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0019e] =  Ifd35529b44c957737bf422127283c08e['h0033c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0019f] =  Ifd35529b44c957737bf422127283c08e['h0033e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001a0] =  Ifd35529b44c957737bf422127283c08e['h00340] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001a1] =  Ifd35529b44c957737bf422127283c08e['h00342] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001a2] =  Ifd35529b44c957737bf422127283c08e['h00344] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001a3] =  Ifd35529b44c957737bf422127283c08e['h00346] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001a4] =  Ifd35529b44c957737bf422127283c08e['h00348] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001a5] =  Ifd35529b44c957737bf422127283c08e['h0034a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001a6] =  Ifd35529b44c957737bf422127283c08e['h0034c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001a7] =  Ifd35529b44c957737bf422127283c08e['h0034e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001a8] =  Ifd35529b44c957737bf422127283c08e['h00350] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001a9] =  Ifd35529b44c957737bf422127283c08e['h00352] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001aa] =  Ifd35529b44c957737bf422127283c08e['h00354] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001ab] =  Ifd35529b44c957737bf422127283c08e['h00356] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001ac] =  Ifd35529b44c957737bf422127283c08e['h00358] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001ad] =  Ifd35529b44c957737bf422127283c08e['h0035a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001ae] =  Ifd35529b44c957737bf422127283c08e['h0035c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001af] =  Ifd35529b44c957737bf422127283c08e['h0035e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001b0] =  Ifd35529b44c957737bf422127283c08e['h00360] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001b1] =  Ifd35529b44c957737bf422127283c08e['h00362] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001b2] =  Ifd35529b44c957737bf422127283c08e['h00364] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001b3] =  Ifd35529b44c957737bf422127283c08e['h00366] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001b4] =  Ifd35529b44c957737bf422127283c08e['h00368] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001b5] =  Ifd35529b44c957737bf422127283c08e['h0036a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001b6] =  Ifd35529b44c957737bf422127283c08e['h0036c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001b7] =  Ifd35529b44c957737bf422127283c08e['h0036e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001b8] =  Ifd35529b44c957737bf422127283c08e['h00370] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001b9] =  Ifd35529b44c957737bf422127283c08e['h00372] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001ba] =  Ifd35529b44c957737bf422127283c08e['h00374] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001bb] =  Ifd35529b44c957737bf422127283c08e['h00376] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001bc] =  Ifd35529b44c957737bf422127283c08e['h00378] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001bd] =  Ifd35529b44c957737bf422127283c08e['h0037a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001be] =  Ifd35529b44c957737bf422127283c08e['h0037c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001bf] =  Ifd35529b44c957737bf422127283c08e['h0037e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001c0] =  Ifd35529b44c957737bf422127283c08e['h00380] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001c1] =  Ifd35529b44c957737bf422127283c08e['h00382] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001c2] =  Ifd35529b44c957737bf422127283c08e['h00384] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001c3] =  Ifd35529b44c957737bf422127283c08e['h00386] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001c4] =  Ifd35529b44c957737bf422127283c08e['h00388] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001c5] =  Ifd35529b44c957737bf422127283c08e['h0038a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001c6] =  Ifd35529b44c957737bf422127283c08e['h0038c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001c7] =  Ifd35529b44c957737bf422127283c08e['h0038e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001c8] =  Ifd35529b44c957737bf422127283c08e['h00390] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001c9] =  Ifd35529b44c957737bf422127283c08e['h00392] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001ca] =  Ifd35529b44c957737bf422127283c08e['h00394] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001cb] =  Ifd35529b44c957737bf422127283c08e['h00396] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001cc] =  Ifd35529b44c957737bf422127283c08e['h00398] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001cd] =  Ifd35529b44c957737bf422127283c08e['h0039a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001ce] =  Ifd35529b44c957737bf422127283c08e['h0039c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001cf] =  Ifd35529b44c957737bf422127283c08e['h0039e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001d0] =  Ifd35529b44c957737bf422127283c08e['h003a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001d1] =  Ifd35529b44c957737bf422127283c08e['h003a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001d2] =  Ifd35529b44c957737bf422127283c08e['h003a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001d3] =  Ifd35529b44c957737bf422127283c08e['h003a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001d4] =  Ifd35529b44c957737bf422127283c08e['h003a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001d5] =  Ifd35529b44c957737bf422127283c08e['h003aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001d6] =  Ifd35529b44c957737bf422127283c08e['h003ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001d7] =  Ifd35529b44c957737bf422127283c08e['h003ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001d8] =  Ifd35529b44c957737bf422127283c08e['h003b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001d9] =  Ifd35529b44c957737bf422127283c08e['h003b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001da] =  Ifd35529b44c957737bf422127283c08e['h003b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001db] =  Ifd35529b44c957737bf422127283c08e['h003b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001dc] =  Ifd35529b44c957737bf422127283c08e['h003b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001dd] =  Ifd35529b44c957737bf422127283c08e['h003ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001de] =  Ifd35529b44c957737bf422127283c08e['h003bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001df] =  Ifd35529b44c957737bf422127283c08e['h003be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001e0] =  Ifd35529b44c957737bf422127283c08e['h003c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001e1] =  Ifd35529b44c957737bf422127283c08e['h003c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001e2] =  Ifd35529b44c957737bf422127283c08e['h003c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001e3] =  Ifd35529b44c957737bf422127283c08e['h003c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001e4] =  Ifd35529b44c957737bf422127283c08e['h003c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001e5] =  Ifd35529b44c957737bf422127283c08e['h003ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001e6] =  Ifd35529b44c957737bf422127283c08e['h003cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001e7] =  Ifd35529b44c957737bf422127283c08e['h003ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001e8] =  Ifd35529b44c957737bf422127283c08e['h003d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001e9] =  Ifd35529b44c957737bf422127283c08e['h003d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001ea] =  Ifd35529b44c957737bf422127283c08e['h003d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001eb] =  Ifd35529b44c957737bf422127283c08e['h003d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001ec] =  Ifd35529b44c957737bf422127283c08e['h003d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001ed] =  Ifd35529b44c957737bf422127283c08e['h003da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001ee] =  Ifd35529b44c957737bf422127283c08e['h003dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001ef] =  Ifd35529b44c957737bf422127283c08e['h003de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001f0] =  Ifd35529b44c957737bf422127283c08e['h003e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001f1] =  Ifd35529b44c957737bf422127283c08e['h003e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001f2] =  Ifd35529b44c957737bf422127283c08e['h003e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001f3] =  Ifd35529b44c957737bf422127283c08e['h003e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001f4] =  Ifd35529b44c957737bf422127283c08e['h003e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001f5] =  Ifd35529b44c957737bf422127283c08e['h003ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001f6] =  Ifd35529b44c957737bf422127283c08e['h003ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001f7] =  Ifd35529b44c957737bf422127283c08e['h003ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001f8] =  Ifd35529b44c957737bf422127283c08e['h003f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001f9] =  Ifd35529b44c957737bf422127283c08e['h003f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001fa] =  Ifd35529b44c957737bf422127283c08e['h003f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001fb] =  Ifd35529b44c957737bf422127283c08e['h003f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001fc] =  Ifd35529b44c957737bf422127283c08e['h003f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001fd] =  Ifd35529b44c957737bf422127283c08e['h003fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001fe] =  Ifd35529b44c957737bf422127283c08e['h003fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h001ff] =  Ifd35529b44c957737bf422127283c08e['h003fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00200] =  Ifd35529b44c957737bf422127283c08e['h00400] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00201] =  Ifd35529b44c957737bf422127283c08e['h00402] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00202] =  Ifd35529b44c957737bf422127283c08e['h00404] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00203] =  Ifd35529b44c957737bf422127283c08e['h00406] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00204] =  Ifd35529b44c957737bf422127283c08e['h00408] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00205] =  Ifd35529b44c957737bf422127283c08e['h0040a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00206] =  Ifd35529b44c957737bf422127283c08e['h0040c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00207] =  Ifd35529b44c957737bf422127283c08e['h0040e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00208] =  Ifd35529b44c957737bf422127283c08e['h00410] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00209] =  Ifd35529b44c957737bf422127283c08e['h00412] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0020a] =  Ifd35529b44c957737bf422127283c08e['h00414] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0020b] =  Ifd35529b44c957737bf422127283c08e['h00416] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0020c] =  Ifd35529b44c957737bf422127283c08e['h00418] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0020d] =  Ifd35529b44c957737bf422127283c08e['h0041a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0020e] =  Ifd35529b44c957737bf422127283c08e['h0041c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0020f] =  Ifd35529b44c957737bf422127283c08e['h0041e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00210] =  Ifd35529b44c957737bf422127283c08e['h00420] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00211] =  Ifd35529b44c957737bf422127283c08e['h00422] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00212] =  Ifd35529b44c957737bf422127283c08e['h00424] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00213] =  Ifd35529b44c957737bf422127283c08e['h00426] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00214] =  Ifd35529b44c957737bf422127283c08e['h00428] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00215] =  Ifd35529b44c957737bf422127283c08e['h0042a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00216] =  Ifd35529b44c957737bf422127283c08e['h0042c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00217] =  Ifd35529b44c957737bf422127283c08e['h0042e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00218] =  Ifd35529b44c957737bf422127283c08e['h00430] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00219] =  Ifd35529b44c957737bf422127283c08e['h00432] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0021a] =  Ifd35529b44c957737bf422127283c08e['h00434] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0021b] =  Ifd35529b44c957737bf422127283c08e['h00436] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0021c] =  Ifd35529b44c957737bf422127283c08e['h00438] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0021d] =  Ifd35529b44c957737bf422127283c08e['h0043a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0021e] =  Ifd35529b44c957737bf422127283c08e['h0043c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0021f] =  Ifd35529b44c957737bf422127283c08e['h0043e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00220] =  Ifd35529b44c957737bf422127283c08e['h00440] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00221] =  Ifd35529b44c957737bf422127283c08e['h00442] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00222] =  Ifd35529b44c957737bf422127283c08e['h00444] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00223] =  Ifd35529b44c957737bf422127283c08e['h00446] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00224] =  Ifd35529b44c957737bf422127283c08e['h00448] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00225] =  Ifd35529b44c957737bf422127283c08e['h0044a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00226] =  Ifd35529b44c957737bf422127283c08e['h0044c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00227] =  Ifd35529b44c957737bf422127283c08e['h0044e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00228] =  Ifd35529b44c957737bf422127283c08e['h00450] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00229] =  Ifd35529b44c957737bf422127283c08e['h00452] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0022a] =  Ifd35529b44c957737bf422127283c08e['h00454] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0022b] =  Ifd35529b44c957737bf422127283c08e['h00456] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0022c] =  Ifd35529b44c957737bf422127283c08e['h00458] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0022d] =  Ifd35529b44c957737bf422127283c08e['h0045a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0022e] =  Ifd35529b44c957737bf422127283c08e['h0045c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0022f] =  Ifd35529b44c957737bf422127283c08e['h0045e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00230] =  Ifd35529b44c957737bf422127283c08e['h00460] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00231] =  Ifd35529b44c957737bf422127283c08e['h00462] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00232] =  Ifd35529b44c957737bf422127283c08e['h00464] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00233] =  Ifd35529b44c957737bf422127283c08e['h00466] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00234] =  Ifd35529b44c957737bf422127283c08e['h00468] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00235] =  Ifd35529b44c957737bf422127283c08e['h0046a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00236] =  Ifd35529b44c957737bf422127283c08e['h0046c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00237] =  Ifd35529b44c957737bf422127283c08e['h0046e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00238] =  Ifd35529b44c957737bf422127283c08e['h00470] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00239] =  Ifd35529b44c957737bf422127283c08e['h00472] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0023a] =  Ifd35529b44c957737bf422127283c08e['h00474] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0023b] =  Ifd35529b44c957737bf422127283c08e['h00476] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0023c] =  Ifd35529b44c957737bf422127283c08e['h00478] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0023d] =  Ifd35529b44c957737bf422127283c08e['h0047a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0023e] =  Ifd35529b44c957737bf422127283c08e['h0047c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0023f] =  Ifd35529b44c957737bf422127283c08e['h0047e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00240] =  Ifd35529b44c957737bf422127283c08e['h00480] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00241] =  Ifd35529b44c957737bf422127283c08e['h00482] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00242] =  Ifd35529b44c957737bf422127283c08e['h00484] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00243] =  Ifd35529b44c957737bf422127283c08e['h00486] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00244] =  Ifd35529b44c957737bf422127283c08e['h00488] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00245] =  Ifd35529b44c957737bf422127283c08e['h0048a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00246] =  Ifd35529b44c957737bf422127283c08e['h0048c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00247] =  Ifd35529b44c957737bf422127283c08e['h0048e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00248] =  Ifd35529b44c957737bf422127283c08e['h00490] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00249] =  Ifd35529b44c957737bf422127283c08e['h00492] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0024a] =  Ifd35529b44c957737bf422127283c08e['h00494] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0024b] =  Ifd35529b44c957737bf422127283c08e['h00496] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0024c] =  Ifd35529b44c957737bf422127283c08e['h00498] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0024d] =  Ifd35529b44c957737bf422127283c08e['h0049a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0024e] =  Ifd35529b44c957737bf422127283c08e['h0049c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0024f] =  Ifd35529b44c957737bf422127283c08e['h0049e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00250] =  Ifd35529b44c957737bf422127283c08e['h004a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00251] =  Ifd35529b44c957737bf422127283c08e['h004a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00252] =  Ifd35529b44c957737bf422127283c08e['h004a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00253] =  Ifd35529b44c957737bf422127283c08e['h004a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00254] =  Ifd35529b44c957737bf422127283c08e['h004a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00255] =  Ifd35529b44c957737bf422127283c08e['h004aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00256] =  Ifd35529b44c957737bf422127283c08e['h004ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00257] =  Ifd35529b44c957737bf422127283c08e['h004ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00258] =  Ifd35529b44c957737bf422127283c08e['h004b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00259] =  Ifd35529b44c957737bf422127283c08e['h004b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0025a] =  Ifd35529b44c957737bf422127283c08e['h004b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0025b] =  Ifd35529b44c957737bf422127283c08e['h004b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0025c] =  Ifd35529b44c957737bf422127283c08e['h004b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0025d] =  Ifd35529b44c957737bf422127283c08e['h004ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0025e] =  Ifd35529b44c957737bf422127283c08e['h004bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0025f] =  Ifd35529b44c957737bf422127283c08e['h004be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00260] =  Ifd35529b44c957737bf422127283c08e['h004c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00261] =  Ifd35529b44c957737bf422127283c08e['h004c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00262] =  Ifd35529b44c957737bf422127283c08e['h004c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00263] =  Ifd35529b44c957737bf422127283c08e['h004c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00264] =  Ifd35529b44c957737bf422127283c08e['h004c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00265] =  Ifd35529b44c957737bf422127283c08e['h004ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00266] =  Ifd35529b44c957737bf422127283c08e['h004cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00267] =  Ifd35529b44c957737bf422127283c08e['h004ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00268] =  Ifd35529b44c957737bf422127283c08e['h004d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00269] =  Ifd35529b44c957737bf422127283c08e['h004d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0026a] =  Ifd35529b44c957737bf422127283c08e['h004d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0026b] =  Ifd35529b44c957737bf422127283c08e['h004d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0026c] =  Ifd35529b44c957737bf422127283c08e['h004d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0026d] =  Ifd35529b44c957737bf422127283c08e['h004da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0026e] =  Ifd35529b44c957737bf422127283c08e['h004dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0026f] =  Ifd35529b44c957737bf422127283c08e['h004de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00270] =  Ifd35529b44c957737bf422127283c08e['h004e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00271] =  Ifd35529b44c957737bf422127283c08e['h004e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00272] =  Ifd35529b44c957737bf422127283c08e['h004e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00273] =  Ifd35529b44c957737bf422127283c08e['h004e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00274] =  Ifd35529b44c957737bf422127283c08e['h004e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00275] =  Ifd35529b44c957737bf422127283c08e['h004ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00276] =  Ifd35529b44c957737bf422127283c08e['h004ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00277] =  Ifd35529b44c957737bf422127283c08e['h004ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00278] =  Ifd35529b44c957737bf422127283c08e['h004f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00279] =  Ifd35529b44c957737bf422127283c08e['h004f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0027a] =  Ifd35529b44c957737bf422127283c08e['h004f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0027b] =  Ifd35529b44c957737bf422127283c08e['h004f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0027c] =  Ifd35529b44c957737bf422127283c08e['h004f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0027d] =  Ifd35529b44c957737bf422127283c08e['h004fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0027e] =  Ifd35529b44c957737bf422127283c08e['h004fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0027f] =  Ifd35529b44c957737bf422127283c08e['h004fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00280] =  Ifd35529b44c957737bf422127283c08e['h00500] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00281] =  Ifd35529b44c957737bf422127283c08e['h00502] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00282] =  Ifd35529b44c957737bf422127283c08e['h00504] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00283] =  Ifd35529b44c957737bf422127283c08e['h00506] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00284] =  Ifd35529b44c957737bf422127283c08e['h00508] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00285] =  Ifd35529b44c957737bf422127283c08e['h0050a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00286] =  Ifd35529b44c957737bf422127283c08e['h0050c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00287] =  Ifd35529b44c957737bf422127283c08e['h0050e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00288] =  Ifd35529b44c957737bf422127283c08e['h00510] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00289] =  Ifd35529b44c957737bf422127283c08e['h00512] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0028a] =  Ifd35529b44c957737bf422127283c08e['h00514] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0028b] =  Ifd35529b44c957737bf422127283c08e['h00516] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0028c] =  Ifd35529b44c957737bf422127283c08e['h00518] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0028d] =  Ifd35529b44c957737bf422127283c08e['h0051a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0028e] =  Ifd35529b44c957737bf422127283c08e['h0051c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0028f] =  Ifd35529b44c957737bf422127283c08e['h0051e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00290] =  Ifd35529b44c957737bf422127283c08e['h00520] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00291] =  Ifd35529b44c957737bf422127283c08e['h00522] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00292] =  Ifd35529b44c957737bf422127283c08e['h00524] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00293] =  Ifd35529b44c957737bf422127283c08e['h00526] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00294] =  Ifd35529b44c957737bf422127283c08e['h00528] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00295] =  Ifd35529b44c957737bf422127283c08e['h0052a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00296] =  Ifd35529b44c957737bf422127283c08e['h0052c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00297] =  Ifd35529b44c957737bf422127283c08e['h0052e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00298] =  Ifd35529b44c957737bf422127283c08e['h00530] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00299] =  Ifd35529b44c957737bf422127283c08e['h00532] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0029a] =  Ifd35529b44c957737bf422127283c08e['h00534] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0029b] =  Ifd35529b44c957737bf422127283c08e['h00536] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0029c] =  Ifd35529b44c957737bf422127283c08e['h00538] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0029d] =  Ifd35529b44c957737bf422127283c08e['h0053a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0029e] =  Ifd35529b44c957737bf422127283c08e['h0053c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0029f] =  Ifd35529b44c957737bf422127283c08e['h0053e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002a0] =  Ifd35529b44c957737bf422127283c08e['h00540] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002a1] =  Ifd35529b44c957737bf422127283c08e['h00542] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002a2] =  Ifd35529b44c957737bf422127283c08e['h00544] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002a3] =  Ifd35529b44c957737bf422127283c08e['h00546] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002a4] =  Ifd35529b44c957737bf422127283c08e['h00548] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002a5] =  Ifd35529b44c957737bf422127283c08e['h0054a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002a6] =  Ifd35529b44c957737bf422127283c08e['h0054c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002a7] =  Ifd35529b44c957737bf422127283c08e['h0054e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002a8] =  Ifd35529b44c957737bf422127283c08e['h00550] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002a9] =  Ifd35529b44c957737bf422127283c08e['h00552] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002aa] =  Ifd35529b44c957737bf422127283c08e['h00554] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002ab] =  Ifd35529b44c957737bf422127283c08e['h00556] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002ac] =  Ifd35529b44c957737bf422127283c08e['h00558] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002ad] =  Ifd35529b44c957737bf422127283c08e['h0055a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002ae] =  Ifd35529b44c957737bf422127283c08e['h0055c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002af] =  Ifd35529b44c957737bf422127283c08e['h0055e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002b0] =  Ifd35529b44c957737bf422127283c08e['h00560] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002b1] =  Ifd35529b44c957737bf422127283c08e['h00562] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002b2] =  Ifd35529b44c957737bf422127283c08e['h00564] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002b3] =  Ifd35529b44c957737bf422127283c08e['h00566] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002b4] =  Ifd35529b44c957737bf422127283c08e['h00568] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002b5] =  Ifd35529b44c957737bf422127283c08e['h0056a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002b6] =  Ifd35529b44c957737bf422127283c08e['h0056c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002b7] =  Ifd35529b44c957737bf422127283c08e['h0056e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002b8] =  Ifd35529b44c957737bf422127283c08e['h00570] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002b9] =  Ifd35529b44c957737bf422127283c08e['h00572] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002ba] =  Ifd35529b44c957737bf422127283c08e['h00574] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002bb] =  Ifd35529b44c957737bf422127283c08e['h00576] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002bc] =  Ifd35529b44c957737bf422127283c08e['h00578] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002bd] =  Ifd35529b44c957737bf422127283c08e['h0057a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002be] =  Ifd35529b44c957737bf422127283c08e['h0057c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002bf] =  Ifd35529b44c957737bf422127283c08e['h0057e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002c0] =  Ifd35529b44c957737bf422127283c08e['h00580] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002c1] =  Ifd35529b44c957737bf422127283c08e['h00582] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002c2] =  Ifd35529b44c957737bf422127283c08e['h00584] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002c3] =  Ifd35529b44c957737bf422127283c08e['h00586] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002c4] =  Ifd35529b44c957737bf422127283c08e['h00588] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002c5] =  Ifd35529b44c957737bf422127283c08e['h0058a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002c6] =  Ifd35529b44c957737bf422127283c08e['h0058c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002c7] =  Ifd35529b44c957737bf422127283c08e['h0058e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002c8] =  Ifd35529b44c957737bf422127283c08e['h00590] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002c9] =  Ifd35529b44c957737bf422127283c08e['h00592] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002ca] =  Ifd35529b44c957737bf422127283c08e['h00594] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002cb] =  Ifd35529b44c957737bf422127283c08e['h00596] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002cc] =  Ifd35529b44c957737bf422127283c08e['h00598] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002cd] =  Ifd35529b44c957737bf422127283c08e['h0059a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002ce] =  Ifd35529b44c957737bf422127283c08e['h0059c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002cf] =  Ifd35529b44c957737bf422127283c08e['h0059e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002d0] =  Ifd35529b44c957737bf422127283c08e['h005a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002d1] =  Ifd35529b44c957737bf422127283c08e['h005a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002d2] =  Ifd35529b44c957737bf422127283c08e['h005a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002d3] =  Ifd35529b44c957737bf422127283c08e['h005a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002d4] =  Ifd35529b44c957737bf422127283c08e['h005a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002d5] =  Ifd35529b44c957737bf422127283c08e['h005aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002d6] =  Ifd35529b44c957737bf422127283c08e['h005ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002d7] =  Ifd35529b44c957737bf422127283c08e['h005ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002d8] =  Ifd35529b44c957737bf422127283c08e['h005b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002d9] =  Ifd35529b44c957737bf422127283c08e['h005b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002da] =  Ifd35529b44c957737bf422127283c08e['h005b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002db] =  Ifd35529b44c957737bf422127283c08e['h005b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002dc] =  Ifd35529b44c957737bf422127283c08e['h005b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002dd] =  Ifd35529b44c957737bf422127283c08e['h005ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002de] =  Ifd35529b44c957737bf422127283c08e['h005bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002df] =  Ifd35529b44c957737bf422127283c08e['h005be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002e0] =  Ifd35529b44c957737bf422127283c08e['h005c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002e1] =  Ifd35529b44c957737bf422127283c08e['h005c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002e2] =  Ifd35529b44c957737bf422127283c08e['h005c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002e3] =  Ifd35529b44c957737bf422127283c08e['h005c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002e4] =  Ifd35529b44c957737bf422127283c08e['h005c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002e5] =  Ifd35529b44c957737bf422127283c08e['h005ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002e6] =  Ifd35529b44c957737bf422127283c08e['h005cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002e7] =  Ifd35529b44c957737bf422127283c08e['h005ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002e8] =  Ifd35529b44c957737bf422127283c08e['h005d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002e9] =  Ifd35529b44c957737bf422127283c08e['h005d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002ea] =  Ifd35529b44c957737bf422127283c08e['h005d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002eb] =  Ifd35529b44c957737bf422127283c08e['h005d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002ec] =  Ifd35529b44c957737bf422127283c08e['h005d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002ed] =  Ifd35529b44c957737bf422127283c08e['h005da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002ee] =  Ifd35529b44c957737bf422127283c08e['h005dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002ef] =  Ifd35529b44c957737bf422127283c08e['h005de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002f0] =  Ifd35529b44c957737bf422127283c08e['h005e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002f1] =  Ifd35529b44c957737bf422127283c08e['h005e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002f2] =  Ifd35529b44c957737bf422127283c08e['h005e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002f3] =  Ifd35529b44c957737bf422127283c08e['h005e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002f4] =  Ifd35529b44c957737bf422127283c08e['h005e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002f5] =  Ifd35529b44c957737bf422127283c08e['h005ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002f6] =  Ifd35529b44c957737bf422127283c08e['h005ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002f7] =  Ifd35529b44c957737bf422127283c08e['h005ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002f8] =  Ifd35529b44c957737bf422127283c08e['h005f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002f9] =  Ifd35529b44c957737bf422127283c08e['h005f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002fa] =  Ifd35529b44c957737bf422127283c08e['h005f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002fb] =  Ifd35529b44c957737bf422127283c08e['h005f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002fc] =  Ifd35529b44c957737bf422127283c08e['h005f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002fd] =  Ifd35529b44c957737bf422127283c08e['h005fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002fe] =  Ifd35529b44c957737bf422127283c08e['h005fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h002ff] =  Ifd35529b44c957737bf422127283c08e['h005fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00300] =  Ifd35529b44c957737bf422127283c08e['h00600] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00301] =  Ifd35529b44c957737bf422127283c08e['h00602] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00302] =  Ifd35529b44c957737bf422127283c08e['h00604] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00303] =  Ifd35529b44c957737bf422127283c08e['h00606] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00304] =  Ifd35529b44c957737bf422127283c08e['h00608] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00305] =  Ifd35529b44c957737bf422127283c08e['h0060a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00306] =  Ifd35529b44c957737bf422127283c08e['h0060c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00307] =  Ifd35529b44c957737bf422127283c08e['h0060e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00308] =  Ifd35529b44c957737bf422127283c08e['h00610] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00309] =  Ifd35529b44c957737bf422127283c08e['h00612] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0030a] =  Ifd35529b44c957737bf422127283c08e['h00614] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0030b] =  Ifd35529b44c957737bf422127283c08e['h00616] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0030c] =  Ifd35529b44c957737bf422127283c08e['h00618] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0030d] =  Ifd35529b44c957737bf422127283c08e['h0061a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0030e] =  Ifd35529b44c957737bf422127283c08e['h0061c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0030f] =  Ifd35529b44c957737bf422127283c08e['h0061e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00310] =  Ifd35529b44c957737bf422127283c08e['h00620] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00311] =  Ifd35529b44c957737bf422127283c08e['h00622] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00312] =  Ifd35529b44c957737bf422127283c08e['h00624] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00313] =  Ifd35529b44c957737bf422127283c08e['h00626] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00314] =  Ifd35529b44c957737bf422127283c08e['h00628] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00315] =  Ifd35529b44c957737bf422127283c08e['h0062a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00316] =  Ifd35529b44c957737bf422127283c08e['h0062c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00317] =  Ifd35529b44c957737bf422127283c08e['h0062e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00318] =  Ifd35529b44c957737bf422127283c08e['h00630] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00319] =  Ifd35529b44c957737bf422127283c08e['h00632] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0031a] =  Ifd35529b44c957737bf422127283c08e['h00634] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0031b] =  Ifd35529b44c957737bf422127283c08e['h00636] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0031c] =  Ifd35529b44c957737bf422127283c08e['h00638] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0031d] =  Ifd35529b44c957737bf422127283c08e['h0063a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0031e] =  Ifd35529b44c957737bf422127283c08e['h0063c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0031f] =  Ifd35529b44c957737bf422127283c08e['h0063e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00320] =  Ifd35529b44c957737bf422127283c08e['h00640] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00321] =  Ifd35529b44c957737bf422127283c08e['h00642] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00322] =  Ifd35529b44c957737bf422127283c08e['h00644] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00323] =  Ifd35529b44c957737bf422127283c08e['h00646] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00324] =  Ifd35529b44c957737bf422127283c08e['h00648] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00325] =  Ifd35529b44c957737bf422127283c08e['h0064a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00326] =  Ifd35529b44c957737bf422127283c08e['h0064c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00327] =  Ifd35529b44c957737bf422127283c08e['h0064e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00328] =  Ifd35529b44c957737bf422127283c08e['h00650] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00329] =  Ifd35529b44c957737bf422127283c08e['h00652] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0032a] =  Ifd35529b44c957737bf422127283c08e['h00654] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0032b] =  Ifd35529b44c957737bf422127283c08e['h00656] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0032c] =  Ifd35529b44c957737bf422127283c08e['h00658] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0032d] =  Ifd35529b44c957737bf422127283c08e['h0065a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0032e] =  Ifd35529b44c957737bf422127283c08e['h0065c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0032f] =  Ifd35529b44c957737bf422127283c08e['h0065e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00330] =  Ifd35529b44c957737bf422127283c08e['h00660] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00331] =  Ifd35529b44c957737bf422127283c08e['h00662] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00332] =  Ifd35529b44c957737bf422127283c08e['h00664] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00333] =  Ifd35529b44c957737bf422127283c08e['h00666] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00334] =  Ifd35529b44c957737bf422127283c08e['h00668] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00335] =  Ifd35529b44c957737bf422127283c08e['h0066a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00336] =  Ifd35529b44c957737bf422127283c08e['h0066c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00337] =  Ifd35529b44c957737bf422127283c08e['h0066e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00338] =  Ifd35529b44c957737bf422127283c08e['h00670] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00339] =  Ifd35529b44c957737bf422127283c08e['h00672] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0033a] =  Ifd35529b44c957737bf422127283c08e['h00674] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0033b] =  Ifd35529b44c957737bf422127283c08e['h00676] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0033c] =  Ifd35529b44c957737bf422127283c08e['h00678] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0033d] =  Ifd35529b44c957737bf422127283c08e['h0067a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0033e] =  Ifd35529b44c957737bf422127283c08e['h0067c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0033f] =  Ifd35529b44c957737bf422127283c08e['h0067e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00340] =  Ifd35529b44c957737bf422127283c08e['h00680] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00341] =  Ifd35529b44c957737bf422127283c08e['h00682] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00342] =  Ifd35529b44c957737bf422127283c08e['h00684] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00343] =  Ifd35529b44c957737bf422127283c08e['h00686] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00344] =  Ifd35529b44c957737bf422127283c08e['h00688] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00345] =  Ifd35529b44c957737bf422127283c08e['h0068a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00346] =  Ifd35529b44c957737bf422127283c08e['h0068c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00347] =  Ifd35529b44c957737bf422127283c08e['h0068e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00348] =  Ifd35529b44c957737bf422127283c08e['h00690] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00349] =  Ifd35529b44c957737bf422127283c08e['h00692] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0034a] =  Ifd35529b44c957737bf422127283c08e['h00694] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0034b] =  Ifd35529b44c957737bf422127283c08e['h00696] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0034c] =  Ifd35529b44c957737bf422127283c08e['h00698] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0034d] =  Ifd35529b44c957737bf422127283c08e['h0069a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0034e] =  Ifd35529b44c957737bf422127283c08e['h0069c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0034f] =  Ifd35529b44c957737bf422127283c08e['h0069e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00350] =  Ifd35529b44c957737bf422127283c08e['h006a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00351] =  Ifd35529b44c957737bf422127283c08e['h006a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00352] =  Ifd35529b44c957737bf422127283c08e['h006a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00353] =  Ifd35529b44c957737bf422127283c08e['h006a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00354] =  Ifd35529b44c957737bf422127283c08e['h006a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00355] =  Ifd35529b44c957737bf422127283c08e['h006aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00356] =  Ifd35529b44c957737bf422127283c08e['h006ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00357] =  Ifd35529b44c957737bf422127283c08e['h006ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00358] =  Ifd35529b44c957737bf422127283c08e['h006b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00359] =  Ifd35529b44c957737bf422127283c08e['h006b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0035a] =  Ifd35529b44c957737bf422127283c08e['h006b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0035b] =  Ifd35529b44c957737bf422127283c08e['h006b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0035c] =  Ifd35529b44c957737bf422127283c08e['h006b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0035d] =  Ifd35529b44c957737bf422127283c08e['h006ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0035e] =  Ifd35529b44c957737bf422127283c08e['h006bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0035f] =  Ifd35529b44c957737bf422127283c08e['h006be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00360] =  Ifd35529b44c957737bf422127283c08e['h006c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00361] =  Ifd35529b44c957737bf422127283c08e['h006c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00362] =  Ifd35529b44c957737bf422127283c08e['h006c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00363] =  Ifd35529b44c957737bf422127283c08e['h006c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00364] =  Ifd35529b44c957737bf422127283c08e['h006c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00365] =  Ifd35529b44c957737bf422127283c08e['h006ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00366] =  Ifd35529b44c957737bf422127283c08e['h006cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00367] =  Ifd35529b44c957737bf422127283c08e['h006ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00368] =  Ifd35529b44c957737bf422127283c08e['h006d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00369] =  Ifd35529b44c957737bf422127283c08e['h006d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0036a] =  Ifd35529b44c957737bf422127283c08e['h006d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0036b] =  Ifd35529b44c957737bf422127283c08e['h006d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0036c] =  Ifd35529b44c957737bf422127283c08e['h006d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0036d] =  Ifd35529b44c957737bf422127283c08e['h006da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0036e] =  Ifd35529b44c957737bf422127283c08e['h006dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0036f] =  Ifd35529b44c957737bf422127283c08e['h006de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00370] =  Ifd35529b44c957737bf422127283c08e['h006e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00371] =  Ifd35529b44c957737bf422127283c08e['h006e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00372] =  Ifd35529b44c957737bf422127283c08e['h006e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00373] =  Ifd35529b44c957737bf422127283c08e['h006e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00374] =  Ifd35529b44c957737bf422127283c08e['h006e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00375] =  Ifd35529b44c957737bf422127283c08e['h006ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00376] =  Ifd35529b44c957737bf422127283c08e['h006ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00377] =  Ifd35529b44c957737bf422127283c08e['h006ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00378] =  Ifd35529b44c957737bf422127283c08e['h006f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00379] =  Ifd35529b44c957737bf422127283c08e['h006f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0037a] =  Ifd35529b44c957737bf422127283c08e['h006f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0037b] =  Ifd35529b44c957737bf422127283c08e['h006f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0037c] =  Ifd35529b44c957737bf422127283c08e['h006f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0037d] =  Ifd35529b44c957737bf422127283c08e['h006fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0037e] =  Ifd35529b44c957737bf422127283c08e['h006fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0037f] =  Ifd35529b44c957737bf422127283c08e['h006fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00380] =  Ifd35529b44c957737bf422127283c08e['h00700] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00381] =  Ifd35529b44c957737bf422127283c08e['h00702] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00382] =  Ifd35529b44c957737bf422127283c08e['h00704] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00383] =  Ifd35529b44c957737bf422127283c08e['h00706] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00384] =  Ifd35529b44c957737bf422127283c08e['h00708] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00385] =  Ifd35529b44c957737bf422127283c08e['h0070a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00386] =  Ifd35529b44c957737bf422127283c08e['h0070c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00387] =  Ifd35529b44c957737bf422127283c08e['h0070e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00388] =  Ifd35529b44c957737bf422127283c08e['h00710] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00389] =  Ifd35529b44c957737bf422127283c08e['h00712] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0038a] =  Ifd35529b44c957737bf422127283c08e['h00714] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0038b] =  Ifd35529b44c957737bf422127283c08e['h00716] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0038c] =  Ifd35529b44c957737bf422127283c08e['h00718] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0038d] =  Ifd35529b44c957737bf422127283c08e['h0071a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0038e] =  Ifd35529b44c957737bf422127283c08e['h0071c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0038f] =  Ifd35529b44c957737bf422127283c08e['h0071e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00390] =  Ifd35529b44c957737bf422127283c08e['h00720] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00391] =  Ifd35529b44c957737bf422127283c08e['h00722] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00392] =  Ifd35529b44c957737bf422127283c08e['h00724] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00393] =  Ifd35529b44c957737bf422127283c08e['h00726] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00394] =  Ifd35529b44c957737bf422127283c08e['h00728] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00395] =  Ifd35529b44c957737bf422127283c08e['h0072a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00396] =  Ifd35529b44c957737bf422127283c08e['h0072c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00397] =  Ifd35529b44c957737bf422127283c08e['h0072e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00398] =  Ifd35529b44c957737bf422127283c08e['h00730] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00399] =  Ifd35529b44c957737bf422127283c08e['h00732] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0039a] =  Ifd35529b44c957737bf422127283c08e['h00734] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0039b] =  Ifd35529b44c957737bf422127283c08e['h00736] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0039c] =  Ifd35529b44c957737bf422127283c08e['h00738] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0039d] =  Ifd35529b44c957737bf422127283c08e['h0073a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0039e] =  Ifd35529b44c957737bf422127283c08e['h0073c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0039f] =  Ifd35529b44c957737bf422127283c08e['h0073e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003a0] =  Ifd35529b44c957737bf422127283c08e['h00740] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003a1] =  Ifd35529b44c957737bf422127283c08e['h00742] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003a2] =  Ifd35529b44c957737bf422127283c08e['h00744] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003a3] =  Ifd35529b44c957737bf422127283c08e['h00746] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003a4] =  Ifd35529b44c957737bf422127283c08e['h00748] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003a5] =  Ifd35529b44c957737bf422127283c08e['h0074a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003a6] =  Ifd35529b44c957737bf422127283c08e['h0074c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003a7] =  Ifd35529b44c957737bf422127283c08e['h0074e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003a8] =  Ifd35529b44c957737bf422127283c08e['h00750] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003a9] =  Ifd35529b44c957737bf422127283c08e['h00752] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003aa] =  Ifd35529b44c957737bf422127283c08e['h00754] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003ab] =  Ifd35529b44c957737bf422127283c08e['h00756] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003ac] =  Ifd35529b44c957737bf422127283c08e['h00758] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003ad] =  Ifd35529b44c957737bf422127283c08e['h0075a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003ae] =  Ifd35529b44c957737bf422127283c08e['h0075c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003af] =  Ifd35529b44c957737bf422127283c08e['h0075e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003b0] =  Ifd35529b44c957737bf422127283c08e['h00760] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003b1] =  Ifd35529b44c957737bf422127283c08e['h00762] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003b2] =  Ifd35529b44c957737bf422127283c08e['h00764] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003b3] =  Ifd35529b44c957737bf422127283c08e['h00766] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003b4] =  Ifd35529b44c957737bf422127283c08e['h00768] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003b5] =  Ifd35529b44c957737bf422127283c08e['h0076a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003b6] =  Ifd35529b44c957737bf422127283c08e['h0076c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003b7] =  Ifd35529b44c957737bf422127283c08e['h0076e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003b8] =  Ifd35529b44c957737bf422127283c08e['h00770] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003b9] =  Ifd35529b44c957737bf422127283c08e['h00772] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003ba] =  Ifd35529b44c957737bf422127283c08e['h00774] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003bb] =  Ifd35529b44c957737bf422127283c08e['h00776] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003bc] =  Ifd35529b44c957737bf422127283c08e['h00778] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003bd] =  Ifd35529b44c957737bf422127283c08e['h0077a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003be] =  Ifd35529b44c957737bf422127283c08e['h0077c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003bf] =  Ifd35529b44c957737bf422127283c08e['h0077e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003c0] =  Ifd35529b44c957737bf422127283c08e['h00780] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003c1] =  Ifd35529b44c957737bf422127283c08e['h00782] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003c2] =  Ifd35529b44c957737bf422127283c08e['h00784] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003c3] =  Ifd35529b44c957737bf422127283c08e['h00786] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003c4] =  Ifd35529b44c957737bf422127283c08e['h00788] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003c5] =  Ifd35529b44c957737bf422127283c08e['h0078a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003c6] =  Ifd35529b44c957737bf422127283c08e['h0078c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003c7] =  Ifd35529b44c957737bf422127283c08e['h0078e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003c8] =  Ifd35529b44c957737bf422127283c08e['h00790] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003c9] =  Ifd35529b44c957737bf422127283c08e['h00792] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003ca] =  Ifd35529b44c957737bf422127283c08e['h00794] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003cb] =  Ifd35529b44c957737bf422127283c08e['h00796] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003cc] =  Ifd35529b44c957737bf422127283c08e['h00798] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003cd] =  Ifd35529b44c957737bf422127283c08e['h0079a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003ce] =  Ifd35529b44c957737bf422127283c08e['h0079c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003cf] =  Ifd35529b44c957737bf422127283c08e['h0079e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003d0] =  Ifd35529b44c957737bf422127283c08e['h007a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003d1] =  Ifd35529b44c957737bf422127283c08e['h007a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003d2] =  Ifd35529b44c957737bf422127283c08e['h007a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003d3] =  Ifd35529b44c957737bf422127283c08e['h007a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003d4] =  Ifd35529b44c957737bf422127283c08e['h007a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003d5] =  Ifd35529b44c957737bf422127283c08e['h007aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003d6] =  Ifd35529b44c957737bf422127283c08e['h007ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003d7] =  Ifd35529b44c957737bf422127283c08e['h007ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003d8] =  Ifd35529b44c957737bf422127283c08e['h007b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003d9] =  Ifd35529b44c957737bf422127283c08e['h007b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003da] =  Ifd35529b44c957737bf422127283c08e['h007b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003db] =  Ifd35529b44c957737bf422127283c08e['h007b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003dc] =  Ifd35529b44c957737bf422127283c08e['h007b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003dd] =  Ifd35529b44c957737bf422127283c08e['h007ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003de] =  Ifd35529b44c957737bf422127283c08e['h007bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003df] =  Ifd35529b44c957737bf422127283c08e['h007be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003e0] =  Ifd35529b44c957737bf422127283c08e['h007c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003e1] =  Ifd35529b44c957737bf422127283c08e['h007c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003e2] =  Ifd35529b44c957737bf422127283c08e['h007c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003e3] =  Ifd35529b44c957737bf422127283c08e['h007c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003e4] =  Ifd35529b44c957737bf422127283c08e['h007c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003e5] =  Ifd35529b44c957737bf422127283c08e['h007ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003e6] =  Ifd35529b44c957737bf422127283c08e['h007cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003e7] =  Ifd35529b44c957737bf422127283c08e['h007ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003e8] =  Ifd35529b44c957737bf422127283c08e['h007d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003e9] =  Ifd35529b44c957737bf422127283c08e['h007d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003ea] =  Ifd35529b44c957737bf422127283c08e['h007d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003eb] =  Ifd35529b44c957737bf422127283c08e['h007d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003ec] =  Ifd35529b44c957737bf422127283c08e['h007d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003ed] =  Ifd35529b44c957737bf422127283c08e['h007da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003ee] =  Ifd35529b44c957737bf422127283c08e['h007dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003ef] =  Ifd35529b44c957737bf422127283c08e['h007de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003f0] =  Ifd35529b44c957737bf422127283c08e['h007e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003f1] =  Ifd35529b44c957737bf422127283c08e['h007e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003f2] =  Ifd35529b44c957737bf422127283c08e['h007e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003f3] =  Ifd35529b44c957737bf422127283c08e['h007e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003f4] =  Ifd35529b44c957737bf422127283c08e['h007e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003f5] =  Ifd35529b44c957737bf422127283c08e['h007ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003f6] =  Ifd35529b44c957737bf422127283c08e['h007ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003f7] =  Ifd35529b44c957737bf422127283c08e['h007ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003f8] =  Ifd35529b44c957737bf422127283c08e['h007f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003f9] =  Ifd35529b44c957737bf422127283c08e['h007f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003fa] =  Ifd35529b44c957737bf422127283c08e['h007f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003fb] =  Ifd35529b44c957737bf422127283c08e['h007f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003fc] =  Ifd35529b44c957737bf422127283c08e['h007f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003fd] =  Ifd35529b44c957737bf422127283c08e['h007fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003fe] =  Ifd35529b44c957737bf422127283c08e['h007fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h003ff] =  Ifd35529b44c957737bf422127283c08e['h007fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00400] =  Ifd35529b44c957737bf422127283c08e['h00800] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00401] =  Ifd35529b44c957737bf422127283c08e['h00802] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00402] =  Ifd35529b44c957737bf422127283c08e['h00804] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00403] =  Ifd35529b44c957737bf422127283c08e['h00806] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00404] =  Ifd35529b44c957737bf422127283c08e['h00808] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00405] =  Ifd35529b44c957737bf422127283c08e['h0080a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00406] =  Ifd35529b44c957737bf422127283c08e['h0080c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00407] =  Ifd35529b44c957737bf422127283c08e['h0080e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00408] =  Ifd35529b44c957737bf422127283c08e['h00810] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00409] =  Ifd35529b44c957737bf422127283c08e['h00812] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0040a] =  Ifd35529b44c957737bf422127283c08e['h00814] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0040b] =  Ifd35529b44c957737bf422127283c08e['h00816] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0040c] =  Ifd35529b44c957737bf422127283c08e['h00818] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0040d] =  Ifd35529b44c957737bf422127283c08e['h0081a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0040e] =  Ifd35529b44c957737bf422127283c08e['h0081c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0040f] =  Ifd35529b44c957737bf422127283c08e['h0081e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00410] =  Ifd35529b44c957737bf422127283c08e['h00820] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00411] =  Ifd35529b44c957737bf422127283c08e['h00822] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00412] =  Ifd35529b44c957737bf422127283c08e['h00824] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00413] =  Ifd35529b44c957737bf422127283c08e['h00826] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00414] =  Ifd35529b44c957737bf422127283c08e['h00828] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00415] =  Ifd35529b44c957737bf422127283c08e['h0082a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00416] =  Ifd35529b44c957737bf422127283c08e['h0082c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00417] =  Ifd35529b44c957737bf422127283c08e['h0082e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00418] =  Ifd35529b44c957737bf422127283c08e['h00830] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00419] =  Ifd35529b44c957737bf422127283c08e['h00832] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0041a] =  Ifd35529b44c957737bf422127283c08e['h00834] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0041b] =  Ifd35529b44c957737bf422127283c08e['h00836] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0041c] =  Ifd35529b44c957737bf422127283c08e['h00838] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0041d] =  Ifd35529b44c957737bf422127283c08e['h0083a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0041e] =  Ifd35529b44c957737bf422127283c08e['h0083c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0041f] =  Ifd35529b44c957737bf422127283c08e['h0083e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00420] =  Ifd35529b44c957737bf422127283c08e['h00840] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00421] =  Ifd35529b44c957737bf422127283c08e['h00842] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00422] =  Ifd35529b44c957737bf422127283c08e['h00844] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00423] =  Ifd35529b44c957737bf422127283c08e['h00846] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00424] =  Ifd35529b44c957737bf422127283c08e['h00848] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00425] =  Ifd35529b44c957737bf422127283c08e['h0084a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00426] =  Ifd35529b44c957737bf422127283c08e['h0084c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00427] =  Ifd35529b44c957737bf422127283c08e['h0084e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00428] =  Ifd35529b44c957737bf422127283c08e['h00850] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00429] =  Ifd35529b44c957737bf422127283c08e['h00852] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0042a] =  Ifd35529b44c957737bf422127283c08e['h00854] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0042b] =  Ifd35529b44c957737bf422127283c08e['h00856] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0042c] =  Ifd35529b44c957737bf422127283c08e['h00858] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0042d] =  Ifd35529b44c957737bf422127283c08e['h0085a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0042e] =  Ifd35529b44c957737bf422127283c08e['h0085c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0042f] =  Ifd35529b44c957737bf422127283c08e['h0085e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00430] =  Ifd35529b44c957737bf422127283c08e['h00860] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00431] =  Ifd35529b44c957737bf422127283c08e['h00862] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00432] =  Ifd35529b44c957737bf422127283c08e['h00864] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00433] =  Ifd35529b44c957737bf422127283c08e['h00866] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00434] =  Ifd35529b44c957737bf422127283c08e['h00868] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00435] =  Ifd35529b44c957737bf422127283c08e['h0086a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00436] =  Ifd35529b44c957737bf422127283c08e['h0086c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00437] =  Ifd35529b44c957737bf422127283c08e['h0086e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00438] =  Ifd35529b44c957737bf422127283c08e['h00870] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00439] =  Ifd35529b44c957737bf422127283c08e['h00872] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0043a] =  Ifd35529b44c957737bf422127283c08e['h00874] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0043b] =  Ifd35529b44c957737bf422127283c08e['h00876] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0043c] =  Ifd35529b44c957737bf422127283c08e['h00878] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0043d] =  Ifd35529b44c957737bf422127283c08e['h0087a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0043e] =  Ifd35529b44c957737bf422127283c08e['h0087c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0043f] =  Ifd35529b44c957737bf422127283c08e['h0087e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00440] =  Ifd35529b44c957737bf422127283c08e['h00880] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00441] =  Ifd35529b44c957737bf422127283c08e['h00882] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00442] =  Ifd35529b44c957737bf422127283c08e['h00884] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00443] =  Ifd35529b44c957737bf422127283c08e['h00886] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00444] =  Ifd35529b44c957737bf422127283c08e['h00888] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00445] =  Ifd35529b44c957737bf422127283c08e['h0088a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00446] =  Ifd35529b44c957737bf422127283c08e['h0088c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00447] =  Ifd35529b44c957737bf422127283c08e['h0088e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00448] =  Ifd35529b44c957737bf422127283c08e['h00890] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00449] =  Ifd35529b44c957737bf422127283c08e['h00892] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0044a] =  Ifd35529b44c957737bf422127283c08e['h00894] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0044b] =  Ifd35529b44c957737bf422127283c08e['h00896] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0044c] =  Ifd35529b44c957737bf422127283c08e['h00898] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0044d] =  Ifd35529b44c957737bf422127283c08e['h0089a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0044e] =  Ifd35529b44c957737bf422127283c08e['h0089c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0044f] =  Ifd35529b44c957737bf422127283c08e['h0089e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00450] =  Ifd35529b44c957737bf422127283c08e['h008a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00451] =  Ifd35529b44c957737bf422127283c08e['h008a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00452] =  Ifd35529b44c957737bf422127283c08e['h008a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00453] =  Ifd35529b44c957737bf422127283c08e['h008a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00454] =  Ifd35529b44c957737bf422127283c08e['h008a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00455] =  Ifd35529b44c957737bf422127283c08e['h008aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00456] =  Ifd35529b44c957737bf422127283c08e['h008ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00457] =  Ifd35529b44c957737bf422127283c08e['h008ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00458] =  Ifd35529b44c957737bf422127283c08e['h008b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00459] =  Ifd35529b44c957737bf422127283c08e['h008b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0045a] =  Ifd35529b44c957737bf422127283c08e['h008b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0045b] =  Ifd35529b44c957737bf422127283c08e['h008b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0045c] =  Ifd35529b44c957737bf422127283c08e['h008b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0045d] =  Ifd35529b44c957737bf422127283c08e['h008ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0045e] =  Ifd35529b44c957737bf422127283c08e['h008bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0045f] =  Ifd35529b44c957737bf422127283c08e['h008be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00460] =  Ifd35529b44c957737bf422127283c08e['h008c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00461] =  Ifd35529b44c957737bf422127283c08e['h008c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00462] =  Ifd35529b44c957737bf422127283c08e['h008c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00463] =  Ifd35529b44c957737bf422127283c08e['h008c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00464] =  Ifd35529b44c957737bf422127283c08e['h008c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00465] =  Ifd35529b44c957737bf422127283c08e['h008ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00466] =  Ifd35529b44c957737bf422127283c08e['h008cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00467] =  Ifd35529b44c957737bf422127283c08e['h008ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00468] =  Ifd35529b44c957737bf422127283c08e['h008d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00469] =  Ifd35529b44c957737bf422127283c08e['h008d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0046a] =  Ifd35529b44c957737bf422127283c08e['h008d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0046b] =  Ifd35529b44c957737bf422127283c08e['h008d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0046c] =  Ifd35529b44c957737bf422127283c08e['h008d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0046d] =  Ifd35529b44c957737bf422127283c08e['h008da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0046e] =  Ifd35529b44c957737bf422127283c08e['h008dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0046f] =  Ifd35529b44c957737bf422127283c08e['h008de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00470] =  Ifd35529b44c957737bf422127283c08e['h008e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00471] =  Ifd35529b44c957737bf422127283c08e['h008e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00472] =  Ifd35529b44c957737bf422127283c08e['h008e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00473] =  Ifd35529b44c957737bf422127283c08e['h008e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00474] =  Ifd35529b44c957737bf422127283c08e['h008e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00475] =  Ifd35529b44c957737bf422127283c08e['h008ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00476] =  Ifd35529b44c957737bf422127283c08e['h008ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00477] =  Ifd35529b44c957737bf422127283c08e['h008ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00478] =  Ifd35529b44c957737bf422127283c08e['h008f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00479] =  Ifd35529b44c957737bf422127283c08e['h008f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0047a] =  Ifd35529b44c957737bf422127283c08e['h008f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0047b] =  Ifd35529b44c957737bf422127283c08e['h008f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0047c] =  Ifd35529b44c957737bf422127283c08e['h008f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0047d] =  Ifd35529b44c957737bf422127283c08e['h008fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0047e] =  Ifd35529b44c957737bf422127283c08e['h008fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0047f] =  Ifd35529b44c957737bf422127283c08e['h008fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00480] =  Ifd35529b44c957737bf422127283c08e['h00900] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00481] =  Ifd35529b44c957737bf422127283c08e['h00902] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00482] =  Ifd35529b44c957737bf422127283c08e['h00904] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00483] =  Ifd35529b44c957737bf422127283c08e['h00906] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00484] =  Ifd35529b44c957737bf422127283c08e['h00908] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00485] =  Ifd35529b44c957737bf422127283c08e['h0090a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00486] =  Ifd35529b44c957737bf422127283c08e['h0090c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00487] =  Ifd35529b44c957737bf422127283c08e['h0090e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00488] =  Ifd35529b44c957737bf422127283c08e['h00910] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00489] =  Ifd35529b44c957737bf422127283c08e['h00912] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0048a] =  Ifd35529b44c957737bf422127283c08e['h00914] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0048b] =  Ifd35529b44c957737bf422127283c08e['h00916] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0048c] =  Ifd35529b44c957737bf422127283c08e['h00918] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0048d] =  Ifd35529b44c957737bf422127283c08e['h0091a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0048e] =  Ifd35529b44c957737bf422127283c08e['h0091c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0048f] =  Ifd35529b44c957737bf422127283c08e['h0091e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00490] =  Ifd35529b44c957737bf422127283c08e['h00920] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00491] =  Ifd35529b44c957737bf422127283c08e['h00922] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00492] =  Ifd35529b44c957737bf422127283c08e['h00924] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00493] =  Ifd35529b44c957737bf422127283c08e['h00926] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00494] =  Ifd35529b44c957737bf422127283c08e['h00928] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00495] =  Ifd35529b44c957737bf422127283c08e['h0092a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00496] =  Ifd35529b44c957737bf422127283c08e['h0092c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00497] =  Ifd35529b44c957737bf422127283c08e['h0092e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00498] =  Ifd35529b44c957737bf422127283c08e['h00930] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00499] =  Ifd35529b44c957737bf422127283c08e['h00932] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0049a] =  Ifd35529b44c957737bf422127283c08e['h00934] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0049b] =  Ifd35529b44c957737bf422127283c08e['h00936] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0049c] =  Ifd35529b44c957737bf422127283c08e['h00938] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0049d] =  Ifd35529b44c957737bf422127283c08e['h0093a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0049e] =  Ifd35529b44c957737bf422127283c08e['h0093c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0049f] =  Ifd35529b44c957737bf422127283c08e['h0093e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004a0] =  Ifd35529b44c957737bf422127283c08e['h00940] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004a1] =  Ifd35529b44c957737bf422127283c08e['h00942] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004a2] =  Ifd35529b44c957737bf422127283c08e['h00944] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004a3] =  Ifd35529b44c957737bf422127283c08e['h00946] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004a4] =  Ifd35529b44c957737bf422127283c08e['h00948] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004a5] =  Ifd35529b44c957737bf422127283c08e['h0094a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004a6] =  Ifd35529b44c957737bf422127283c08e['h0094c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004a7] =  Ifd35529b44c957737bf422127283c08e['h0094e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004a8] =  Ifd35529b44c957737bf422127283c08e['h00950] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004a9] =  Ifd35529b44c957737bf422127283c08e['h00952] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004aa] =  Ifd35529b44c957737bf422127283c08e['h00954] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004ab] =  Ifd35529b44c957737bf422127283c08e['h00956] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004ac] =  Ifd35529b44c957737bf422127283c08e['h00958] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004ad] =  Ifd35529b44c957737bf422127283c08e['h0095a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004ae] =  Ifd35529b44c957737bf422127283c08e['h0095c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004af] =  Ifd35529b44c957737bf422127283c08e['h0095e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004b0] =  Ifd35529b44c957737bf422127283c08e['h00960] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004b1] =  Ifd35529b44c957737bf422127283c08e['h00962] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004b2] =  Ifd35529b44c957737bf422127283c08e['h00964] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004b3] =  Ifd35529b44c957737bf422127283c08e['h00966] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004b4] =  Ifd35529b44c957737bf422127283c08e['h00968] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004b5] =  Ifd35529b44c957737bf422127283c08e['h0096a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004b6] =  Ifd35529b44c957737bf422127283c08e['h0096c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004b7] =  Ifd35529b44c957737bf422127283c08e['h0096e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004b8] =  Ifd35529b44c957737bf422127283c08e['h00970] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004b9] =  Ifd35529b44c957737bf422127283c08e['h00972] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004ba] =  Ifd35529b44c957737bf422127283c08e['h00974] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004bb] =  Ifd35529b44c957737bf422127283c08e['h00976] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004bc] =  Ifd35529b44c957737bf422127283c08e['h00978] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004bd] =  Ifd35529b44c957737bf422127283c08e['h0097a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004be] =  Ifd35529b44c957737bf422127283c08e['h0097c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004bf] =  Ifd35529b44c957737bf422127283c08e['h0097e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004c0] =  Ifd35529b44c957737bf422127283c08e['h00980] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004c1] =  Ifd35529b44c957737bf422127283c08e['h00982] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004c2] =  Ifd35529b44c957737bf422127283c08e['h00984] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004c3] =  Ifd35529b44c957737bf422127283c08e['h00986] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004c4] =  Ifd35529b44c957737bf422127283c08e['h00988] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004c5] =  Ifd35529b44c957737bf422127283c08e['h0098a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004c6] =  Ifd35529b44c957737bf422127283c08e['h0098c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004c7] =  Ifd35529b44c957737bf422127283c08e['h0098e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004c8] =  Ifd35529b44c957737bf422127283c08e['h00990] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004c9] =  Ifd35529b44c957737bf422127283c08e['h00992] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004ca] =  Ifd35529b44c957737bf422127283c08e['h00994] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004cb] =  Ifd35529b44c957737bf422127283c08e['h00996] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004cc] =  Ifd35529b44c957737bf422127283c08e['h00998] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004cd] =  Ifd35529b44c957737bf422127283c08e['h0099a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004ce] =  Ifd35529b44c957737bf422127283c08e['h0099c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004cf] =  Ifd35529b44c957737bf422127283c08e['h0099e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004d0] =  Ifd35529b44c957737bf422127283c08e['h009a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004d1] =  Ifd35529b44c957737bf422127283c08e['h009a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004d2] =  Ifd35529b44c957737bf422127283c08e['h009a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004d3] =  Ifd35529b44c957737bf422127283c08e['h009a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004d4] =  Ifd35529b44c957737bf422127283c08e['h009a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004d5] =  Ifd35529b44c957737bf422127283c08e['h009aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004d6] =  Ifd35529b44c957737bf422127283c08e['h009ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004d7] =  Ifd35529b44c957737bf422127283c08e['h009ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004d8] =  Ifd35529b44c957737bf422127283c08e['h009b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004d9] =  Ifd35529b44c957737bf422127283c08e['h009b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004da] =  Ifd35529b44c957737bf422127283c08e['h009b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004db] =  Ifd35529b44c957737bf422127283c08e['h009b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004dc] =  Ifd35529b44c957737bf422127283c08e['h009b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004dd] =  Ifd35529b44c957737bf422127283c08e['h009ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004de] =  Ifd35529b44c957737bf422127283c08e['h009bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004df] =  Ifd35529b44c957737bf422127283c08e['h009be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004e0] =  Ifd35529b44c957737bf422127283c08e['h009c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004e1] =  Ifd35529b44c957737bf422127283c08e['h009c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004e2] =  Ifd35529b44c957737bf422127283c08e['h009c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004e3] =  Ifd35529b44c957737bf422127283c08e['h009c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004e4] =  Ifd35529b44c957737bf422127283c08e['h009c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004e5] =  Ifd35529b44c957737bf422127283c08e['h009ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004e6] =  Ifd35529b44c957737bf422127283c08e['h009cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004e7] =  Ifd35529b44c957737bf422127283c08e['h009ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004e8] =  Ifd35529b44c957737bf422127283c08e['h009d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004e9] =  Ifd35529b44c957737bf422127283c08e['h009d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004ea] =  Ifd35529b44c957737bf422127283c08e['h009d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004eb] =  Ifd35529b44c957737bf422127283c08e['h009d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004ec] =  Ifd35529b44c957737bf422127283c08e['h009d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004ed] =  Ifd35529b44c957737bf422127283c08e['h009da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004ee] =  Ifd35529b44c957737bf422127283c08e['h009dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004ef] =  Ifd35529b44c957737bf422127283c08e['h009de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004f0] =  Ifd35529b44c957737bf422127283c08e['h009e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004f1] =  Ifd35529b44c957737bf422127283c08e['h009e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004f2] =  Ifd35529b44c957737bf422127283c08e['h009e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004f3] =  Ifd35529b44c957737bf422127283c08e['h009e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004f4] =  Ifd35529b44c957737bf422127283c08e['h009e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004f5] =  Ifd35529b44c957737bf422127283c08e['h009ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004f6] =  Ifd35529b44c957737bf422127283c08e['h009ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004f7] =  Ifd35529b44c957737bf422127283c08e['h009ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004f8] =  Ifd35529b44c957737bf422127283c08e['h009f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004f9] =  Ifd35529b44c957737bf422127283c08e['h009f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004fa] =  Ifd35529b44c957737bf422127283c08e['h009f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004fb] =  Ifd35529b44c957737bf422127283c08e['h009f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004fc] =  Ifd35529b44c957737bf422127283c08e['h009f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004fd] =  Ifd35529b44c957737bf422127283c08e['h009fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004fe] =  Ifd35529b44c957737bf422127283c08e['h009fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h004ff] =  Ifd35529b44c957737bf422127283c08e['h009fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00500] =  Ifd35529b44c957737bf422127283c08e['h00a00] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00501] =  Ifd35529b44c957737bf422127283c08e['h00a02] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00502] =  Ifd35529b44c957737bf422127283c08e['h00a04] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00503] =  Ifd35529b44c957737bf422127283c08e['h00a06] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00504] =  Ifd35529b44c957737bf422127283c08e['h00a08] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00505] =  Ifd35529b44c957737bf422127283c08e['h00a0a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00506] =  Ifd35529b44c957737bf422127283c08e['h00a0c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00507] =  Ifd35529b44c957737bf422127283c08e['h00a0e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00508] =  Ifd35529b44c957737bf422127283c08e['h00a10] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00509] =  Ifd35529b44c957737bf422127283c08e['h00a12] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0050a] =  Ifd35529b44c957737bf422127283c08e['h00a14] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0050b] =  Ifd35529b44c957737bf422127283c08e['h00a16] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0050c] =  Ifd35529b44c957737bf422127283c08e['h00a18] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0050d] =  Ifd35529b44c957737bf422127283c08e['h00a1a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0050e] =  Ifd35529b44c957737bf422127283c08e['h00a1c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0050f] =  Ifd35529b44c957737bf422127283c08e['h00a1e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00510] =  Ifd35529b44c957737bf422127283c08e['h00a20] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00511] =  Ifd35529b44c957737bf422127283c08e['h00a22] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00512] =  Ifd35529b44c957737bf422127283c08e['h00a24] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00513] =  Ifd35529b44c957737bf422127283c08e['h00a26] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00514] =  Ifd35529b44c957737bf422127283c08e['h00a28] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00515] =  Ifd35529b44c957737bf422127283c08e['h00a2a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00516] =  Ifd35529b44c957737bf422127283c08e['h00a2c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00517] =  Ifd35529b44c957737bf422127283c08e['h00a2e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00518] =  Ifd35529b44c957737bf422127283c08e['h00a30] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00519] =  Ifd35529b44c957737bf422127283c08e['h00a32] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0051a] =  Ifd35529b44c957737bf422127283c08e['h00a34] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0051b] =  Ifd35529b44c957737bf422127283c08e['h00a36] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0051c] =  Ifd35529b44c957737bf422127283c08e['h00a38] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0051d] =  Ifd35529b44c957737bf422127283c08e['h00a3a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0051e] =  Ifd35529b44c957737bf422127283c08e['h00a3c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0051f] =  Ifd35529b44c957737bf422127283c08e['h00a3e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00520] =  Ifd35529b44c957737bf422127283c08e['h00a40] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00521] =  Ifd35529b44c957737bf422127283c08e['h00a42] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00522] =  Ifd35529b44c957737bf422127283c08e['h00a44] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00523] =  Ifd35529b44c957737bf422127283c08e['h00a46] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00524] =  Ifd35529b44c957737bf422127283c08e['h00a48] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00525] =  Ifd35529b44c957737bf422127283c08e['h00a4a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00526] =  Ifd35529b44c957737bf422127283c08e['h00a4c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00527] =  Ifd35529b44c957737bf422127283c08e['h00a4e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00528] =  Ifd35529b44c957737bf422127283c08e['h00a50] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00529] =  Ifd35529b44c957737bf422127283c08e['h00a52] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0052a] =  Ifd35529b44c957737bf422127283c08e['h00a54] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0052b] =  Ifd35529b44c957737bf422127283c08e['h00a56] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0052c] =  Ifd35529b44c957737bf422127283c08e['h00a58] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0052d] =  Ifd35529b44c957737bf422127283c08e['h00a5a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0052e] =  Ifd35529b44c957737bf422127283c08e['h00a5c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0052f] =  Ifd35529b44c957737bf422127283c08e['h00a5e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00530] =  Ifd35529b44c957737bf422127283c08e['h00a60] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00531] =  Ifd35529b44c957737bf422127283c08e['h00a62] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00532] =  Ifd35529b44c957737bf422127283c08e['h00a64] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00533] =  Ifd35529b44c957737bf422127283c08e['h00a66] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00534] =  Ifd35529b44c957737bf422127283c08e['h00a68] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00535] =  Ifd35529b44c957737bf422127283c08e['h00a6a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00536] =  Ifd35529b44c957737bf422127283c08e['h00a6c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00537] =  Ifd35529b44c957737bf422127283c08e['h00a6e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00538] =  Ifd35529b44c957737bf422127283c08e['h00a70] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00539] =  Ifd35529b44c957737bf422127283c08e['h00a72] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0053a] =  Ifd35529b44c957737bf422127283c08e['h00a74] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0053b] =  Ifd35529b44c957737bf422127283c08e['h00a76] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0053c] =  Ifd35529b44c957737bf422127283c08e['h00a78] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0053d] =  Ifd35529b44c957737bf422127283c08e['h00a7a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0053e] =  Ifd35529b44c957737bf422127283c08e['h00a7c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0053f] =  Ifd35529b44c957737bf422127283c08e['h00a7e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00540] =  Ifd35529b44c957737bf422127283c08e['h00a80] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00541] =  Ifd35529b44c957737bf422127283c08e['h00a82] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00542] =  Ifd35529b44c957737bf422127283c08e['h00a84] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00543] =  Ifd35529b44c957737bf422127283c08e['h00a86] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00544] =  Ifd35529b44c957737bf422127283c08e['h00a88] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00545] =  Ifd35529b44c957737bf422127283c08e['h00a8a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00546] =  Ifd35529b44c957737bf422127283c08e['h00a8c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00547] =  Ifd35529b44c957737bf422127283c08e['h00a8e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00548] =  Ifd35529b44c957737bf422127283c08e['h00a90] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00549] =  Ifd35529b44c957737bf422127283c08e['h00a92] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0054a] =  Ifd35529b44c957737bf422127283c08e['h00a94] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0054b] =  Ifd35529b44c957737bf422127283c08e['h00a96] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0054c] =  Ifd35529b44c957737bf422127283c08e['h00a98] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0054d] =  Ifd35529b44c957737bf422127283c08e['h00a9a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0054e] =  Ifd35529b44c957737bf422127283c08e['h00a9c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0054f] =  Ifd35529b44c957737bf422127283c08e['h00a9e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00550] =  Ifd35529b44c957737bf422127283c08e['h00aa0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00551] =  Ifd35529b44c957737bf422127283c08e['h00aa2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00552] =  Ifd35529b44c957737bf422127283c08e['h00aa4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00553] =  Ifd35529b44c957737bf422127283c08e['h00aa6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00554] =  Ifd35529b44c957737bf422127283c08e['h00aa8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00555] =  Ifd35529b44c957737bf422127283c08e['h00aaa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00556] =  Ifd35529b44c957737bf422127283c08e['h00aac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00557] =  Ifd35529b44c957737bf422127283c08e['h00aae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00558] =  Ifd35529b44c957737bf422127283c08e['h00ab0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00559] =  Ifd35529b44c957737bf422127283c08e['h00ab2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0055a] =  Ifd35529b44c957737bf422127283c08e['h00ab4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0055b] =  Ifd35529b44c957737bf422127283c08e['h00ab6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0055c] =  Ifd35529b44c957737bf422127283c08e['h00ab8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0055d] =  Ifd35529b44c957737bf422127283c08e['h00aba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0055e] =  Ifd35529b44c957737bf422127283c08e['h00abc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0055f] =  Ifd35529b44c957737bf422127283c08e['h00abe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00560] =  Ifd35529b44c957737bf422127283c08e['h00ac0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00561] =  Ifd35529b44c957737bf422127283c08e['h00ac2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00562] =  Ifd35529b44c957737bf422127283c08e['h00ac4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00563] =  Ifd35529b44c957737bf422127283c08e['h00ac6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00564] =  Ifd35529b44c957737bf422127283c08e['h00ac8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00565] =  Ifd35529b44c957737bf422127283c08e['h00aca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00566] =  Ifd35529b44c957737bf422127283c08e['h00acc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00567] =  Ifd35529b44c957737bf422127283c08e['h00ace] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00568] =  Ifd35529b44c957737bf422127283c08e['h00ad0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00569] =  Ifd35529b44c957737bf422127283c08e['h00ad2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0056a] =  Ifd35529b44c957737bf422127283c08e['h00ad4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0056b] =  Ifd35529b44c957737bf422127283c08e['h00ad6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0056c] =  Ifd35529b44c957737bf422127283c08e['h00ad8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0056d] =  Ifd35529b44c957737bf422127283c08e['h00ada] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0056e] =  Ifd35529b44c957737bf422127283c08e['h00adc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0056f] =  Ifd35529b44c957737bf422127283c08e['h00ade] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00570] =  Ifd35529b44c957737bf422127283c08e['h00ae0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00571] =  Ifd35529b44c957737bf422127283c08e['h00ae2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00572] =  Ifd35529b44c957737bf422127283c08e['h00ae4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00573] =  Ifd35529b44c957737bf422127283c08e['h00ae6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00574] =  Ifd35529b44c957737bf422127283c08e['h00ae8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00575] =  Ifd35529b44c957737bf422127283c08e['h00aea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00576] =  Ifd35529b44c957737bf422127283c08e['h00aec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00577] =  Ifd35529b44c957737bf422127283c08e['h00aee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00578] =  Ifd35529b44c957737bf422127283c08e['h00af0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00579] =  Ifd35529b44c957737bf422127283c08e['h00af2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0057a] =  Ifd35529b44c957737bf422127283c08e['h00af4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0057b] =  Ifd35529b44c957737bf422127283c08e['h00af6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0057c] =  Ifd35529b44c957737bf422127283c08e['h00af8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0057d] =  Ifd35529b44c957737bf422127283c08e['h00afa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0057e] =  Ifd35529b44c957737bf422127283c08e['h00afc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0057f] =  Ifd35529b44c957737bf422127283c08e['h00afe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00580] =  Ifd35529b44c957737bf422127283c08e['h00b00] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00581] =  Ifd35529b44c957737bf422127283c08e['h00b02] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00582] =  Ifd35529b44c957737bf422127283c08e['h00b04] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00583] =  Ifd35529b44c957737bf422127283c08e['h00b06] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00584] =  Ifd35529b44c957737bf422127283c08e['h00b08] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00585] =  Ifd35529b44c957737bf422127283c08e['h00b0a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00586] =  Ifd35529b44c957737bf422127283c08e['h00b0c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00587] =  Ifd35529b44c957737bf422127283c08e['h00b0e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00588] =  Ifd35529b44c957737bf422127283c08e['h00b10] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00589] =  Ifd35529b44c957737bf422127283c08e['h00b12] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0058a] =  Ifd35529b44c957737bf422127283c08e['h00b14] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0058b] =  Ifd35529b44c957737bf422127283c08e['h00b16] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0058c] =  Ifd35529b44c957737bf422127283c08e['h00b18] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0058d] =  Ifd35529b44c957737bf422127283c08e['h00b1a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0058e] =  Ifd35529b44c957737bf422127283c08e['h00b1c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0058f] =  Ifd35529b44c957737bf422127283c08e['h00b1e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00590] =  Ifd35529b44c957737bf422127283c08e['h00b20] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00591] =  Ifd35529b44c957737bf422127283c08e['h00b22] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00592] =  Ifd35529b44c957737bf422127283c08e['h00b24] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00593] =  Ifd35529b44c957737bf422127283c08e['h00b26] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00594] =  Ifd35529b44c957737bf422127283c08e['h00b28] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00595] =  Ifd35529b44c957737bf422127283c08e['h00b2a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00596] =  Ifd35529b44c957737bf422127283c08e['h00b2c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00597] =  Ifd35529b44c957737bf422127283c08e['h00b2e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00598] =  Ifd35529b44c957737bf422127283c08e['h00b30] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00599] =  Ifd35529b44c957737bf422127283c08e['h00b32] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0059a] =  Ifd35529b44c957737bf422127283c08e['h00b34] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0059b] =  Ifd35529b44c957737bf422127283c08e['h00b36] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0059c] =  Ifd35529b44c957737bf422127283c08e['h00b38] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0059d] =  Ifd35529b44c957737bf422127283c08e['h00b3a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0059e] =  Ifd35529b44c957737bf422127283c08e['h00b3c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0059f] =  Ifd35529b44c957737bf422127283c08e['h00b3e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005a0] =  Ifd35529b44c957737bf422127283c08e['h00b40] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005a1] =  Ifd35529b44c957737bf422127283c08e['h00b42] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005a2] =  Ifd35529b44c957737bf422127283c08e['h00b44] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005a3] =  Ifd35529b44c957737bf422127283c08e['h00b46] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005a4] =  Ifd35529b44c957737bf422127283c08e['h00b48] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005a5] =  Ifd35529b44c957737bf422127283c08e['h00b4a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005a6] =  Ifd35529b44c957737bf422127283c08e['h00b4c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005a7] =  Ifd35529b44c957737bf422127283c08e['h00b4e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005a8] =  Ifd35529b44c957737bf422127283c08e['h00b50] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005a9] =  Ifd35529b44c957737bf422127283c08e['h00b52] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005aa] =  Ifd35529b44c957737bf422127283c08e['h00b54] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005ab] =  Ifd35529b44c957737bf422127283c08e['h00b56] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005ac] =  Ifd35529b44c957737bf422127283c08e['h00b58] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005ad] =  Ifd35529b44c957737bf422127283c08e['h00b5a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005ae] =  Ifd35529b44c957737bf422127283c08e['h00b5c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005af] =  Ifd35529b44c957737bf422127283c08e['h00b5e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005b0] =  Ifd35529b44c957737bf422127283c08e['h00b60] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005b1] =  Ifd35529b44c957737bf422127283c08e['h00b62] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005b2] =  Ifd35529b44c957737bf422127283c08e['h00b64] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005b3] =  Ifd35529b44c957737bf422127283c08e['h00b66] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005b4] =  Ifd35529b44c957737bf422127283c08e['h00b68] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005b5] =  Ifd35529b44c957737bf422127283c08e['h00b6a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005b6] =  Ifd35529b44c957737bf422127283c08e['h00b6c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005b7] =  Ifd35529b44c957737bf422127283c08e['h00b6e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005b8] =  Ifd35529b44c957737bf422127283c08e['h00b70] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005b9] =  Ifd35529b44c957737bf422127283c08e['h00b72] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005ba] =  Ifd35529b44c957737bf422127283c08e['h00b74] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005bb] =  Ifd35529b44c957737bf422127283c08e['h00b76] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005bc] =  Ifd35529b44c957737bf422127283c08e['h00b78] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005bd] =  Ifd35529b44c957737bf422127283c08e['h00b7a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005be] =  Ifd35529b44c957737bf422127283c08e['h00b7c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005bf] =  Ifd35529b44c957737bf422127283c08e['h00b7e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005c0] =  Ifd35529b44c957737bf422127283c08e['h00b80] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005c1] =  Ifd35529b44c957737bf422127283c08e['h00b82] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005c2] =  Ifd35529b44c957737bf422127283c08e['h00b84] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005c3] =  Ifd35529b44c957737bf422127283c08e['h00b86] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005c4] =  Ifd35529b44c957737bf422127283c08e['h00b88] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005c5] =  Ifd35529b44c957737bf422127283c08e['h00b8a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005c6] =  Ifd35529b44c957737bf422127283c08e['h00b8c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005c7] =  Ifd35529b44c957737bf422127283c08e['h00b8e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005c8] =  Ifd35529b44c957737bf422127283c08e['h00b90] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005c9] =  Ifd35529b44c957737bf422127283c08e['h00b92] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005ca] =  Ifd35529b44c957737bf422127283c08e['h00b94] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005cb] =  Ifd35529b44c957737bf422127283c08e['h00b96] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005cc] =  Ifd35529b44c957737bf422127283c08e['h00b98] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005cd] =  Ifd35529b44c957737bf422127283c08e['h00b9a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005ce] =  Ifd35529b44c957737bf422127283c08e['h00b9c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005cf] =  Ifd35529b44c957737bf422127283c08e['h00b9e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005d0] =  Ifd35529b44c957737bf422127283c08e['h00ba0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005d1] =  Ifd35529b44c957737bf422127283c08e['h00ba2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005d2] =  Ifd35529b44c957737bf422127283c08e['h00ba4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005d3] =  Ifd35529b44c957737bf422127283c08e['h00ba6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005d4] =  Ifd35529b44c957737bf422127283c08e['h00ba8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005d5] =  Ifd35529b44c957737bf422127283c08e['h00baa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005d6] =  Ifd35529b44c957737bf422127283c08e['h00bac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005d7] =  Ifd35529b44c957737bf422127283c08e['h00bae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005d8] =  Ifd35529b44c957737bf422127283c08e['h00bb0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005d9] =  Ifd35529b44c957737bf422127283c08e['h00bb2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005da] =  Ifd35529b44c957737bf422127283c08e['h00bb4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005db] =  Ifd35529b44c957737bf422127283c08e['h00bb6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005dc] =  Ifd35529b44c957737bf422127283c08e['h00bb8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005dd] =  Ifd35529b44c957737bf422127283c08e['h00bba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005de] =  Ifd35529b44c957737bf422127283c08e['h00bbc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005df] =  Ifd35529b44c957737bf422127283c08e['h00bbe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005e0] =  Ifd35529b44c957737bf422127283c08e['h00bc0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005e1] =  Ifd35529b44c957737bf422127283c08e['h00bc2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005e2] =  Ifd35529b44c957737bf422127283c08e['h00bc4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005e3] =  Ifd35529b44c957737bf422127283c08e['h00bc6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005e4] =  Ifd35529b44c957737bf422127283c08e['h00bc8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005e5] =  Ifd35529b44c957737bf422127283c08e['h00bca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005e6] =  Ifd35529b44c957737bf422127283c08e['h00bcc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005e7] =  Ifd35529b44c957737bf422127283c08e['h00bce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005e8] =  Ifd35529b44c957737bf422127283c08e['h00bd0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005e9] =  Ifd35529b44c957737bf422127283c08e['h00bd2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005ea] =  Ifd35529b44c957737bf422127283c08e['h00bd4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005eb] =  Ifd35529b44c957737bf422127283c08e['h00bd6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005ec] =  Ifd35529b44c957737bf422127283c08e['h00bd8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005ed] =  Ifd35529b44c957737bf422127283c08e['h00bda] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005ee] =  Ifd35529b44c957737bf422127283c08e['h00bdc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005ef] =  Ifd35529b44c957737bf422127283c08e['h00bde] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005f0] =  Ifd35529b44c957737bf422127283c08e['h00be0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005f1] =  Ifd35529b44c957737bf422127283c08e['h00be2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005f2] =  Ifd35529b44c957737bf422127283c08e['h00be4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005f3] =  Ifd35529b44c957737bf422127283c08e['h00be6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005f4] =  Ifd35529b44c957737bf422127283c08e['h00be8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005f5] =  Ifd35529b44c957737bf422127283c08e['h00bea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005f6] =  Ifd35529b44c957737bf422127283c08e['h00bec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005f7] =  Ifd35529b44c957737bf422127283c08e['h00bee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005f8] =  Ifd35529b44c957737bf422127283c08e['h00bf0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005f9] =  Ifd35529b44c957737bf422127283c08e['h00bf2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005fa] =  Ifd35529b44c957737bf422127283c08e['h00bf4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005fb] =  Ifd35529b44c957737bf422127283c08e['h00bf6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005fc] =  Ifd35529b44c957737bf422127283c08e['h00bf8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005fd] =  Ifd35529b44c957737bf422127283c08e['h00bfa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005fe] =  Ifd35529b44c957737bf422127283c08e['h00bfc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h005ff] =  Ifd35529b44c957737bf422127283c08e['h00bfe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00600] =  Ifd35529b44c957737bf422127283c08e['h00c00] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00601] =  Ifd35529b44c957737bf422127283c08e['h00c02] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00602] =  Ifd35529b44c957737bf422127283c08e['h00c04] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00603] =  Ifd35529b44c957737bf422127283c08e['h00c06] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00604] =  Ifd35529b44c957737bf422127283c08e['h00c08] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00605] =  Ifd35529b44c957737bf422127283c08e['h00c0a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00606] =  Ifd35529b44c957737bf422127283c08e['h00c0c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00607] =  Ifd35529b44c957737bf422127283c08e['h00c0e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00608] =  Ifd35529b44c957737bf422127283c08e['h00c10] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00609] =  Ifd35529b44c957737bf422127283c08e['h00c12] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0060a] =  Ifd35529b44c957737bf422127283c08e['h00c14] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0060b] =  Ifd35529b44c957737bf422127283c08e['h00c16] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0060c] =  Ifd35529b44c957737bf422127283c08e['h00c18] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0060d] =  Ifd35529b44c957737bf422127283c08e['h00c1a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0060e] =  Ifd35529b44c957737bf422127283c08e['h00c1c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0060f] =  Ifd35529b44c957737bf422127283c08e['h00c1e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00610] =  Ifd35529b44c957737bf422127283c08e['h00c20] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00611] =  Ifd35529b44c957737bf422127283c08e['h00c22] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00612] =  Ifd35529b44c957737bf422127283c08e['h00c24] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00613] =  Ifd35529b44c957737bf422127283c08e['h00c26] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00614] =  Ifd35529b44c957737bf422127283c08e['h00c28] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00615] =  Ifd35529b44c957737bf422127283c08e['h00c2a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00616] =  Ifd35529b44c957737bf422127283c08e['h00c2c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00617] =  Ifd35529b44c957737bf422127283c08e['h00c2e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00618] =  Ifd35529b44c957737bf422127283c08e['h00c30] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00619] =  Ifd35529b44c957737bf422127283c08e['h00c32] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0061a] =  Ifd35529b44c957737bf422127283c08e['h00c34] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0061b] =  Ifd35529b44c957737bf422127283c08e['h00c36] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0061c] =  Ifd35529b44c957737bf422127283c08e['h00c38] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0061d] =  Ifd35529b44c957737bf422127283c08e['h00c3a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0061e] =  Ifd35529b44c957737bf422127283c08e['h00c3c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0061f] =  Ifd35529b44c957737bf422127283c08e['h00c3e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00620] =  Ifd35529b44c957737bf422127283c08e['h00c40] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00621] =  Ifd35529b44c957737bf422127283c08e['h00c42] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00622] =  Ifd35529b44c957737bf422127283c08e['h00c44] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00623] =  Ifd35529b44c957737bf422127283c08e['h00c46] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00624] =  Ifd35529b44c957737bf422127283c08e['h00c48] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00625] =  Ifd35529b44c957737bf422127283c08e['h00c4a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00626] =  Ifd35529b44c957737bf422127283c08e['h00c4c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00627] =  Ifd35529b44c957737bf422127283c08e['h00c4e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00628] =  Ifd35529b44c957737bf422127283c08e['h00c50] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00629] =  Ifd35529b44c957737bf422127283c08e['h00c52] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0062a] =  Ifd35529b44c957737bf422127283c08e['h00c54] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0062b] =  Ifd35529b44c957737bf422127283c08e['h00c56] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0062c] =  Ifd35529b44c957737bf422127283c08e['h00c58] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0062d] =  Ifd35529b44c957737bf422127283c08e['h00c5a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0062e] =  Ifd35529b44c957737bf422127283c08e['h00c5c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0062f] =  Ifd35529b44c957737bf422127283c08e['h00c5e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00630] =  Ifd35529b44c957737bf422127283c08e['h00c60] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00631] =  Ifd35529b44c957737bf422127283c08e['h00c62] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00632] =  Ifd35529b44c957737bf422127283c08e['h00c64] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00633] =  Ifd35529b44c957737bf422127283c08e['h00c66] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00634] =  Ifd35529b44c957737bf422127283c08e['h00c68] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00635] =  Ifd35529b44c957737bf422127283c08e['h00c6a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00636] =  Ifd35529b44c957737bf422127283c08e['h00c6c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00637] =  Ifd35529b44c957737bf422127283c08e['h00c6e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00638] =  Ifd35529b44c957737bf422127283c08e['h00c70] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00639] =  Ifd35529b44c957737bf422127283c08e['h00c72] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0063a] =  Ifd35529b44c957737bf422127283c08e['h00c74] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0063b] =  Ifd35529b44c957737bf422127283c08e['h00c76] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0063c] =  Ifd35529b44c957737bf422127283c08e['h00c78] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0063d] =  Ifd35529b44c957737bf422127283c08e['h00c7a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0063e] =  Ifd35529b44c957737bf422127283c08e['h00c7c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0063f] =  Ifd35529b44c957737bf422127283c08e['h00c7e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00640] =  Ifd35529b44c957737bf422127283c08e['h00c80] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00641] =  Ifd35529b44c957737bf422127283c08e['h00c82] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00642] =  Ifd35529b44c957737bf422127283c08e['h00c84] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00643] =  Ifd35529b44c957737bf422127283c08e['h00c86] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00644] =  Ifd35529b44c957737bf422127283c08e['h00c88] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00645] =  Ifd35529b44c957737bf422127283c08e['h00c8a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00646] =  Ifd35529b44c957737bf422127283c08e['h00c8c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00647] =  Ifd35529b44c957737bf422127283c08e['h00c8e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00648] =  Ifd35529b44c957737bf422127283c08e['h00c90] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00649] =  Ifd35529b44c957737bf422127283c08e['h00c92] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0064a] =  Ifd35529b44c957737bf422127283c08e['h00c94] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0064b] =  Ifd35529b44c957737bf422127283c08e['h00c96] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0064c] =  Ifd35529b44c957737bf422127283c08e['h00c98] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0064d] =  Ifd35529b44c957737bf422127283c08e['h00c9a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0064e] =  Ifd35529b44c957737bf422127283c08e['h00c9c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0064f] =  Ifd35529b44c957737bf422127283c08e['h00c9e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00650] =  Ifd35529b44c957737bf422127283c08e['h00ca0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00651] =  Ifd35529b44c957737bf422127283c08e['h00ca2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00652] =  Ifd35529b44c957737bf422127283c08e['h00ca4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00653] =  Ifd35529b44c957737bf422127283c08e['h00ca6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00654] =  Ifd35529b44c957737bf422127283c08e['h00ca8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00655] =  Ifd35529b44c957737bf422127283c08e['h00caa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00656] =  Ifd35529b44c957737bf422127283c08e['h00cac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00657] =  Ifd35529b44c957737bf422127283c08e['h00cae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00658] =  Ifd35529b44c957737bf422127283c08e['h00cb0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00659] =  Ifd35529b44c957737bf422127283c08e['h00cb2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0065a] =  Ifd35529b44c957737bf422127283c08e['h00cb4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0065b] =  Ifd35529b44c957737bf422127283c08e['h00cb6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0065c] =  Ifd35529b44c957737bf422127283c08e['h00cb8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0065d] =  Ifd35529b44c957737bf422127283c08e['h00cba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0065e] =  Ifd35529b44c957737bf422127283c08e['h00cbc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0065f] =  Ifd35529b44c957737bf422127283c08e['h00cbe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00660] =  Ifd35529b44c957737bf422127283c08e['h00cc0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00661] =  Ifd35529b44c957737bf422127283c08e['h00cc2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00662] =  Ifd35529b44c957737bf422127283c08e['h00cc4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00663] =  Ifd35529b44c957737bf422127283c08e['h00cc6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00664] =  Ifd35529b44c957737bf422127283c08e['h00cc8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00665] =  Ifd35529b44c957737bf422127283c08e['h00cca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00666] =  Ifd35529b44c957737bf422127283c08e['h00ccc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00667] =  Ifd35529b44c957737bf422127283c08e['h00cce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00668] =  Ifd35529b44c957737bf422127283c08e['h00cd0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00669] =  Ifd35529b44c957737bf422127283c08e['h00cd2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0066a] =  Ifd35529b44c957737bf422127283c08e['h00cd4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0066b] =  Ifd35529b44c957737bf422127283c08e['h00cd6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0066c] =  Ifd35529b44c957737bf422127283c08e['h00cd8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0066d] =  Ifd35529b44c957737bf422127283c08e['h00cda] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0066e] =  Ifd35529b44c957737bf422127283c08e['h00cdc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0066f] =  Ifd35529b44c957737bf422127283c08e['h00cde] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00670] =  Ifd35529b44c957737bf422127283c08e['h00ce0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00671] =  Ifd35529b44c957737bf422127283c08e['h00ce2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00672] =  Ifd35529b44c957737bf422127283c08e['h00ce4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00673] =  Ifd35529b44c957737bf422127283c08e['h00ce6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00674] =  Ifd35529b44c957737bf422127283c08e['h00ce8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00675] =  Ifd35529b44c957737bf422127283c08e['h00cea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00676] =  Ifd35529b44c957737bf422127283c08e['h00cec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00677] =  Ifd35529b44c957737bf422127283c08e['h00cee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00678] =  Ifd35529b44c957737bf422127283c08e['h00cf0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00679] =  Ifd35529b44c957737bf422127283c08e['h00cf2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0067a] =  Ifd35529b44c957737bf422127283c08e['h00cf4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0067b] =  Ifd35529b44c957737bf422127283c08e['h00cf6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0067c] =  Ifd35529b44c957737bf422127283c08e['h00cf8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0067d] =  Ifd35529b44c957737bf422127283c08e['h00cfa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0067e] =  Ifd35529b44c957737bf422127283c08e['h00cfc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0067f] =  Ifd35529b44c957737bf422127283c08e['h00cfe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00680] =  Ifd35529b44c957737bf422127283c08e['h00d00] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00681] =  Ifd35529b44c957737bf422127283c08e['h00d02] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00682] =  Ifd35529b44c957737bf422127283c08e['h00d04] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00683] =  Ifd35529b44c957737bf422127283c08e['h00d06] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00684] =  Ifd35529b44c957737bf422127283c08e['h00d08] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00685] =  Ifd35529b44c957737bf422127283c08e['h00d0a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00686] =  Ifd35529b44c957737bf422127283c08e['h00d0c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00687] =  Ifd35529b44c957737bf422127283c08e['h00d0e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00688] =  Ifd35529b44c957737bf422127283c08e['h00d10] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00689] =  Ifd35529b44c957737bf422127283c08e['h00d12] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0068a] =  Ifd35529b44c957737bf422127283c08e['h00d14] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0068b] =  Ifd35529b44c957737bf422127283c08e['h00d16] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0068c] =  Ifd35529b44c957737bf422127283c08e['h00d18] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0068d] =  Ifd35529b44c957737bf422127283c08e['h00d1a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0068e] =  Ifd35529b44c957737bf422127283c08e['h00d1c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0068f] =  Ifd35529b44c957737bf422127283c08e['h00d1e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00690] =  Ifd35529b44c957737bf422127283c08e['h00d20] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00691] =  Ifd35529b44c957737bf422127283c08e['h00d22] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00692] =  Ifd35529b44c957737bf422127283c08e['h00d24] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00693] =  Ifd35529b44c957737bf422127283c08e['h00d26] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00694] =  Ifd35529b44c957737bf422127283c08e['h00d28] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00695] =  Ifd35529b44c957737bf422127283c08e['h00d2a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00696] =  Ifd35529b44c957737bf422127283c08e['h00d2c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00697] =  Ifd35529b44c957737bf422127283c08e['h00d2e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00698] =  Ifd35529b44c957737bf422127283c08e['h00d30] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00699] =  Ifd35529b44c957737bf422127283c08e['h00d32] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0069a] =  Ifd35529b44c957737bf422127283c08e['h00d34] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0069b] =  Ifd35529b44c957737bf422127283c08e['h00d36] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0069c] =  Ifd35529b44c957737bf422127283c08e['h00d38] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0069d] =  Ifd35529b44c957737bf422127283c08e['h00d3a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0069e] =  Ifd35529b44c957737bf422127283c08e['h00d3c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0069f] =  Ifd35529b44c957737bf422127283c08e['h00d3e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006a0] =  Ifd35529b44c957737bf422127283c08e['h00d40] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006a1] =  Ifd35529b44c957737bf422127283c08e['h00d42] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006a2] =  Ifd35529b44c957737bf422127283c08e['h00d44] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006a3] =  Ifd35529b44c957737bf422127283c08e['h00d46] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006a4] =  Ifd35529b44c957737bf422127283c08e['h00d48] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006a5] =  Ifd35529b44c957737bf422127283c08e['h00d4a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006a6] =  Ifd35529b44c957737bf422127283c08e['h00d4c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006a7] =  Ifd35529b44c957737bf422127283c08e['h00d4e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006a8] =  Ifd35529b44c957737bf422127283c08e['h00d50] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006a9] =  Ifd35529b44c957737bf422127283c08e['h00d52] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006aa] =  Ifd35529b44c957737bf422127283c08e['h00d54] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006ab] =  Ifd35529b44c957737bf422127283c08e['h00d56] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006ac] =  Ifd35529b44c957737bf422127283c08e['h00d58] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006ad] =  Ifd35529b44c957737bf422127283c08e['h00d5a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006ae] =  Ifd35529b44c957737bf422127283c08e['h00d5c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006af] =  Ifd35529b44c957737bf422127283c08e['h00d5e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006b0] =  Ifd35529b44c957737bf422127283c08e['h00d60] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006b1] =  Ifd35529b44c957737bf422127283c08e['h00d62] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006b2] =  Ifd35529b44c957737bf422127283c08e['h00d64] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006b3] =  Ifd35529b44c957737bf422127283c08e['h00d66] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006b4] =  Ifd35529b44c957737bf422127283c08e['h00d68] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006b5] =  Ifd35529b44c957737bf422127283c08e['h00d6a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006b6] =  Ifd35529b44c957737bf422127283c08e['h00d6c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006b7] =  Ifd35529b44c957737bf422127283c08e['h00d6e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006b8] =  Ifd35529b44c957737bf422127283c08e['h00d70] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006b9] =  Ifd35529b44c957737bf422127283c08e['h00d72] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006ba] =  Ifd35529b44c957737bf422127283c08e['h00d74] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006bb] =  Ifd35529b44c957737bf422127283c08e['h00d76] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006bc] =  Ifd35529b44c957737bf422127283c08e['h00d78] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006bd] =  Ifd35529b44c957737bf422127283c08e['h00d7a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006be] =  Ifd35529b44c957737bf422127283c08e['h00d7c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006bf] =  Ifd35529b44c957737bf422127283c08e['h00d7e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006c0] =  Ifd35529b44c957737bf422127283c08e['h00d80] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006c1] =  Ifd35529b44c957737bf422127283c08e['h00d82] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006c2] =  Ifd35529b44c957737bf422127283c08e['h00d84] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006c3] =  Ifd35529b44c957737bf422127283c08e['h00d86] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006c4] =  Ifd35529b44c957737bf422127283c08e['h00d88] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006c5] =  Ifd35529b44c957737bf422127283c08e['h00d8a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006c6] =  Ifd35529b44c957737bf422127283c08e['h00d8c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006c7] =  Ifd35529b44c957737bf422127283c08e['h00d8e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006c8] =  Ifd35529b44c957737bf422127283c08e['h00d90] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006c9] =  Ifd35529b44c957737bf422127283c08e['h00d92] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006ca] =  Ifd35529b44c957737bf422127283c08e['h00d94] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006cb] =  Ifd35529b44c957737bf422127283c08e['h00d96] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006cc] =  Ifd35529b44c957737bf422127283c08e['h00d98] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006cd] =  Ifd35529b44c957737bf422127283c08e['h00d9a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006ce] =  Ifd35529b44c957737bf422127283c08e['h00d9c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006cf] =  Ifd35529b44c957737bf422127283c08e['h00d9e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006d0] =  Ifd35529b44c957737bf422127283c08e['h00da0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006d1] =  Ifd35529b44c957737bf422127283c08e['h00da2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006d2] =  Ifd35529b44c957737bf422127283c08e['h00da4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006d3] =  Ifd35529b44c957737bf422127283c08e['h00da6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006d4] =  Ifd35529b44c957737bf422127283c08e['h00da8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006d5] =  Ifd35529b44c957737bf422127283c08e['h00daa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006d6] =  Ifd35529b44c957737bf422127283c08e['h00dac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006d7] =  Ifd35529b44c957737bf422127283c08e['h00dae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006d8] =  Ifd35529b44c957737bf422127283c08e['h00db0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006d9] =  Ifd35529b44c957737bf422127283c08e['h00db2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006da] =  Ifd35529b44c957737bf422127283c08e['h00db4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006db] =  Ifd35529b44c957737bf422127283c08e['h00db6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006dc] =  Ifd35529b44c957737bf422127283c08e['h00db8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006dd] =  Ifd35529b44c957737bf422127283c08e['h00dba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006de] =  Ifd35529b44c957737bf422127283c08e['h00dbc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006df] =  Ifd35529b44c957737bf422127283c08e['h00dbe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006e0] =  Ifd35529b44c957737bf422127283c08e['h00dc0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006e1] =  Ifd35529b44c957737bf422127283c08e['h00dc2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006e2] =  Ifd35529b44c957737bf422127283c08e['h00dc4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006e3] =  Ifd35529b44c957737bf422127283c08e['h00dc6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006e4] =  Ifd35529b44c957737bf422127283c08e['h00dc8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006e5] =  Ifd35529b44c957737bf422127283c08e['h00dca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006e6] =  Ifd35529b44c957737bf422127283c08e['h00dcc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006e7] =  Ifd35529b44c957737bf422127283c08e['h00dce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006e8] =  Ifd35529b44c957737bf422127283c08e['h00dd0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006e9] =  Ifd35529b44c957737bf422127283c08e['h00dd2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006ea] =  Ifd35529b44c957737bf422127283c08e['h00dd4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006eb] =  Ifd35529b44c957737bf422127283c08e['h00dd6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006ec] =  Ifd35529b44c957737bf422127283c08e['h00dd8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006ed] =  Ifd35529b44c957737bf422127283c08e['h00dda] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006ee] =  Ifd35529b44c957737bf422127283c08e['h00ddc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006ef] =  Ifd35529b44c957737bf422127283c08e['h00dde] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006f0] =  Ifd35529b44c957737bf422127283c08e['h00de0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006f1] =  Ifd35529b44c957737bf422127283c08e['h00de2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006f2] =  Ifd35529b44c957737bf422127283c08e['h00de4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006f3] =  Ifd35529b44c957737bf422127283c08e['h00de6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006f4] =  Ifd35529b44c957737bf422127283c08e['h00de8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006f5] =  Ifd35529b44c957737bf422127283c08e['h00dea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006f6] =  Ifd35529b44c957737bf422127283c08e['h00dec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006f7] =  Ifd35529b44c957737bf422127283c08e['h00dee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006f8] =  Ifd35529b44c957737bf422127283c08e['h00df0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006f9] =  Ifd35529b44c957737bf422127283c08e['h00df2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006fa] =  Ifd35529b44c957737bf422127283c08e['h00df4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006fb] =  Ifd35529b44c957737bf422127283c08e['h00df6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006fc] =  Ifd35529b44c957737bf422127283c08e['h00df8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006fd] =  Ifd35529b44c957737bf422127283c08e['h00dfa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006fe] =  Ifd35529b44c957737bf422127283c08e['h00dfc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h006ff] =  Ifd35529b44c957737bf422127283c08e['h00dfe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00700] =  Ifd35529b44c957737bf422127283c08e['h00e00] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00701] =  Ifd35529b44c957737bf422127283c08e['h00e02] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00702] =  Ifd35529b44c957737bf422127283c08e['h00e04] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00703] =  Ifd35529b44c957737bf422127283c08e['h00e06] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00704] =  Ifd35529b44c957737bf422127283c08e['h00e08] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00705] =  Ifd35529b44c957737bf422127283c08e['h00e0a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00706] =  Ifd35529b44c957737bf422127283c08e['h00e0c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00707] =  Ifd35529b44c957737bf422127283c08e['h00e0e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00708] =  Ifd35529b44c957737bf422127283c08e['h00e10] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00709] =  Ifd35529b44c957737bf422127283c08e['h00e12] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0070a] =  Ifd35529b44c957737bf422127283c08e['h00e14] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0070b] =  Ifd35529b44c957737bf422127283c08e['h00e16] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0070c] =  Ifd35529b44c957737bf422127283c08e['h00e18] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0070d] =  Ifd35529b44c957737bf422127283c08e['h00e1a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0070e] =  Ifd35529b44c957737bf422127283c08e['h00e1c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0070f] =  Ifd35529b44c957737bf422127283c08e['h00e1e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00710] =  Ifd35529b44c957737bf422127283c08e['h00e20] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00711] =  Ifd35529b44c957737bf422127283c08e['h00e22] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00712] =  Ifd35529b44c957737bf422127283c08e['h00e24] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00713] =  Ifd35529b44c957737bf422127283c08e['h00e26] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00714] =  Ifd35529b44c957737bf422127283c08e['h00e28] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00715] =  Ifd35529b44c957737bf422127283c08e['h00e2a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00716] =  Ifd35529b44c957737bf422127283c08e['h00e2c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00717] =  Ifd35529b44c957737bf422127283c08e['h00e2e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00718] =  Ifd35529b44c957737bf422127283c08e['h00e30] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00719] =  Ifd35529b44c957737bf422127283c08e['h00e32] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0071a] =  Ifd35529b44c957737bf422127283c08e['h00e34] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0071b] =  Ifd35529b44c957737bf422127283c08e['h00e36] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0071c] =  Ifd35529b44c957737bf422127283c08e['h00e38] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0071d] =  Ifd35529b44c957737bf422127283c08e['h00e3a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0071e] =  Ifd35529b44c957737bf422127283c08e['h00e3c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0071f] =  Ifd35529b44c957737bf422127283c08e['h00e3e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00720] =  Ifd35529b44c957737bf422127283c08e['h00e40] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00721] =  Ifd35529b44c957737bf422127283c08e['h00e42] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00722] =  Ifd35529b44c957737bf422127283c08e['h00e44] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00723] =  Ifd35529b44c957737bf422127283c08e['h00e46] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00724] =  Ifd35529b44c957737bf422127283c08e['h00e48] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00725] =  Ifd35529b44c957737bf422127283c08e['h00e4a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00726] =  Ifd35529b44c957737bf422127283c08e['h00e4c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00727] =  Ifd35529b44c957737bf422127283c08e['h00e4e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00728] =  Ifd35529b44c957737bf422127283c08e['h00e50] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00729] =  Ifd35529b44c957737bf422127283c08e['h00e52] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0072a] =  Ifd35529b44c957737bf422127283c08e['h00e54] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0072b] =  Ifd35529b44c957737bf422127283c08e['h00e56] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0072c] =  Ifd35529b44c957737bf422127283c08e['h00e58] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0072d] =  Ifd35529b44c957737bf422127283c08e['h00e5a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0072e] =  Ifd35529b44c957737bf422127283c08e['h00e5c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0072f] =  Ifd35529b44c957737bf422127283c08e['h00e5e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00730] =  Ifd35529b44c957737bf422127283c08e['h00e60] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00731] =  Ifd35529b44c957737bf422127283c08e['h00e62] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00732] =  Ifd35529b44c957737bf422127283c08e['h00e64] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00733] =  Ifd35529b44c957737bf422127283c08e['h00e66] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00734] =  Ifd35529b44c957737bf422127283c08e['h00e68] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00735] =  Ifd35529b44c957737bf422127283c08e['h00e6a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00736] =  Ifd35529b44c957737bf422127283c08e['h00e6c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00737] =  Ifd35529b44c957737bf422127283c08e['h00e6e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00738] =  Ifd35529b44c957737bf422127283c08e['h00e70] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00739] =  Ifd35529b44c957737bf422127283c08e['h00e72] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0073a] =  Ifd35529b44c957737bf422127283c08e['h00e74] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0073b] =  Ifd35529b44c957737bf422127283c08e['h00e76] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0073c] =  Ifd35529b44c957737bf422127283c08e['h00e78] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0073d] =  Ifd35529b44c957737bf422127283c08e['h00e7a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0073e] =  Ifd35529b44c957737bf422127283c08e['h00e7c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0073f] =  Ifd35529b44c957737bf422127283c08e['h00e7e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00740] =  Ifd35529b44c957737bf422127283c08e['h00e80] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00741] =  Ifd35529b44c957737bf422127283c08e['h00e82] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00742] =  Ifd35529b44c957737bf422127283c08e['h00e84] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00743] =  Ifd35529b44c957737bf422127283c08e['h00e86] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00744] =  Ifd35529b44c957737bf422127283c08e['h00e88] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00745] =  Ifd35529b44c957737bf422127283c08e['h00e8a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00746] =  Ifd35529b44c957737bf422127283c08e['h00e8c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00747] =  Ifd35529b44c957737bf422127283c08e['h00e8e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00748] =  Ifd35529b44c957737bf422127283c08e['h00e90] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00749] =  Ifd35529b44c957737bf422127283c08e['h00e92] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0074a] =  Ifd35529b44c957737bf422127283c08e['h00e94] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0074b] =  Ifd35529b44c957737bf422127283c08e['h00e96] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0074c] =  Ifd35529b44c957737bf422127283c08e['h00e98] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0074d] =  Ifd35529b44c957737bf422127283c08e['h00e9a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0074e] =  Ifd35529b44c957737bf422127283c08e['h00e9c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0074f] =  Ifd35529b44c957737bf422127283c08e['h00e9e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00750] =  Ifd35529b44c957737bf422127283c08e['h00ea0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00751] =  Ifd35529b44c957737bf422127283c08e['h00ea2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00752] =  Ifd35529b44c957737bf422127283c08e['h00ea4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00753] =  Ifd35529b44c957737bf422127283c08e['h00ea6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00754] =  Ifd35529b44c957737bf422127283c08e['h00ea8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00755] =  Ifd35529b44c957737bf422127283c08e['h00eaa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00756] =  Ifd35529b44c957737bf422127283c08e['h00eac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00757] =  Ifd35529b44c957737bf422127283c08e['h00eae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00758] =  Ifd35529b44c957737bf422127283c08e['h00eb0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00759] =  Ifd35529b44c957737bf422127283c08e['h00eb2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0075a] =  Ifd35529b44c957737bf422127283c08e['h00eb4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0075b] =  Ifd35529b44c957737bf422127283c08e['h00eb6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0075c] =  Ifd35529b44c957737bf422127283c08e['h00eb8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0075d] =  Ifd35529b44c957737bf422127283c08e['h00eba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0075e] =  Ifd35529b44c957737bf422127283c08e['h00ebc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0075f] =  Ifd35529b44c957737bf422127283c08e['h00ebe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00760] =  Ifd35529b44c957737bf422127283c08e['h00ec0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00761] =  Ifd35529b44c957737bf422127283c08e['h00ec2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00762] =  Ifd35529b44c957737bf422127283c08e['h00ec4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00763] =  Ifd35529b44c957737bf422127283c08e['h00ec6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00764] =  Ifd35529b44c957737bf422127283c08e['h00ec8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00765] =  Ifd35529b44c957737bf422127283c08e['h00eca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00766] =  Ifd35529b44c957737bf422127283c08e['h00ecc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00767] =  Ifd35529b44c957737bf422127283c08e['h00ece] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00768] =  Ifd35529b44c957737bf422127283c08e['h00ed0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00769] =  Ifd35529b44c957737bf422127283c08e['h00ed2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0076a] =  Ifd35529b44c957737bf422127283c08e['h00ed4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0076b] =  Ifd35529b44c957737bf422127283c08e['h00ed6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0076c] =  Ifd35529b44c957737bf422127283c08e['h00ed8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0076d] =  Ifd35529b44c957737bf422127283c08e['h00eda] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0076e] =  Ifd35529b44c957737bf422127283c08e['h00edc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0076f] =  Ifd35529b44c957737bf422127283c08e['h00ede] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00770] =  Ifd35529b44c957737bf422127283c08e['h00ee0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00771] =  Ifd35529b44c957737bf422127283c08e['h00ee2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00772] =  Ifd35529b44c957737bf422127283c08e['h00ee4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00773] =  Ifd35529b44c957737bf422127283c08e['h00ee6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00774] =  Ifd35529b44c957737bf422127283c08e['h00ee8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00775] =  Ifd35529b44c957737bf422127283c08e['h00eea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00776] =  Ifd35529b44c957737bf422127283c08e['h00eec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00777] =  Ifd35529b44c957737bf422127283c08e['h00eee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00778] =  Ifd35529b44c957737bf422127283c08e['h00ef0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00779] =  Ifd35529b44c957737bf422127283c08e['h00ef2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0077a] =  Ifd35529b44c957737bf422127283c08e['h00ef4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0077b] =  Ifd35529b44c957737bf422127283c08e['h00ef6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0077c] =  Ifd35529b44c957737bf422127283c08e['h00ef8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0077d] =  Ifd35529b44c957737bf422127283c08e['h00efa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0077e] =  Ifd35529b44c957737bf422127283c08e['h00efc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0077f] =  Ifd35529b44c957737bf422127283c08e['h00efe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00780] =  Ifd35529b44c957737bf422127283c08e['h00f00] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00781] =  Ifd35529b44c957737bf422127283c08e['h00f02] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00782] =  Ifd35529b44c957737bf422127283c08e['h00f04] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00783] =  Ifd35529b44c957737bf422127283c08e['h00f06] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00784] =  Ifd35529b44c957737bf422127283c08e['h00f08] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00785] =  Ifd35529b44c957737bf422127283c08e['h00f0a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00786] =  Ifd35529b44c957737bf422127283c08e['h00f0c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00787] =  Ifd35529b44c957737bf422127283c08e['h00f0e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00788] =  Ifd35529b44c957737bf422127283c08e['h00f10] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00789] =  Ifd35529b44c957737bf422127283c08e['h00f12] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0078a] =  Ifd35529b44c957737bf422127283c08e['h00f14] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0078b] =  Ifd35529b44c957737bf422127283c08e['h00f16] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0078c] =  Ifd35529b44c957737bf422127283c08e['h00f18] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0078d] =  Ifd35529b44c957737bf422127283c08e['h00f1a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0078e] =  Ifd35529b44c957737bf422127283c08e['h00f1c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0078f] =  Ifd35529b44c957737bf422127283c08e['h00f1e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00790] =  Ifd35529b44c957737bf422127283c08e['h00f20] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00791] =  Ifd35529b44c957737bf422127283c08e['h00f22] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00792] =  Ifd35529b44c957737bf422127283c08e['h00f24] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00793] =  Ifd35529b44c957737bf422127283c08e['h00f26] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00794] =  Ifd35529b44c957737bf422127283c08e['h00f28] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00795] =  Ifd35529b44c957737bf422127283c08e['h00f2a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00796] =  Ifd35529b44c957737bf422127283c08e['h00f2c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00797] =  Ifd35529b44c957737bf422127283c08e['h00f2e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00798] =  Ifd35529b44c957737bf422127283c08e['h00f30] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00799] =  Ifd35529b44c957737bf422127283c08e['h00f32] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0079a] =  Ifd35529b44c957737bf422127283c08e['h00f34] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0079b] =  Ifd35529b44c957737bf422127283c08e['h00f36] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0079c] =  Ifd35529b44c957737bf422127283c08e['h00f38] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0079d] =  Ifd35529b44c957737bf422127283c08e['h00f3a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0079e] =  Ifd35529b44c957737bf422127283c08e['h00f3c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0079f] =  Ifd35529b44c957737bf422127283c08e['h00f3e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007a0] =  Ifd35529b44c957737bf422127283c08e['h00f40] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007a1] =  Ifd35529b44c957737bf422127283c08e['h00f42] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007a2] =  Ifd35529b44c957737bf422127283c08e['h00f44] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007a3] =  Ifd35529b44c957737bf422127283c08e['h00f46] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007a4] =  Ifd35529b44c957737bf422127283c08e['h00f48] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007a5] =  Ifd35529b44c957737bf422127283c08e['h00f4a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007a6] =  Ifd35529b44c957737bf422127283c08e['h00f4c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007a7] =  Ifd35529b44c957737bf422127283c08e['h00f4e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007a8] =  Ifd35529b44c957737bf422127283c08e['h00f50] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007a9] =  Ifd35529b44c957737bf422127283c08e['h00f52] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007aa] =  Ifd35529b44c957737bf422127283c08e['h00f54] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007ab] =  Ifd35529b44c957737bf422127283c08e['h00f56] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007ac] =  Ifd35529b44c957737bf422127283c08e['h00f58] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007ad] =  Ifd35529b44c957737bf422127283c08e['h00f5a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007ae] =  Ifd35529b44c957737bf422127283c08e['h00f5c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007af] =  Ifd35529b44c957737bf422127283c08e['h00f5e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007b0] =  Ifd35529b44c957737bf422127283c08e['h00f60] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007b1] =  Ifd35529b44c957737bf422127283c08e['h00f62] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007b2] =  Ifd35529b44c957737bf422127283c08e['h00f64] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007b3] =  Ifd35529b44c957737bf422127283c08e['h00f66] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007b4] =  Ifd35529b44c957737bf422127283c08e['h00f68] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007b5] =  Ifd35529b44c957737bf422127283c08e['h00f6a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007b6] =  Ifd35529b44c957737bf422127283c08e['h00f6c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007b7] =  Ifd35529b44c957737bf422127283c08e['h00f6e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007b8] =  Ifd35529b44c957737bf422127283c08e['h00f70] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007b9] =  Ifd35529b44c957737bf422127283c08e['h00f72] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007ba] =  Ifd35529b44c957737bf422127283c08e['h00f74] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007bb] =  Ifd35529b44c957737bf422127283c08e['h00f76] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007bc] =  Ifd35529b44c957737bf422127283c08e['h00f78] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007bd] =  Ifd35529b44c957737bf422127283c08e['h00f7a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007be] =  Ifd35529b44c957737bf422127283c08e['h00f7c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007bf] =  Ifd35529b44c957737bf422127283c08e['h00f7e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007c0] =  Ifd35529b44c957737bf422127283c08e['h00f80] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007c1] =  Ifd35529b44c957737bf422127283c08e['h00f82] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007c2] =  Ifd35529b44c957737bf422127283c08e['h00f84] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007c3] =  Ifd35529b44c957737bf422127283c08e['h00f86] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007c4] =  Ifd35529b44c957737bf422127283c08e['h00f88] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007c5] =  Ifd35529b44c957737bf422127283c08e['h00f8a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007c6] =  Ifd35529b44c957737bf422127283c08e['h00f8c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007c7] =  Ifd35529b44c957737bf422127283c08e['h00f8e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007c8] =  Ifd35529b44c957737bf422127283c08e['h00f90] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007c9] =  Ifd35529b44c957737bf422127283c08e['h00f92] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007ca] =  Ifd35529b44c957737bf422127283c08e['h00f94] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007cb] =  Ifd35529b44c957737bf422127283c08e['h00f96] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007cc] =  Ifd35529b44c957737bf422127283c08e['h00f98] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007cd] =  Ifd35529b44c957737bf422127283c08e['h00f9a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007ce] =  Ifd35529b44c957737bf422127283c08e['h00f9c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007cf] =  Ifd35529b44c957737bf422127283c08e['h00f9e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007d0] =  Ifd35529b44c957737bf422127283c08e['h00fa0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007d1] =  Ifd35529b44c957737bf422127283c08e['h00fa2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007d2] =  Ifd35529b44c957737bf422127283c08e['h00fa4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007d3] =  Ifd35529b44c957737bf422127283c08e['h00fa6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007d4] =  Ifd35529b44c957737bf422127283c08e['h00fa8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007d5] =  Ifd35529b44c957737bf422127283c08e['h00faa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007d6] =  Ifd35529b44c957737bf422127283c08e['h00fac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007d7] =  Ifd35529b44c957737bf422127283c08e['h00fae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007d8] =  Ifd35529b44c957737bf422127283c08e['h00fb0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007d9] =  Ifd35529b44c957737bf422127283c08e['h00fb2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007da] =  Ifd35529b44c957737bf422127283c08e['h00fb4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007db] =  Ifd35529b44c957737bf422127283c08e['h00fb6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007dc] =  Ifd35529b44c957737bf422127283c08e['h00fb8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007dd] =  Ifd35529b44c957737bf422127283c08e['h00fba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007de] =  Ifd35529b44c957737bf422127283c08e['h00fbc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007df] =  Ifd35529b44c957737bf422127283c08e['h00fbe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007e0] =  Ifd35529b44c957737bf422127283c08e['h00fc0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007e1] =  Ifd35529b44c957737bf422127283c08e['h00fc2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007e2] =  Ifd35529b44c957737bf422127283c08e['h00fc4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007e3] =  Ifd35529b44c957737bf422127283c08e['h00fc6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007e4] =  Ifd35529b44c957737bf422127283c08e['h00fc8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007e5] =  Ifd35529b44c957737bf422127283c08e['h00fca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007e6] =  Ifd35529b44c957737bf422127283c08e['h00fcc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007e7] =  Ifd35529b44c957737bf422127283c08e['h00fce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007e8] =  Ifd35529b44c957737bf422127283c08e['h00fd0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007e9] =  Ifd35529b44c957737bf422127283c08e['h00fd2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007ea] =  Ifd35529b44c957737bf422127283c08e['h00fd4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007eb] =  Ifd35529b44c957737bf422127283c08e['h00fd6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007ec] =  Ifd35529b44c957737bf422127283c08e['h00fd8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007ed] =  Ifd35529b44c957737bf422127283c08e['h00fda] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007ee] =  Ifd35529b44c957737bf422127283c08e['h00fdc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007ef] =  Ifd35529b44c957737bf422127283c08e['h00fde] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007f0] =  Ifd35529b44c957737bf422127283c08e['h00fe0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007f1] =  Ifd35529b44c957737bf422127283c08e['h00fe2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007f2] =  Ifd35529b44c957737bf422127283c08e['h00fe4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007f3] =  Ifd35529b44c957737bf422127283c08e['h00fe6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007f4] =  Ifd35529b44c957737bf422127283c08e['h00fe8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007f5] =  Ifd35529b44c957737bf422127283c08e['h00fea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007f6] =  Ifd35529b44c957737bf422127283c08e['h00fec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007f7] =  Ifd35529b44c957737bf422127283c08e['h00fee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007f8] =  Ifd35529b44c957737bf422127283c08e['h00ff0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007f9] =  Ifd35529b44c957737bf422127283c08e['h00ff2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007fa] =  Ifd35529b44c957737bf422127283c08e['h00ff4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007fb] =  Ifd35529b44c957737bf422127283c08e['h00ff6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007fc] =  Ifd35529b44c957737bf422127283c08e['h00ff8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007fd] =  Ifd35529b44c957737bf422127283c08e['h00ffa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007fe] =  Ifd35529b44c957737bf422127283c08e['h00ffc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h007ff] =  Ifd35529b44c957737bf422127283c08e['h00ffe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00800] =  Ifd35529b44c957737bf422127283c08e['h01000] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00801] =  Ifd35529b44c957737bf422127283c08e['h01002] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00802] =  Ifd35529b44c957737bf422127283c08e['h01004] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00803] =  Ifd35529b44c957737bf422127283c08e['h01006] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00804] =  Ifd35529b44c957737bf422127283c08e['h01008] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00805] =  Ifd35529b44c957737bf422127283c08e['h0100a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00806] =  Ifd35529b44c957737bf422127283c08e['h0100c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00807] =  Ifd35529b44c957737bf422127283c08e['h0100e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00808] =  Ifd35529b44c957737bf422127283c08e['h01010] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00809] =  Ifd35529b44c957737bf422127283c08e['h01012] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0080a] =  Ifd35529b44c957737bf422127283c08e['h01014] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0080b] =  Ifd35529b44c957737bf422127283c08e['h01016] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0080c] =  Ifd35529b44c957737bf422127283c08e['h01018] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0080d] =  Ifd35529b44c957737bf422127283c08e['h0101a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0080e] =  Ifd35529b44c957737bf422127283c08e['h0101c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0080f] =  Ifd35529b44c957737bf422127283c08e['h0101e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00810] =  Ifd35529b44c957737bf422127283c08e['h01020] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00811] =  Ifd35529b44c957737bf422127283c08e['h01022] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00812] =  Ifd35529b44c957737bf422127283c08e['h01024] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00813] =  Ifd35529b44c957737bf422127283c08e['h01026] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00814] =  Ifd35529b44c957737bf422127283c08e['h01028] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00815] =  Ifd35529b44c957737bf422127283c08e['h0102a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00816] =  Ifd35529b44c957737bf422127283c08e['h0102c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00817] =  Ifd35529b44c957737bf422127283c08e['h0102e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00818] =  Ifd35529b44c957737bf422127283c08e['h01030] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00819] =  Ifd35529b44c957737bf422127283c08e['h01032] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0081a] =  Ifd35529b44c957737bf422127283c08e['h01034] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0081b] =  Ifd35529b44c957737bf422127283c08e['h01036] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0081c] =  Ifd35529b44c957737bf422127283c08e['h01038] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0081d] =  Ifd35529b44c957737bf422127283c08e['h0103a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0081e] =  Ifd35529b44c957737bf422127283c08e['h0103c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0081f] =  Ifd35529b44c957737bf422127283c08e['h0103e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00820] =  Ifd35529b44c957737bf422127283c08e['h01040] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00821] =  Ifd35529b44c957737bf422127283c08e['h01042] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00822] =  Ifd35529b44c957737bf422127283c08e['h01044] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00823] =  Ifd35529b44c957737bf422127283c08e['h01046] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00824] =  Ifd35529b44c957737bf422127283c08e['h01048] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00825] =  Ifd35529b44c957737bf422127283c08e['h0104a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00826] =  Ifd35529b44c957737bf422127283c08e['h0104c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00827] =  Ifd35529b44c957737bf422127283c08e['h0104e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00828] =  Ifd35529b44c957737bf422127283c08e['h01050] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00829] =  Ifd35529b44c957737bf422127283c08e['h01052] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0082a] =  Ifd35529b44c957737bf422127283c08e['h01054] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0082b] =  Ifd35529b44c957737bf422127283c08e['h01056] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0082c] =  Ifd35529b44c957737bf422127283c08e['h01058] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0082d] =  Ifd35529b44c957737bf422127283c08e['h0105a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0082e] =  Ifd35529b44c957737bf422127283c08e['h0105c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0082f] =  Ifd35529b44c957737bf422127283c08e['h0105e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00830] =  Ifd35529b44c957737bf422127283c08e['h01060] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00831] =  Ifd35529b44c957737bf422127283c08e['h01062] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00832] =  Ifd35529b44c957737bf422127283c08e['h01064] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00833] =  Ifd35529b44c957737bf422127283c08e['h01066] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00834] =  Ifd35529b44c957737bf422127283c08e['h01068] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00835] =  Ifd35529b44c957737bf422127283c08e['h0106a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00836] =  Ifd35529b44c957737bf422127283c08e['h0106c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00837] =  Ifd35529b44c957737bf422127283c08e['h0106e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00838] =  Ifd35529b44c957737bf422127283c08e['h01070] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00839] =  Ifd35529b44c957737bf422127283c08e['h01072] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0083a] =  Ifd35529b44c957737bf422127283c08e['h01074] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0083b] =  Ifd35529b44c957737bf422127283c08e['h01076] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0083c] =  Ifd35529b44c957737bf422127283c08e['h01078] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0083d] =  Ifd35529b44c957737bf422127283c08e['h0107a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0083e] =  Ifd35529b44c957737bf422127283c08e['h0107c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0083f] =  Ifd35529b44c957737bf422127283c08e['h0107e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00840] =  Ifd35529b44c957737bf422127283c08e['h01080] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00841] =  Ifd35529b44c957737bf422127283c08e['h01082] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00842] =  Ifd35529b44c957737bf422127283c08e['h01084] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00843] =  Ifd35529b44c957737bf422127283c08e['h01086] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00844] =  Ifd35529b44c957737bf422127283c08e['h01088] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00845] =  Ifd35529b44c957737bf422127283c08e['h0108a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00846] =  Ifd35529b44c957737bf422127283c08e['h0108c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00847] =  Ifd35529b44c957737bf422127283c08e['h0108e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00848] =  Ifd35529b44c957737bf422127283c08e['h01090] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00849] =  Ifd35529b44c957737bf422127283c08e['h01092] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0084a] =  Ifd35529b44c957737bf422127283c08e['h01094] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0084b] =  Ifd35529b44c957737bf422127283c08e['h01096] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0084c] =  Ifd35529b44c957737bf422127283c08e['h01098] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0084d] =  Ifd35529b44c957737bf422127283c08e['h0109a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0084e] =  Ifd35529b44c957737bf422127283c08e['h0109c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0084f] =  Ifd35529b44c957737bf422127283c08e['h0109e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00850] =  Ifd35529b44c957737bf422127283c08e['h010a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00851] =  Ifd35529b44c957737bf422127283c08e['h010a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00852] =  Ifd35529b44c957737bf422127283c08e['h010a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00853] =  Ifd35529b44c957737bf422127283c08e['h010a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00854] =  Ifd35529b44c957737bf422127283c08e['h010a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00855] =  Ifd35529b44c957737bf422127283c08e['h010aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00856] =  Ifd35529b44c957737bf422127283c08e['h010ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00857] =  Ifd35529b44c957737bf422127283c08e['h010ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00858] =  Ifd35529b44c957737bf422127283c08e['h010b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00859] =  Ifd35529b44c957737bf422127283c08e['h010b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0085a] =  Ifd35529b44c957737bf422127283c08e['h010b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0085b] =  Ifd35529b44c957737bf422127283c08e['h010b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0085c] =  Ifd35529b44c957737bf422127283c08e['h010b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0085d] =  Ifd35529b44c957737bf422127283c08e['h010ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0085e] =  Ifd35529b44c957737bf422127283c08e['h010bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0085f] =  Ifd35529b44c957737bf422127283c08e['h010be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00860] =  Ifd35529b44c957737bf422127283c08e['h010c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00861] =  Ifd35529b44c957737bf422127283c08e['h010c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00862] =  Ifd35529b44c957737bf422127283c08e['h010c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00863] =  Ifd35529b44c957737bf422127283c08e['h010c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00864] =  Ifd35529b44c957737bf422127283c08e['h010c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00865] =  Ifd35529b44c957737bf422127283c08e['h010ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00866] =  Ifd35529b44c957737bf422127283c08e['h010cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00867] =  Ifd35529b44c957737bf422127283c08e['h010ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00868] =  Ifd35529b44c957737bf422127283c08e['h010d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00869] =  Ifd35529b44c957737bf422127283c08e['h010d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0086a] =  Ifd35529b44c957737bf422127283c08e['h010d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0086b] =  Ifd35529b44c957737bf422127283c08e['h010d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0086c] =  Ifd35529b44c957737bf422127283c08e['h010d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0086d] =  Ifd35529b44c957737bf422127283c08e['h010da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0086e] =  Ifd35529b44c957737bf422127283c08e['h010dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0086f] =  Ifd35529b44c957737bf422127283c08e['h010de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00870] =  Ifd35529b44c957737bf422127283c08e['h010e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00871] =  Ifd35529b44c957737bf422127283c08e['h010e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00872] =  Ifd35529b44c957737bf422127283c08e['h010e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00873] =  Ifd35529b44c957737bf422127283c08e['h010e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00874] =  Ifd35529b44c957737bf422127283c08e['h010e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00875] =  Ifd35529b44c957737bf422127283c08e['h010ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00876] =  Ifd35529b44c957737bf422127283c08e['h010ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00877] =  Ifd35529b44c957737bf422127283c08e['h010ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00878] =  Ifd35529b44c957737bf422127283c08e['h010f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00879] =  Ifd35529b44c957737bf422127283c08e['h010f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0087a] =  Ifd35529b44c957737bf422127283c08e['h010f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0087b] =  Ifd35529b44c957737bf422127283c08e['h010f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0087c] =  Ifd35529b44c957737bf422127283c08e['h010f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0087d] =  Ifd35529b44c957737bf422127283c08e['h010fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0087e] =  Ifd35529b44c957737bf422127283c08e['h010fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0087f] =  Ifd35529b44c957737bf422127283c08e['h010fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00880] =  Ifd35529b44c957737bf422127283c08e['h01100] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00881] =  Ifd35529b44c957737bf422127283c08e['h01102] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00882] =  Ifd35529b44c957737bf422127283c08e['h01104] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00883] =  Ifd35529b44c957737bf422127283c08e['h01106] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00884] =  Ifd35529b44c957737bf422127283c08e['h01108] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00885] =  Ifd35529b44c957737bf422127283c08e['h0110a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00886] =  Ifd35529b44c957737bf422127283c08e['h0110c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00887] =  Ifd35529b44c957737bf422127283c08e['h0110e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00888] =  Ifd35529b44c957737bf422127283c08e['h01110] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00889] =  Ifd35529b44c957737bf422127283c08e['h01112] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0088a] =  Ifd35529b44c957737bf422127283c08e['h01114] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0088b] =  Ifd35529b44c957737bf422127283c08e['h01116] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0088c] =  Ifd35529b44c957737bf422127283c08e['h01118] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0088d] =  Ifd35529b44c957737bf422127283c08e['h0111a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0088e] =  Ifd35529b44c957737bf422127283c08e['h0111c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0088f] =  Ifd35529b44c957737bf422127283c08e['h0111e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00890] =  Ifd35529b44c957737bf422127283c08e['h01120] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00891] =  Ifd35529b44c957737bf422127283c08e['h01122] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00892] =  Ifd35529b44c957737bf422127283c08e['h01124] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00893] =  Ifd35529b44c957737bf422127283c08e['h01126] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00894] =  Ifd35529b44c957737bf422127283c08e['h01128] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00895] =  Ifd35529b44c957737bf422127283c08e['h0112a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00896] =  Ifd35529b44c957737bf422127283c08e['h0112c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00897] =  Ifd35529b44c957737bf422127283c08e['h0112e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00898] =  Ifd35529b44c957737bf422127283c08e['h01130] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00899] =  Ifd35529b44c957737bf422127283c08e['h01132] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0089a] =  Ifd35529b44c957737bf422127283c08e['h01134] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0089b] =  Ifd35529b44c957737bf422127283c08e['h01136] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0089c] =  Ifd35529b44c957737bf422127283c08e['h01138] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0089d] =  Ifd35529b44c957737bf422127283c08e['h0113a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0089e] =  Ifd35529b44c957737bf422127283c08e['h0113c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0089f] =  Ifd35529b44c957737bf422127283c08e['h0113e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008a0] =  Ifd35529b44c957737bf422127283c08e['h01140] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008a1] =  Ifd35529b44c957737bf422127283c08e['h01142] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008a2] =  Ifd35529b44c957737bf422127283c08e['h01144] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008a3] =  Ifd35529b44c957737bf422127283c08e['h01146] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008a4] =  Ifd35529b44c957737bf422127283c08e['h01148] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008a5] =  Ifd35529b44c957737bf422127283c08e['h0114a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008a6] =  Ifd35529b44c957737bf422127283c08e['h0114c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008a7] =  Ifd35529b44c957737bf422127283c08e['h0114e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008a8] =  Ifd35529b44c957737bf422127283c08e['h01150] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008a9] =  Ifd35529b44c957737bf422127283c08e['h01152] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008aa] =  Ifd35529b44c957737bf422127283c08e['h01154] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008ab] =  Ifd35529b44c957737bf422127283c08e['h01156] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008ac] =  Ifd35529b44c957737bf422127283c08e['h01158] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008ad] =  Ifd35529b44c957737bf422127283c08e['h0115a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008ae] =  Ifd35529b44c957737bf422127283c08e['h0115c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008af] =  Ifd35529b44c957737bf422127283c08e['h0115e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008b0] =  Ifd35529b44c957737bf422127283c08e['h01160] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008b1] =  Ifd35529b44c957737bf422127283c08e['h01162] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008b2] =  Ifd35529b44c957737bf422127283c08e['h01164] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008b3] =  Ifd35529b44c957737bf422127283c08e['h01166] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008b4] =  Ifd35529b44c957737bf422127283c08e['h01168] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008b5] =  Ifd35529b44c957737bf422127283c08e['h0116a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008b6] =  Ifd35529b44c957737bf422127283c08e['h0116c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008b7] =  Ifd35529b44c957737bf422127283c08e['h0116e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008b8] =  Ifd35529b44c957737bf422127283c08e['h01170] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008b9] =  Ifd35529b44c957737bf422127283c08e['h01172] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008ba] =  Ifd35529b44c957737bf422127283c08e['h01174] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008bb] =  Ifd35529b44c957737bf422127283c08e['h01176] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008bc] =  Ifd35529b44c957737bf422127283c08e['h01178] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008bd] =  Ifd35529b44c957737bf422127283c08e['h0117a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008be] =  Ifd35529b44c957737bf422127283c08e['h0117c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008bf] =  Ifd35529b44c957737bf422127283c08e['h0117e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008c0] =  Ifd35529b44c957737bf422127283c08e['h01180] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008c1] =  Ifd35529b44c957737bf422127283c08e['h01182] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008c2] =  Ifd35529b44c957737bf422127283c08e['h01184] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008c3] =  Ifd35529b44c957737bf422127283c08e['h01186] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008c4] =  Ifd35529b44c957737bf422127283c08e['h01188] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008c5] =  Ifd35529b44c957737bf422127283c08e['h0118a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008c6] =  Ifd35529b44c957737bf422127283c08e['h0118c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008c7] =  Ifd35529b44c957737bf422127283c08e['h0118e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008c8] =  Ifd35529b44c957737bf422127283c08e['h01190] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008c9] =  Ifd35529b44c957737bf422127283c08e['h01192] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008ca] =  Ifd35529b44c957737bf422127283c08e['h01194] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008cb] =  Ifd35529b44c957737bf422127283c08e['h01196] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008cc] =  Ifd35529b44c957737bf422127283c08e['h01198] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008cd] =  Ifd35529b44c957737bf422127283c08e['h0119a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008ce] =  Ifd35529b44c957737bf422127283c08e['h0119c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008cf] =  Ifd35529b44c957737bf422127283c08e['h0119e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008d0] =  Ifd35529b44c957737bf422127283c08e['h011a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008d1] =  Ifd35529b44c957737bf422127283c08e['h011a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008d2] =  Ifd35529b44c957737bf422127283c08e['h011a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008d3] =  Ifd35529b44c957737bf422127283c08e['h011a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008d4] =  Ifd35529b44c957737bf422127283c08e['h011a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008d5] =  Ifd35529b44c957737bf422127283c08e['h011aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008d6] =  Ifd35529b44c957737bf422127283c08e['h011ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008d7] =  Ifd35529b44c957737bf422127283c08e['h011ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008d8] =  Ifd35529b44c957737bf422127283c08e['h011b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008d9] =  Ifd35529b44c957737bf422127283c08e['h011b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008da] =  Ifd35529b44c957737bf422127283c08e['h011b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008db] =  Ifd35529b44c957737bf422127283c08e['h011b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008dc] =  Ifd35529b44c957737bf422127283c08e['h011b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008dd] =  Ifd35529b44c957737bf422127283c08e['h011ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008de] =  Ifd35529b44c957737bf422127283c08e['h011bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008df] =  Ifd35529b44c957737bf422127283c08e['h011be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008e0] =  Ifd35529b44c957737bf422127283c08e['h011c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008e1] =  Ifd35529b44c957737bf422127283c08e['h011c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008e2] =  Ifd35529b44c957737bf422127283c08e['h011c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008e3] =  Ifd35529b44c957737bf422127283c08e['h011c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008e4] =  Ifd35529b44c957737bf422127283c08e['h011c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008e5] =  Ifd35529b44c957737bf422127283c08e['h011ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008e6] =  Ifd35529b44c957737bf422127283c08e['h011cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008e7] =  Ifd35529b44c957737bf422127283c08e['h011ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008e8] =  Ifd35529b44c957737bf422127283c08e['h011d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008e9] =  Ifd35529b44c957737bf422127283c08e['h011d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008ea] =  Ifd35529b44c957737bf422127283c08e['h011d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008eb] =  Ifd35529b44c957737bf422127283c08e['h011d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008ec] =  Ifd35529b44c957737bf422127283c08e['h011d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008ed] =  Ifd35529b44c957737bf422127283c08e['h011da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008ee] =  Ifd35529b44c957737bf422127283c08e['h011dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008ef] =  Ifd35529b44c957737bf422127283c08e['h011de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008f0] =  Ifd35529b44c957737bf422127283c08e['h011e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008f1] =  Ifd35529b44c957737bf422127283c08e['h011e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008f2] =  Ifd35529b44c957737bf422127283c08e['h011e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008f3] =  Ifd35529b44c957737bf422127283c08e['h011e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008f4] =  Ifd35529b44c957737bf422127283c08e['h011e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008f5] =  Ifd35529b44c957737bf422127283c08e['h011ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008f6] =  Ifd35529b44c957737bf422127283c08e['h011ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008f7] =  Ifd35529b44c957737bf422127283c08e['h011ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008f8] =  Ifd35529b44c957737bf422127283c08e['h011f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008f9] =  Ifd35529b44c957737bf422127283c08e['h011f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008fa] =  Ifd35529b44c957737bf422127283c08e['h011f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008fb] =  Ifd35529b44c957737bf422127283c08e['h011f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008fc] =  Ifd35529b44c957737bf422127283c08e['h011f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008fd] =  Ifd35529b44c957737bf422127283c08e['h011fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008fe] =  Ifd35529b44c957737bf422127283c08e['h011fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h008ff] =  Ifd35529b44c957737bf422127283c08e['h011fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00900] =  Ifd35529b44c957737bf422127283c08e['h01200] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00901] =  Ifd35529b44c957737bf422127283c08e['h01202] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00902] =  Ifd35529b44c957737bf422127283c08e['h01204] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00903] =  Ifd35529b44c957737bf422127283c08e['h01206] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00904] =  Ifd35529b44c957737bf422127283c08e['h01208] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00905] =  Ifd35529b44c957737bf422127283c08e['h0120a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00906] =  Ifd35529b44c957737bf422127283c08e['h0120c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00907] =  Ifd35529b44c957737bf422127283c08e['h0120e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00908] =  Ifd35529b44c957737bf422127283c08e['h01210] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00909] =  Ifd35529b44c957737bf422127283c08e['h01212] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0090a] =  Ifd35529b44c957737bf422127283c08e['h01214] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0090b] =  Ifd35529b44c957737bf422127283c08e['h01216] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0090c] =  Ifd35529b44c957737bf422127283c08e['h01218] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0090d] =  Ifd35529b44c957737bf422127283c08e['h0121a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0090e] =  Ifd35529b44c957737bf422127283c08e['h0121c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0090f] =  Ifd35529b44c957737bf422127283c08e['h0121e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00910] =  Ifd35529b44c957737bf422127283c08e['h01220] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00911] =  Ifd35529b44c957737bf422127283c08e['h01222] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00912] =  Ifd35529b44c957737bf422127283c08e['h01224] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00913] =  Ifd35529b44c957737bf422127283c08e['h01226] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00914] =  Ifd35529b44c957737bf422127283c08e['h01228] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00915] =  Ifd35529b44c957737bf422127283c08e['h0122a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00916] =  Ifd35529b44c957737bf422127283c08e['h0122c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00917] =  Ifd35529b44c957737bf422127283c08e['h0122e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00918] =  Ifd35529b44c957737bf422127283c08e['h01230] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00919] =  Ifd35529b44c957737bf422127283c08e['h01232] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0091a] =  Ifd35529b44c957737bf422127283c08e['h01234] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0091b] =  Ifd35529b44c957737bf422127283c08e['h01236] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0091c] =  Ifd35529b44c957737bf422127283c08e['h01238] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0091d] =  Ifd35529b44c957737bf422127283c08e['h0123a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0091e] =  Ifd35529b44c957737bf422127283c08e['h0123c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0091f] =  Ifd35529b44c957737bf422127283c08e['h0123e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00920] =  Ifd35529b44c957737bf422127283c08e['h01240] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00921] =  Ifd35529b44c957737bf422127283c08e['h01242] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00922] =  Ifd35529b44c957737bf422127283c08e['h01244] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00923] =  Ifd35529b44c957737bf422127283c08e['h01246] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00924] =  Ifd35529b44c957737bf422127283c08e['h01248] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00925] =  Ifd35529b44c957737bf422127283c08e['h0124a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00926] =  Ifd35529b44c957737bf422127283c08e['h0124c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00927] =  Ifd35529b44c957737bf422127283c08e['h0124e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00928] =  Ifd35529b44c957737bf422127283c08e['h01250] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00929] =  Ifd35529b44c957737bf422127283c08e['h01252] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0092a] =  Ifd35529b44c957737bf422127283c08e['h01254] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0092b] =  Ifd35529b44c957737bf422127283c08e['h01256] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0092c] =  Ifd35529b44c957737bf422127283c08e['h01258] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0092d] =  Ifd35529b44c957737bf422127283c08e['h0125a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0092e] =  Ifd35529b44c957737bf422127283c08e['h0125c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0092f] =  Ifd35529b44c957737bf422127283c08e['h0125e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00930] =  Ifd35529b44c957737bf422127283c08e['h01260] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00931] =  Ifd35529b44c957737bf422127283c08e['h01262] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00932] =  Ifd35529b44c957737bf422127283c08e['h01264] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00933] =  Ifd35529b44c957737bf422127283c08e['h01266] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00934] =  Ifd35529b44c957737bf422127283c08e['h01268] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00935] =  Ifd35529b44c957737bf422127283c08e['h0126a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00936] =  Ifd35529b44c957737bf422127283c08e['h0126c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00937] =  Ifd35529b44c957737bf422127283c08e['h0126e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00938] =  Ifd35529b44c957737bf422127283c08e['h01270] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00939] =  Ifd35529b44c957737bf422127283c08e['h01272] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0093a] =  Ifd35529b44c957737bf422127283c08e['h01274] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0093b] =  Ifd35529b44c957737bf422127283c08e['h01276] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0093c] =  Ifd35529b44c957737bf422127283c08e['h01278] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0093d] =  Ifd35529b44c957737bf422127283c08e['h0127a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0093e] =  Ifd35529b44c957737bf422127283c08e['h0127c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0093f] =  Ifd35529b44c957737bf422127283c08e['h0127e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00940] =  Ifd35529b44c957737bf422127283c08e['h01280] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00941] =  Ifd35529b44c957737bf422127283c08e['h01282] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00942] =  Ifd35529b44c957737bf422127283c08e['h01284] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00943] =  Ifd35529b44c957737bf422127283c08e['h01286] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00944] =  Ifd35529b44c957737bf422127283c08e['h01288] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00945] =  Ifd35529b44c957737bf422127283c08e['h0128a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00946] =  Ifd35529b44c957737bf422127283c08e['h0128c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00947] =  Ifd35529b44c957737bf422127283c08e['h0128e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00948] =  Ifd35529b44c957737bf422127283c08e['h01290] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00949] =  Ifd35529b44c957737bf422127283c08e['h01292] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0094a] =  Ifd35529b44c957737bf422127283c08e['h01294] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0094b] =  Ifd35529b44c957737bf422127283c08e['h01296] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0094c] =  Ifd35529b44c957737bf422127283c08e['h01298] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0094d] =  Ifd35529b44c957737bf422127283c08e['h0129a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0094e] =  Ifd35529b44c957737bf422127283c08e['h0129c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0094f] =  Ifd35529b44c957737bf422127283c08e['h0129e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00950] =  Ifd35529b44c957737bf422127283c08e['h012a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00951] =  Ifd35529b44c957737bf422127283c08e['h012a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00952] =  Ifd35529b44c957737bf422127283c08e['h012a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00953] =  Ifd35529b44c957737bf422127283c08e['h012a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00954] =  Ifd35529b44c957737bf422127283c08e['h012a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00955] =  Ifd35529b44c957737bf422127283c08e['h012aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00956] =  Ifd35529b44c957737bf422127283c08e['h012ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00957] =  Ifd35529b44c957737bf422127283c08e['h012ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00958] =  Ifd35529b44c957737bf422127283c08e['h012b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00959] =  Ifd35529b44c957737bf422127283c08e['h012b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0095a] =  Ifd35529b44c957737bf422127283c08e['h012b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0095b] =  Ifd35529b44c957737bf422127283c08e['h012b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0095c] =  Ifd35529b44c957737bf422127283c08e['h012b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0095d] =  Ifd35529b44c957737bf422127283c08e['h012ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0095e] =  Ifd35529b44c957737bf422127283c08e['h012bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0095f] =  Ifd35529b44c957737bf422127283c08e['h012be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00960] =  Ifd35529b44c957737bf422127283c08e['h012c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00961] =  Ifd35529b44c957737bf422127283c08e['h012c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00962] =  Ifd35529b44c957737bf422127283c08e['h012c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00963] =  Ifd35529b44c957737bf422127283c08e['h012c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00964] =  Ifd35529b44c957737bf422127283c08e['h012c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00965] =  Ifd35529b44c957737bf422127283c08e['h012ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00966] =  Ifd35529b44c957737bf422127283c08e['h012cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00967] =  Ifd35529b44c957737bf422127283c08e['h012ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00968] =  Ifd35529b44c957737bf422127283c08e['h012d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00969] =  Ifd35529b44c957737bf422127283c08e['h012d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0096a] =  Ifd35529b44c957737bf422127283c08e['h012d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0096b] =  Ifd35529b44c957737bf422127283c08e['h012d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0096c] =  Ifd35529b44c957737bf422127283c08e['h012d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0096d] =  Ifd35529b44c957737bf422127283c08e['h012da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0096e] =  Ifd35529b44c957737bf422127283c08e['h012dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0096f] =  Ifd35529b44c957737bf422127283c08e['h012de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00970] =  Ifd35529b44c957737bf422127283c08e['h012e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00971] =  Ifd35529b44c957737bf422127283c08e['h012e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00972] =  Ifd35529b44c957737bf422127283c08e['h012e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00973] =  Ifd35529b44c957737bf422127283c08e['h012e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00974] =  Ifd35529b44c957737bf422127283c08e['h012e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00975] =  Ifd35529b44c957737bf422127283c08e['h012ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00976] =  Ifd35529b44c957737bf422127283c08e['h012ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00977] =  Ifd35529b44c957737bf422127283c08e['h012ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00978] =  Ifd35529b44c957737bf422127283c08e['h012f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00979] =  Ifd35529b44c957737bf422127283c08e['h012f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0097a] =  Ifd35529b44c957737bf422127283c08e['h012f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0097b] =  Ifd35529b44c957737bf422127283c08e['h012f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0097c] =  Ifd35529b44c957737bf422127283c08e['h012f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0097d] =  Ifd35529b44c957737bf422127283c08e['h012fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0097e] =  Ifd35529b44c957737bf422127283c08e['h012fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0097f] =  Ifd35529b44c957737bf422127283c08e['h012fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00980] =  Ifd35529b44c957737bf422127283c08e['h01300] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00981] =  Ifd35529b44c957737bf422127283c08e['h01302] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00982] =  Ifd35529b44c957737bf422127283c08e['h01304] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00983] =  Ifd35529b44c957737bf422127283c08e['h01306] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00984] =  Ifd35529b44c957737bf422127283c08e['h01308] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00985] =  Ifd35529b44c957737bf422127283c08e['h0130a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00986] =  Ifd35529b44c957737bf422127283c08e['h0130c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00987] =  Ifd35529b44c957737bf422127283c08e['h0130e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00988] =  Ifd35529b44c957737bf422127283c08e['h01310] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00989] =  Ifd35529b44c957737bf422127283c08e['h01312] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0098a] =  Ifd35529b44c957737bf422127283c08e['h01314] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0098b] =  Ifd35529b44c957737bf422127283c08e['h01316] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0098c] =  Ifd35529b44c957737bf422127283c08e['h01318] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0098d] =  Ifd35529b44c957737bf422127283c08e['h0131a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0098e] =  Ifd35529b44c957737bf422127283c08e['h0131c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0098f] =  Ifd35529b44c957737bf422127283c08e['h0131e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00990] =  Ifd35529b44c957737bf422127283c08e['h01320] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00991] =  Ifd35529b44c957737bf422127283c08e['h01322] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00992] =  Ifd35529b44c957737bf422127283c08e['h01324] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00993] =  Ifd35529b44c957737bf422127283c08e['h01326] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00994] =  Ifd35529b44c957737bf422127283c08e['h01328] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00995] =  Ifd35529b44c957737bf422127283c08e['h0132a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00996] =  Ifd35529b44c957737bf422127283c08e['h0132c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00997] =  Ifd35529b44c957737bf422127283c08e['h0132e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00998] =  Ifd35529b44c957737bf422127283c08e['h01330] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00999] =  Ifd35529b44c957737bf422127283c08e['h01332] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0099a] =  Ifd35529b44c957737bf422127283c08e['h01334] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0099b] =  Ifd35529b44c957737bf422127283c08e['h01336] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0099c] =  Ifd35529b44c957737bf422127283c08e['h01338] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0099d] =  Ifd35529b44c957737bf422127283c08e['h0133a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0099e] =  Ifd35529b44c957737bf422127283c08e['h0133c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0099f] =  Ifd35529b44c957737bf422127283c08e['h0133e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009a0] =  Ifd35529b44c957737bf422127283c08e['h01340] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009a1] =  Ifd35529b44c957737bf422127283c08e['h01342] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009a2] =  Ifd35529b44c957737bf422127283c08e['h01344] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009a3] =  Ifd35529b44c957737bf422127283c08e['h01346] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009a4] =  Ifd35529b44c957737bf422127283c08e['h01348] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009a5] =  Ifd35529b44c957737bf422127283c08e['h0134a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009a6] =  Ifd35529b44c957737bf422127283c08e['h0134c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009a7] =  Ifd35529b44c957737bf422127283c08e['h0134e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009a8] =  Ifd35529b44c957737bf422127283c08e['h01350] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009a9] =  Ifd35529b44c957737bf422127283c08e['h01352] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009aa] =  Ifd35529b44c957737bf422127283c08e['h01354] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009ab] =  Ifd35529b44c957737bf422127283c08e['h01356] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009ac] =  Ifd35529b44c957737bf422127283c08e['h01358] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009ad] =  Ifd35529b44c957737bf422127283c08e['h0135a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009ae] =  Ifd35529b44c957737bf422127283c08e['h0135c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009af] =  Ifd35529b44c957737bf422127283c08e['h0135e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009b0] =  Ifd35529b44c957737bf422127283c08e['h01360] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009b1] =  Ifd35529b44c957737bf422127283c08e['h01362] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009b2] =  Ifd35529b44c957737bf422127283c08e['h01364] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009b3] =  Ifd35529b44c957737bf422127283c08e['h01366] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009b4] =  Ifd35529b44c957737bf422127283c08e['h01368] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009b5] =  Ifd35529b44c957737bf422127283c08e['h0136a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009b6] =  Ifd35529b44c957737bf422127283c08e['h0136c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009b7] =  Ifd35529b44c957737bf422127283c08e['h0136e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009b8] =  Ifd35529b44c957737bf422127283c08e['h01370] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009b9] =  Ifd35529b44c957737bf422127283c08e['h01372] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009ba] =  Ifd35529b44c957737bf422127283c08e['h01374] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009bb] =  Ifd35529b44c957737bf422127283c08e['h01376] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009bc] =  Ifd35529b44c957737bf422127283c08e['h01378] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009bd] =  Ifd35529b44c957737bf422127283c08e['h0137a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009be] =  Ifd35529b44c957737bf422127283c08e['h0137c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009bf] =  Ifd35529b44c957737bf422127283c08e['h0137e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009c0] =  Ifd35529b44c957737bf422127283c08e['h01380] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009c1] =  Ifd35529b44c957737bf422127283c08e['h01382] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009c2] =  Ifd35529b44c957737bf422127283c08e['h01384] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009c3] =  Ifd35529b44c957737bf422127283c08e['h01386] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009c4] =  Ifd35529b44c957737bf422127283c08e['h01388] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009c5] =  Ifd35529b44c957737bf422127283c08e['h0138a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009c6] =  Ifd35529b44c957737bf422127283c08e['h0138c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009c7] =  Ifd35529b44c957737bf422127283c08e['h0138e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009c8] =  Ifd35529b44c957737bf422127283c08e['h01390] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009c9] =  Ifd35529b44c957737bf422127283c08e['h01392] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009ca] =  Ifd35529b44c957737bf422127283c08e['h01394] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009cb] =  Ifd35529b44c957737bf422127283c08e['h01396] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009cc] =  Ifd35529b44c957737bf422127283c08e['h01398] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009cd] =  Ifd35529b44c957737bf422127283c08e['h0139a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009ce] =  Ifd35529b44c957737bf422127283c08e['h0139c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009cf] =  Ifd35529b44c957737bf422127283c08e['h0139e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009d0] =  Ifd35529b44c957737bf422127283c08e['h013a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009d1] =  Ifd35529b44c957737bf422127283c08e['h013a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009d2] =  Ifd35529b44c957737bf422127283c08e['h013a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009d3] =  Ifd35529b44c957737bf422127283c08e['h013a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009d4] =  Ifd35529b44c957737bf422127283c08e['h013a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009d5] =  Ifd35529b44c957737bf422127283c08e['h013aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009d6] =  Ifd35529b44c957737bf422127283c08e['h013ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009d7] =  Ifd35529b44c957737bf422127283c08e['h013ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009d8] =  Ifd35529b44c957737bf422127283c08e['h013b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009d9] =  Ifd35529b44c957737bf422127283c08e['h013b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009da] =  Ifd35529b44c957737bf422127283c08e['h013b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009db] =  Ifd35529b44c957737bf422127283c08e['h013b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009dc] =  Ifd35529b44c957737bf422127283c08e['h013b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009dd] =  Ifd35529b44c957737bf422127283c08e['h013ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009de] =  Ifd35529b44c957737bf422127283c08e['h013bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009df] =  Ifd35529b44c957737bf422127283c08e['h013be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009e0] =  Ifd35529b44c957737bf422127283c08e['h013c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009e1] =  Ifd35529b44c957737bf422127283c08e['h013c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009e2] =  Ifd35529b44c957737bf422127283c08e['h013c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009e3] =  Ifd35529b44c957737bf422127283c08e['h013c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009e4] =  Ifd35529b44c957737bf422127283c08e['h013c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009e5] =  Ifd35529b44c957737bf422127283c08e['h013ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009e6] =  Ifd35529b44c957737bf422127283c08e['h013cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009e7] =  Ifd35529b44c957737bf422127283c08e['h013ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009e8] =  Ifd35529b44c957737bf422127283c08e['h013d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009e9] =  Ifd35529b44c957737bf422127283c08e['h013d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009ea] =  Ifd35529b44c957737bf422127283c08e['h013d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009eb] =  Ifd35529b44c957737bf422127283c08e['h013d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009ec] =  Ifd35529b44c957737bf422127283c08e['h013d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009ed] =  Ifd35529b44c957737bf422127283c08e['h013da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009ee] =  Ifd35529b44c957737bf422127283c08e['h013dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009ef] =  Ifd35529b44c957737bf422127283c08e['h013de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009f0] =  Ifd35529b44c957737bf422127283c08e['h013e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009f1] =  Ifd35529b44c957737bf422127283c08e['h013e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009f2] =  Ifd35529b44c957737bf422127283c08e['h013e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009f3] =  Ifd35529b44c957737bf422127283c08e['h013e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009f4] =  Ifd35529b44c957737bf422127283c08e['h013e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009f5] =  Ifd35529b44c957737bf422127283c08e['h013ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009f6] =  Ifd35529b44c957737bf422127283c08e['h013ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009f7] =  Ifd35529b44c957737bf422127283c08e['h013ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009f8] =  Ifd35529b44c957737bf422127283c08e['h013f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009f9] =  Ifd35529b44c957737bf422127283c08e['h013f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009fa] =  Ifd35529b44c957737bf422127283c08e['h013f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009fb] =  Ifd35529b44c957737bf422127283c08e['h013f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009fc] =  Ifd35529b44c957737bf422127283c08e['h013f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009fd] =  Ifd35529b44c957737bf422127283c08e['h013fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009fe] =  Ifd35529b44c957737bf422127283c08e['h013fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h009ff] =  Ifd35529b44c957737bf422127283c08e['h013fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a00] =  Ifd35529b44c957737bf422127283c08e['h01400] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a01] =  Ifd35529b44c957737bf422127283c08e['h01402] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a02] =  Ifd35529b44c957737bf422127283c08e['h01404] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a03] =  Ifd35529b44c957737bf422127283c08e['h01406] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a04] =  Ifd35529b44c957737bf422127283c08e['h01408] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a05] =  Ifd35529b44c957737bf422127283c08e['h0140a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a06] =  Ifd35529b44c957737bf422127283c08e['h0140c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a07] =  Ifd35529b44c957737bf422127283c08e['h0140e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a08] =  Ifd35529b44c957737bf422127283c08e['h01410] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a09] =  Ifd35529b44c957737bf422127283c08e['h01412] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a0a] =  Ifd35529b44c957737bf422127283c08e['h01414] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a0b] =  Ifd35529b44c957737bf422127283c08e['h01416] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a0c] =  Ifd35529b44c957737bf422127283c08e['h01418] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a0d] =  Ifd35529b44c957737bf422127283c08e['h0141a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a0e] =  Ifd35529b44c957737bf422127283c08e['h0141c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a0f] =  Ifd35529b44c957737bf422127283c08e['h0141e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a10] =  Ifd35529b44c957737bf422127283c08e['h01420] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a11] =  Ifd35529b44c957737bf422127283c08e['h01422] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a12] =  Ifd35529b44c957737bf422127283c08e['h01424] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a13] =  Ifd35529b44c957737bf422127283c08e['h01426] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a14] =  Ifd35529b44c957737bf422127283c08e['h01428] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a15] =  Ifd35529b44c957737bf422127283c08e['h0142a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a16] =  Ifd35529b44c957737bf422127283c08e['h0142c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a17] =  Ifd35529b44c957737bf422127283c08e['h0142e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a18] =  Ifd35529b44c957737bf422127283c08e['h01430] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a19] =  Ifd35529b44c957737bf422127283c08e['h01432] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a1a] =  Ifd35529b44c957737bf422127283c08e['h01434] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a1b] =  Ifd35529b44c957737bf422127283c08e['h01436] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a1c] =  Ifd35529b44c957737bf422127283c08e['h01438] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a1d] =  Ifd35529b44c957737bf422127283c08e['h0143a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a1e] =  Ifd35529b44c957737bf422127283c08e['h0143c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a1f] =  Ifd35529b44c957737bf422127283c08e['h0143e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a20] =  Ifd35529b44c957737bf422127283c08e['h01440] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a21] =  Ifd35529b44c957737bf422127283c08e['h01442] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a22] =  Ifd35529b44c957737bf422127283c08e['h01444] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a23] =  Ifd35529b44c957737bf422127283c08e['h01446] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a24] =  Ifd35529b44c957737bf422127283c08e['h01448] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a25] =  Ifd35529b44c957737bf422127283c08e['h0144a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a26] =  Ifd35529b44c957737bf422127283c08e['h0144c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a27] =  Ifd35529b44c957737bf422127283c08e['h0144e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a28] =  Ifd35529b44c957737bf422127283c08e['h01450] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a29] =  Ifd35529b44c957737bf422127283c08e['h01452] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a2a] =  Ifd35529b44c957737bf422127283c08e['h01454] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a2b] =  Ifd35529b44c957737bf422127283c08e['h01456] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a2c] =  Ifd35529b44c957737bf422127283c08e['h01458] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a2d] =  Ifd35529b44c957737bf422127283c08e['h0145a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a2e] =  Ifd35529b44c957737bf422127283c08e['h0145c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a2f] =  Ifd35529b44c957737bf422127283c08e['h0145e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a30] =  Ifd35529b44c957737bf422127283c08e['h01460] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a31] =  Ifd35529b44c957737bf422127283c08e['h01462] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a32] =  Ifd35529b44c957737bf422127283c08e['h01464] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a33] =  Ifd35529b44c957737bf422127283c08e['h01466] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a34] =  Ifd35529b44c957737bf422127283c08e['h01468] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a35] =  Ifd35529b44c957737bf422127283c08e['h0146a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a36] =  Ifd35529b44c957737bf422127283c08e['h0146c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a37] =  Ifd35529b44c957737bf422127283c08e['h0146e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a38] =  Ifd35529b44c957737bf422127283c08e['h01470] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a39] =  Ifd35529b44c957737bf422127283c08e['h01472] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a3a] =  Ifd35529b44c957737bf422127283c08e['h01474] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a3b] =  Ifd35529b44c957737bf422127283c08e['h01476] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a3c] =  Ifd35529b44c957737bf422127283c08e['h01478] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a3d] =  Ifd35529b44c957737bf422127283c08e['h0147a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a3e] =  Ifd35529b44c957737bf422127283c08e['h0147c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a3f] =  Ifd35529b44c957737bf422127283c08e['h0147e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a40] =  Ifd35529b44c957737bf422127283c08e['h01480] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a41] =  Ifd35529b44c957737bf422127283c08e['h01482] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a42] =  Ifd35529b44c957737bf422127283c08e['h01484] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a43] =  Ifd35529b44c957737bf422127283c08e['h01486] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a44] =  Ifd35529b44c957737bf422127283c08e['h01488] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a45] =  Ifd35529b44c957737bf422127283c08e['h0148a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a46] =  Ifd35529b44c957737bf422127283c08e['h0148c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a47] =  Ifd35529b44c957737bf422127283c08e['h0148e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a48] =  Ifd35529b44c957737bf422127283c08e['h01490] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a49] =  Ifd35529b44c957737bf422127283c08e['h01492] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a4a] =  Ifd35529b44c957737bf422127283c08e['h01494] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a4b] =  Ifd35529b44c957737bf422127283c08e['h01496] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a4c] =  Ifd35529b44c957737bf422127283c08e['h01498] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a4d] =  Ifd35529b44c957737bf422127283c08e['h0149a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a4e] =  Ifd35529b44c957737bf422127283c08e['h0149c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a4f] =  Ifd35529b44c957737bf422127283c08e['h0149e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a50] =  Ifd35529b44c957737bf422127283c08e['h014a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a51] =  Ifd35529b44c957737bf422127283c08e['h014a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a52] =  Ifd35529b44c957737bf422127283c08e['h014a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a53] =  Ifd35529b44c957737bf422127283c08e['h014a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a54] =  Ifd35529b44c957737bf422127283c08e['h014a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a55] =  Ifd35529b44c957737bf422127283c08e['h014aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a56] =  Ifd35529b44c957737bf422127283c08e['h014ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a57] =  Ifd35529b44c957737bf422127283c08e['h014ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a58] =  Ifd35529b44c957737bf422127283c08e['h014b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a59] =  Ifd35529b44c957737bf422127283c08e['h014b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a5a] =  Ifd35529b44c957737bf422127283c08e['h014b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a5b] =  Ifd35529b44c957737bf422127283c08e['h014b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a5c] =  Ifd35529b44c957737bf422127283c08e['h014b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a5d] =  Ifd35529b44c957737bf422127283c08e['h014ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a5e] =  Ifd35529b44c957737bf422127283c08e['h014bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a5f] =  Ifd35529b44c957737bf422127283c08e['h014be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a60] =  Ifd35529b44c957737bf422127283c08e['h014c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a61] =  Ifd35529b44c957737bf422127283c08e['h014c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a62] =  Ifd35529b44c957737bf422127283c08e['h014c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a63] =  Ifd35529b44c957737bf422127283c08e['h014c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a64] =  Ifd35529b44c957737bf422127283c08e['h014c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a65] =  Ifd35529b44c957737bf422127283c08e['h014ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a66] =  Ifd35529b44c957737bf422127283c08e['h014cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a67] =  Ifd35529b44c957737bf422127283c08e['h014ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a68] =  Ifd35529b44c957737bf422127283c08e['h014d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a69] =  Ifd35529b44c957737bf422127283c08e['h014d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a6a] =  Ifd35529b44c957737bf422127283c08e['h014d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a6b] =  Ifd35529b44c957737bf422127283c08e['h014d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a6c] =  Ifd35529b44c957737bf422127283c08e['h014d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a6d] =  Ifd35529b44c957737bf422127283c08e['h014da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a6e] =  Ifd35529b44c957737bf422127283c08e['h014dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a6f] =  Ifd35529b44c957737bf422127283c08e['h014de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a70] =  Ifd35529b44c957737bf422127283c08e['h014e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a71] =  Ifd35529b44c957737bf422127283c08e['h014e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a72] =  Ifd35529b44c957737bf422127283c08e['h014e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a73] =  Ifd35529b44c957737bf422127283c08e['h014e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a74] =  Ifd35529b44c957737bf422127283c08e['h014e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a75] =  Ifd35529b44c957737bf422127283c08e['h014ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a76] =  Ifd35529b44c957737bf422127283c08e['h014ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a77] =  Ifd35529b44c957737bf422127283c08e['h014ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a78] =  Ifd35529b44c957737bf422127283c08e['h014f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a79] =  Ifd35529b44c957737bf422127283c08e['h014f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a7a] =  Ifd35529b44c957737bf422127283c08e['h014f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a7b] =  Ifd35529b44c957737bf422127283c08e['h014f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a7c] =  Ifd35529b44c957737bf422127283c08e['h014f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a7d] =  Ifd35529b44c957737bf422127283c08e['h014fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a7e] =  Ifd35529b44c957737bf422127283c08e['h014fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a7f] =  Ifd35529b44c957737bf422127283c08e['h014fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a80] =  Ifd35529b44c957737bf422127283c08e['h01500] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a81] =  Ifd35529b44c957737bf422127283c08e['h01502] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a82] =  Ifd35529b44c957737bf422127283c08e['h01504] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a83] =  Ifd35529b44c957737bf422127283c08e['h01506] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a84] =  Ifd35529b44c957737bf422127283c08e['h01508] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a85] =  Ifd35529b44c957737bf422127283c08e['h0150a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a86] =  Ifd35529b44c957737bf422127283c08e['h0150c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a87] =  Ifd35529b44c957737bf422127283c08e['h0150e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a88] =  Ifd35529b44c957737bf422127283c08e['h01510] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a89] =  Ifd35529b44c957737bf422127283c08e['h01512] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a8a] =  Ifd35529b44c957737bf422127283c08e['h01514] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a8b] =  Ifd35529b44c957737bf422127283c08e['h01516] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a8c] =  Ifd35529b44c957737bf422127283c08e['h01518] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a8d] =  Ifd35529b44c957737bf422127283c08e['h0151a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a8e] =  Ifd35529b44c957737bf422127283c08e['h0151c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a8f] =  Ifd35529b44c957737bf422127283c08e['h0151e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a90] =  Ifd35529b44c957737bf422127283c08e['h01520] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a91] =  Ifd35529b44c957737bf422127283c08e['h01522] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a92] =  Ifd35529b44c957737bf422127283c08e['h01524] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a93] =  Ifd35529b44c957737bf422127283c08e['h01526] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a94] =  Ifd35529b44c957737bf422127283c08e['h01528] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a95] =  Ifd35529b44c957737bf422127283c08e['h0152a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a96] =  Ifd35529b44c957737bf422127283c08e['h0152c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a97] =  Ifd35529b44c957737bf422127283c08e['h0152e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a98] =  Ifd35529b44c957737bf422127283c08e['h01530] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a99] =  Ifd35529b44c957737bf422127283c08e['h01532] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a9a] =  Ifd35529b44c957737bf422127283c08e['h01534] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a9b] =  Ifd35529b44c957737bf422127283c08e['h01536] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a9c] =  Ifd35529b44c957737bf422127283c08e['h01538] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a9d] =  Ifd35529b44c957737bf422127283c08e['h0153a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a9e] =  Ifd35529b44c957737bf422127283c08e['h0153c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00a9f] =  Ifd35529b44c957737bf422127283c08e['h0153e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00aa0] =  Ifd35529b44c957737bf422127283c08e['h01540] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00aa1] =  Ifd35529b44c957737bf422127283c08e['h01542] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00aa2] =  Ifd35529b44c957737bf422127283c08e['h01544] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00aa3] =  Ifd35529b44c957737bf422127283c08e['h01546] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00aa4] =  Ifd35529b44c957737bf422127283c08e['h01548] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00aa5] =  Ifd35529b44c957737bf422127283c08e['h0154a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00aa6] =  Ifd35529b44c957737bf422127283c08e['h0154c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00aa7] =  Ifd35529b44c957737bf422127283c08e['h0154e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00aa8] =  Ifd35529b44c957737bf422127283c08e['h01550] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00aa9] =  Ifd35529b44c957737bf422127283c08e['h01552] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00aaa] =  Ifd35529b44c957737bf422127283c08e['h01554] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00aab] =  Ifd35529b44c957737bf422127283c08e['h01556] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00aac] =  Ifd35529b44c957737bf422127283c08e['h01558] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00aad] =  Ifd35529b44c957737bf422127283c08e['h0155a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00aae] =  Ifd35529b44c957737bf422127283c08e['h0155c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00aaf] =  Ifd35529b44c957737bf422127283c08e['h0155e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ab0] =  Ifd35529b44c957737bf422127283c08e['h01560] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ab1] =  Ifd35529b44c957737bf422127283c08e['h01562] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ab2] =  Ifd35529b44c957737bf422127283c08e['h01564] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ab3] =  Ifd35529b44c957737bf422127283c08e['h01566] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ab4] =  Ifd35529b44c957737bf422127283c08e['h01568] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ab5] =  Ifd35529b44c957737bf422127283c08e['h0156a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ab6] =  Ifd35529b44c957737bf422127283c08e['h0156c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ab7] =  Ifd35529b44c957737bf422127283c08e['h0156e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ab8] =  Ifd35529b44c957737bf422127283c08e['h01570] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ab9] =  Ifd35529b44c957737bf422127283c08e['h01572] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00aba] =  Ifd35529b44c957737bf422127283c08e['h01574] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00abb] =  Ifd35529b44c957737bf422127283c08e['h01576] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00abc] =  Ifd35529b44c957737bf422127283c08e['h01578] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00abd] =  Ifd35529b44c957737bf422127283c08e['h0157a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00abe] =  Ifd35529b44c957737bf422127283c08e['h0157c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00abf] =  Ifd35529b44c957737bf422127283c08e['h0157e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ac0] =  Ifd35529b44c957737bf422127283c08e['h01580] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ac1] =  Ifd35529b44c957737bf422127283c08e['h01582] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ac2] =  Ifd35529b44c957737bf422127283c08e['h01584] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ac3] =  Ifd35529b44c957737bf422127283c08e['h01586] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ac4] =  Ifd35529b44c957737bf422127283c08e['h01588] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ac5] =  Ifd35529b44c957737bf422127283c08e['h0158a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ac6] =  Ifd35529b44c957737bf422127283c08e['h0158c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ac7] =  Ifd35529b44c957737bf422127283c08e['h0158e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ac8] =  Ifd35529b44c957737bf422127283c08e['h01590] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ac9] =  Ifd35529b44c957737bf422127283c08e['h01592] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00aca] =  Ifd35529b44c957737bf422127283c08e['h01594] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00acb] =  Ifd35529b44c957737bf422127283c08e['h01596] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00acc] =  Ifd35529b44c957737bf422127283c08e['h01598] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00acd] =  Ifd35529b44c957737bf422127283c08e['h0159a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ace] =  Ifd35529b44c957737bf422127283c08e['h0159c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00acf] =  Ifd35529b44c957737bf422127283c08e['h0159e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ad0] =  Ifd35529b44c957737bf422127283c08e['h015a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ad1] =  Ifd35529b44c957737bf422127283c08e['h015a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ad2] =  Ifd35529b44c957737bf422127283c08e['h015a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ad3] =  Ifd35529b44c957737bf422127283c08e['h015a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ad4] =  Ifd35529b44c957737bf422127283c08e['h015a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ad5] =  Ifd35529b44c957737bf422127283c08e['h015aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ad6] =  Ifd35529b44c957737bf422127283c08e['h015ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ad7] =  Ifd35529b44c957737bf422127283c08e['h015ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ad8] =  Ifd35529b44c957737bf422127283c08e['h015b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ad9] =  Ifd35529b44c957737bf422127283c08e['h015b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ada] =  Ifd35529b44c957737bf422127283c08e['h015b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00adb] =  Ifd35529b44c957737bf422127283c08e['h015b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00adc] =  Ifd35529b44c957737bf422127283c08e['h015b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00add] =  Ifd35529b44c957737bf422127283c08e['h015ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ade] =  Ifd35529b44c957737bf422127283c08e['h015bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00adf] =  Ifd35529b44c957737bf422127283c08e['h015be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ae0] =  Ifd35529b44c957737bf422127283c08e['h015c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ae1] =  Ifd35529b44c957737bf422127283c08e['h015c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ae2] =  Ifd35529b44c957737bf422127283c08e['h015c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ae3] =  Ifd35529b44c957737bf422127283c08e['h015c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ae4] =  Ifd35529b44c957737bf422127283c08e['h015c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ae5] =  Ifd35529b44c957737bf422127283c08e['h015ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ae6] =  Ifd35529b44c957737bf422127283c08e['h015cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ae7] =  Ifd35529b44c957737bf422127283c08e['h015ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ae8] =  Ifd35529b44c957737bf422127283c08e['h015d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ae9] =  Ifd35529b44c957737bf422127283c08e['h015d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00aea] =  Ifd35529b44c957737bf422127283c08e['h015d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00aeb] =  Ifd35529b44c957737bf422127283c08e['h015d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00aec] =  Ifd35529b44c957737bf422127283c08e['h015d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00aed] =  Ifd35529b44c957737bf422127283c08e['h015da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00aee] =  Ifd35529b44c957737bf422127283c08e['h015dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00aef] =  Ifd35529b44c957737bf422127283c08e['h015de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00af0] =  Ifd35529b44c957737bf422127283c08e['h015e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00af1] =  Ifd35529b44c957737bf422127283c08e['h015e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00af2] =  Ifd35529b44c957737bf422127283c08e['h015e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00af3] =  Ifd35529b44c957737bf422127283c08e['h015e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00af4] =  Ifd35529b44c957737bf422127283c08e['h015e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00af5] =  Ifd35529b44c957737bf422127283c08e['h015ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00af6] =  Ifd35529b44c957737bf422127283c08e['h015ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00af7] =  Ifd35529b44c957737bf422127283c08e['h015ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00af8] =  Ifd35529b44c957737bf422127283c08e['h015f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00af9] =  Ifd35529b44c957737bf422127283c08e['h015f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00afa] =  Ifd35529b44c957737bf422127283c08e['h015f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00afb] =  Ifd35529b44c957737bf422127283c08e['h015f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00afc] =  Ifd35529b44c957737bf422127283c08e['h015f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00afd] =  Ifd35529b44c957737bf422127283c08e['h015fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00afe] =  Ifd35529b44c957737bf422127283c08e['h015fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00aff] =  Ifd35529b44c957737bf422127283c08e['h015fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b00] =  Ifd35529b44c957737bf422127283c08e['h01600] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b01] =  Ifd35529b44c957737bf422127283c08e['h01602] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b02] =  Ifd35529b44c957737bf422127283c08e['h01604] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b03] =  Ifd35529b44c957737bf422127283c08e['h01606] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b04] =  Ifd35529b44c957737bf422127283c08e['h01608] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b05] =  Ifd35529b44c957737bf422127283c08e['h0160a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b06] =  Ifd35529b44c957737bf422127283c08e['h0160c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b07] =  Ifd35529b44c957737bf422127283c08e['h0160e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b08] =  Ifd35529b44c957737bf422127283c08e['h01610] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b09] =  Ifd35529b44c957737bf422127283c08e['h01612] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b0a] =  Ifd35529b44c957737bf422127283c08e['h01614] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b0b] =  Ifd35529b44c957737bf422127283c08e['h01616] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b0c] =  Ifd35529b44c957737bf422127283c08e['h01618] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b0d] =  Ifd35529b44c957737bf422127283c08e['h0161a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b0e] =  Ifd35529b44c957737bf422127283c08e['h0161c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b0f] =  Ifd35529b44c957737bf422127283c08e['h0161e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b10] =  Ifd35529b44c957737bf422127283c08e['h01620] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b11] =  Ifd35529b44c957737bf422127283c08e['h01622] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b12] =  Ifd35529b44c957737bf422127283c08e['h01624] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b13] =  Ifd35529b44c957737bf422127283c08e['h01626] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b14] =  Ifd35529b44c957737bf422127283c08e['h01628] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b15] =  Ifd35529b44c957737bf422127283c08e['h0162a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b16] =  Ifd35529b44c957737bf422127283c08e['h0162c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b17] =  Ifd35529b44c957737bf422127283c08e['h0162e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b18] =  Ifd35529b44c957737bf422127283c08e['h01630] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b19] =  Ifd35529b44c957737bf422127283c08e['h01632] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b1a] =  Ifd35529b44c957737bf422127283c08e['h01634] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b1b] =  Ifd35529b44c957737bf422127283c08e['h01636] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b1c] =  Ifd35529b44c957737bf422127283c08e['h01638] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b1d] =  Ifd35529b44c957737bf422127283c08e['h0163a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b1e] =  Ifd35529b44c957737bf422127283c08e['h0163c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b1f] =  Ifd35529b44c957737bf422127283c08e['h0163e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b20] =  Ifd35529b44c957737bf422127283c08e['h01640] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b21] =  Ifd35529b44c957737bf422127283c08e['h01642] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b22] =  Ifd35529b44c957737bf422127283c08e['h01644] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b23] =  Ifd35529b44c957737bf422127283c08e['h01646] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b24] =  Ifd35529b44c957737bf422127283c08e['h01648] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b25] =  Ifd35529b44c957737bf422127283c08e['h0164a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b26] =  Ifd35529b44c957737bf422127283c08e['h0164c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b27] =  Ifd35529b44c957737bf422127283c08e['h0164e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b28] =  Ifd35529b44c957737bf422127283c08e['h01650] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b29] =  Ifd35529b44c957737bf422127283c08e['h01652] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b2a] =  Ifd35529b44c957737bf422127283c08e['h01654] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b2b] =  Ifd35529b44c957737bf422127283c08e['h01656] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b2c] =  Ifd35529b44c957737bf422127283c08e['h01658] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b2d] =  Ifd35529b44c957737bf422127283c08e['h0165a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b2e] =  Ifd35529b44c957737bf422127283c08e['h0165c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b2f] =  Ifd35529b44c957737bf422127283c08e['h0165e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b30] =  Ifd35529b44c957737bf422127283c08e['h01660] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b31] =  Ifd35529b44c957737bf422127283c08e['h01662] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b32] =  Ifd35529b44c957737bf422127283c08e['h01664] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b33] =  Ifd35529b44c957737bf422127283c08e['h01666] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b34] =  Ifd35529b44c957737bf422127283c08e['h01668] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b35] =  Ifd35529b44c957737bf422127283c08e['h0166a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b36] =  Ifd35529b44c957737bf422127283c08e['h0166c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b37] =  Ifd35529b44c957737bf422127283c08e['h0166e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b38] =  Ifd35529b44c957737bf422127283c08e['h01670] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b39] =  Ifd35529b44c957737bf422127283c08e['h01672] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b3a] =  Ifd35529b44c957737bf422127283c08e['h01674] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b3b] =  Ifd35529b44c957737bf422127283c08e['h01676] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b3c] =  Ifd35529b44c957737bf422127283c08e['h01678] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b3d] =  Ifd35529b44c957737bf422127283c08e['h0167a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b3e] =  Ifd35529b44c957737bf422127283c08e['h0167c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b3f] =  Ifd35529b44c957737bf422127283c08e['h0167e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b40] =  Ifd35529b44c957737bf422127283c08e['h01680] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b41] =  Ifd35529b44c957737bf422127283c08e['h01682] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b42] =  Ifd35529b44c957737bf422127283c08e['h01684] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b43] =  Ifd35529b44c957737bf422127283c08e['h01686] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b44] =  Ifd35529b44c957737bf422127283c08e['h01688] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b45] =  Ifd35529b44c957737bf422127283c08e['h0168a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b46] =  Ifd35529b44c957737bf422127283c08e['h0168c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b47] =  Ifd35529b44c957737bf422127283c08e['h0168e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b48] =  Ifd35529b44c957737bf422127283c08e['h01690] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b49] =  Ifd35529b44c957737bf422127283c08e['h01692] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b4a] =  Ifd35529b44c957737bf422127283c08e['h01694] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b4b] =  Ifd35529b44c957737bf422127283c08e['h01696] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b4c] =  Ifd35529b44c957737bf422127283c08e['h01698] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b4d] =  Ifd35529b44c957737bf422127283c08e['h0169a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b4e] =  Ifd35529b44c957737bf422127283c08e['h0169c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b4f] =  Ifd35529b44c957737bf422127283c08e['h0169e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b50] =  Ifd35529b44c957737bf422127283c08e['h016a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b51] =  Ifd35529b44c957737bf422127283c08e['h016a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b52] =  Ifd35529b44c957737bf422127283c08e['h016a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b53] =  Ifd35529b44c957737bf422127283c08e['h016a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b54] =  Ifd35529b44c957737bf422127283c08e['h016a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b55] =  Ifd35529b44c957737bf422127283c08e['h016aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b56] =  Ifd35529b44c957737bf422127283c08e['h016ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b57] =  Ifd35529b44c957737bf422127283c08e['h016ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b58] =  Ifd35529b44c957737bf422127283c08e['h016b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b59] =  Ifd35529b44c957737bf422127283c08e['h016b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b5a] =  Ifd35529b44c957737bf422127283c08e['h016b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b5b] =  Ifd35529b44c957737bf422127283c08e['h016b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b5c] =  Ifd35529b44c957737bf422127283c08e['h016b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b5d] =  Ifd35529b44c957737bf422127283c08e['h016ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b5e] =  Ifd35529b44c957737bf422127283c08e['h016bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b5f] =  Ifd35529b44c957737bf422127283c08e['h016be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b60] =  Ifd35529b44c957737bf422127283c08e['h016c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b61] =  Ifd35529b44c957737bf422127283c08e['h016c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b62] =  Ifd35529b44c957737bf422127283c08e['h016c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b63] =  Ifd35529b44c957737bf422127283c08e['h016c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b64] =  Ifd35529b44c957737bf422127283c08e['h016c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b65] =  Ifd35529b44c957737bf422127283c08e['h016ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b66] =  Ifd35529b44c957737bf422127283c08e['h016cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b67] =  Ifd35529b44c957737bf422127283c08e['h016ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b68] =  Ifd35529b44c957737bf422127283c08e['h016d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b69] =  Ifd35529b44c957737bf422127283c08e['h016d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b6a] =  Ifd35529b44c957737bf422127283c08e['h016d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b6b] =  Ifd35529b44c957737bf422127283c08e['h016d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b6c] =  Ifd35529b44c957737bf422127283c08e['h016d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b6d] =  Ifd35529b44c957737bf422127283c08e['h016da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b6e] =  Ifd35529b44c957737bf422127283c08e['h016dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b6f] =  Ifd35529b44c957737bf422127283c08e['h016de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b70] =  Ifd35529b44c957737bf422127283c08e['h016e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b71] =  Ifd35529b44c957737bf422127283c08e['h016e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b72] =  Ifd35529b44c957737bf422127283c08e['h016e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b73] =  Ifd35529b44c957737bf422127283c08e['h016e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b74] =  Ifd35529b44c957737bf422127283c08e['h016e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b75] =  Ifd35529b44c957737bf422127283c08e['h016ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b76] =  Ifd35529b44c957737bf422127283c08e['h016ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b77] =  Ifd35529b44c957737bf422127283c08e['h016ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b78] =  Ifd35529b44c957737bf422127283c08e['h016f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b79] =  Ifd35529b44c957737bf422127283c08e['h016f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b7a] =  Ifd35529b44c957737bf422127283c08e['h016f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b7b] =  Ifd35529b44c957737bf422127283c08e['h016f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b7c] =  Ifd35529b44c957737bf422127283c08e['h016f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b7d] =  Ifd35529b44c957737bf422127283c08e['h016fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b7e] =  Ifd35529b44c957737bf422127283c08e['h016fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b7f] =  Ifd35529b44c957737bf422127283c08e['h016fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b80] =  Ifd35529b44c957737bf422127283c08e['h01700] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b81] =  Ifd35529b44c957737bf422127283c08e['h01702] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b82] =  Ifd35529b44c957737bf422127283c08e['h01704] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b83] =  Ifd35529b44c957737bf422127283c08e['h01706] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b84] =  Ifd35529b44c957737bf422127283c08e['h01708] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b85] =  Ifd35529b44c957737bf422127283c08e['h0170a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b86] =  Ifd35529b44c957737bf422127283c08e['h0170c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b87] =  Ifd35529b44c957737bf422127283c08e['h0170e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b88] =  Ifd35529b44c957737bf422127283c08e['h01710] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b89] =  Ifd35529b44c957737bf422127283c08e['h01712] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b8a] =  Ifd35529b44c957737bf422127283c08e['h01714] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b8b] =  Ifd35529b44c957737bf422127283c08e['h01716] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b8c] =  Ifd35529b44c957737bf422127283c08e['h01718] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b8d] =  Ifd35529b44c957737bf422127283c08e['h0171a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b8e] =  Ifd35529b44c957737bf422127283c08e['h0171c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b8f] =  Ifd35529b44c957737bf422127283c08e['h0171e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b90] =  Ifd35529b44c957737bf422127283c08e['h01720] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b91] =  Ifd35529b44c957737bf422127283c08e['h01722] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b92] =  Ifd35529b44c957737bf422127283c08e['h01724] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b93] =  Ifd35529b44c957737bf422127283c08e['h01726] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b94] =  Ifd35529b44c957737bf422127283c08e['h01728] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b95] =  Ifd35529b44c957737bf422127283c08e['h0172a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b96] =  Ifd35529b44c957737bf422127283c08e['h0172c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b97] =  Ifd35529b44c957737bf422127283c08e['h0172e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b98] =  Ifd35529b44c957737bf422127283c08e['h01730] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b99] =  Ifd35529b44c957737bf422127283c08e['h01732] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b9a] =  Ifd35529b44c957737bf422127283c08e['h01734] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b9b] =  Ifd35529b44c957737bf422127283c08e['h01736] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b9c] =  Ifd35529b44c957737bf422127283c08e['h01738] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b9d] =  Ifd35529b44c957737bf422127283c08e['h0173a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b9e] =  Ifd35529b44c957737bf422127283c08e['h0173c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00b9f] =  Ifd35529b44c957737bf422127283c08e['h0173e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ba0] =  Ifd35529b44c957737bf422127283c08e['h01740] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ba1] =  Ifd35529b44c957737bf422127283c08e['h01742] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ba2] =  Ifd35529b44c957737bf422127283c08e['h01744] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ba3] =  Ifd35529b44c957737bf422127283c08e['h01746] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ba4] =  Ifd35529b44c957737bf422127283c08e['h01748] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ba5] =  Ifd35529b44c957737bf422127283c08e['h0174a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ba6] =  Ifd35529b44c957737bf422127283c08e['h0174c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ba7] =  Ifd35529b44c957737bf422127283c08e['h0174e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ba8] =  Ifd35529b44c957737bf422127283c08e['h01750] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ba9] =  Ifd35529b44c957737bf422127283c08e['h01752] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00baa] =  Ifd35529b44c957737bf422127283c08e['h01754] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bab] =  Ifd35529b44c957737bf422127283c08e['h01756] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bac] =  Ifd35529b44c957737bf422127283c08e['h01758] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bad] =  Ifd35529b44c957737bf422127283c08e['h0175a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bae] =  Ifd35529b44c957737bf422127283c08e['h0175c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00baf] =  Ifd35529b44c957737bf422127283c08e['h0175e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bb0] =  Ifd35529b44c957737bf422127283c08e['h01760] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bb1] =  Ifd35529b44c957737bf422127283c08e['h01762] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bb2] =  Ifd35529b44c957737bf422127283c08e['h01764] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bb3] =  Ifd35529b44c957737bf422127283c08e['h01766] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bb4] =  Ifd35529b44c957737bf422127283c08e['h01768] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bb5] =  Ifd35529b44c957737bf422127283c08e['h0176a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bb6] =  Ifd35529b44c957737bf422127283c08e['h0176c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bb7] =  Ifd35529b44c957737bf422127283c08e['h0176e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bb8] =  Ifd35529b44c957737bf422127283c08e['h01770] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bb9] =  Ifd35529b44c957737bf422127283c08e['h01772] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bba] =  Ifd35529b44c957737bf422127283c08e['h01774] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bbb] =  Ifd35529b44c957737bf422127283c08e['h01776] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bbc] =  Ifd35529b44c957737bf422127283c08e['h01778] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bbd] =  Ifd35529b44c957737bf422127283c08e['h0177a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bbe] =  Ifd35529b44c957737bf422127283c08e['h0177c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bbf] =  Ifd35529b44c957737bf422127283c08e['h0177e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bc0] =  Ifd35529b44c957737bf422127283c08e['h01780] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bc1] =  Ifd35529b44c957737bf422127283c08e['h01782] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bc2] =  Ifd35529b44c957737bf422127283c08e['h01784] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bc3] =  Ifd35529b44c957737bf422127283c08e['h01786] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bc4] =  Ifd35529b44c957737bf422127283c08e['h01788] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bc5] =  Ifd35529b44c957737bf422127283c08e['h0178a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bc6] =  Ifd35529b44c957737bf422127283c08e['h0178c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bc7] =  Ifd35529b44c957737bf422127283c08e['h0178e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bc8] =  Ifd35529b44c957737bf422127283c08e['h01790] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bc9] =  Ifd35529b44c957737bf422127283c08e['h01792] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bca] =  Ifd35529b44c957737bf422127283c08e['h01794] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bcb] =  Ifd35529b44c957737bf422127283c08e['h01796] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bcc] =  Ifd35529b44c957737bf422127283c08e['h01798] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bcd] =  Ifd35529b44c957737bf422127283c08e['h0179a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bce] =  Ifd35529b44c957737bf422127283c08e['h0179c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bcf] =  Ifd35529b44c957737bf422127283c08e['h0179e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bd0] =  Ifd35529b44c957737bf422127283c08e['h017a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bd1] =  Ifd35529b44c957737bf422127283c08e['h017a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bd2] =  Ifd35529b44c957737bf422127283c08e['h017a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bd3] =  Ifd35529b44c957737bf422127283c08e['h017a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bd4] =  Ifd35529b44c957737bf422127283c08e['h017a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bd5] =  Ifd35529b44c957737bf422127283c08e['h017aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bd6] =  Ifd35529b44c957737bf422127283c08e['h017ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bd7] =  Ifd35529b44c957737bf422127283c08e['h017ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bd8] =  Ifd35529b44c957737bf422127283c08e['h017b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bd9] =  Ifd35529b44c957737bf422127283c08e['h017b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bda] =  Ifd35529b44c957737bf422127283c08e['h017b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bdb] =  Ifd35529b44c957737bf422127283c08e['h017b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bdc] =  Ifd35529b44c957737bf422127283c08e['h017b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bdd] =  Ifd35529b44c957737bf422127283c08e['h017ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bde] =  Ifd35529b44c957737bf422127283c08e['h017bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bdf] =  Ifd35529b44c957737bf422127283c08e['h017be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00be0] =  Ifd35529b44c957737bf422127283c08e['h017c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00be1] =  Ifd35529b44c957737bf422127283c08e['h017c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00be2] =  Ifd35529b44c957737bf422127283c08e['h017c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00be3] =  Ifd35529b44c957737bf422127283c08e['h017c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00be4] =  Ifd35529b44c957737bf422127283c08e['h017c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00be5] =  Ifd35529b44c957737bf422127283c08e['h017ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00be6] =  Ifd35529b44c957737bf422127283c08e['h017cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00be7] =  Ifd35529b44c957737bf422127283c08e['h017ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00be8] =  Ifd35529b44c957737bf422127283c08e['h017d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00be9] =  Ifd35529b44c957737bf422127283c08e['h017d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bea] =  Ifd35529b44c957737bf422127283c08e['h017d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00beb] =  Ifd35529b44c957737bf422127283c08e['h017d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bec] =  Ifd35529b44c957737bf422127283c08e['h017d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bed] =  Ifd35529b44c957737bf422127283c08e['h017da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bee] =  Ifd35529b44c957737bf422127283c08e['h017dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bef] =  Ifd35529b44c957737bf422127283c08e['h017de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bf0] =  Ifd35529b44c957737bf422127283c08e['h017e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bf1] =  Ifd35529b44c957737bf422127283c08e['h017e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bf2] =  Ifd35529b44c957737bf422127283c08e['h017e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bf3] =  Ifd35529b44c957737bf422127283c08e['h017e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bf4] =  Ifd35529b44c957737bf422127283c08e['h017e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bf5] =  Ifd35529b44c957737bf422127283c08e['h017ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bf6] =  Ifd35529b44c957737bf422127283c08e['h017ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bf7] =  Ifd35529b44c957737bf422127283c08e['h017ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bf8] =  Ifd35529b44c957737bf422127283c08e['h017f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bf9] =  Ifd35529b44c957737bf422127283c08e['h017f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bfa] =  Ifd35529b44c957737bf422127283c08e['h017f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bfb] =  Ifd35529b44c957737bf422127283c08e['h017f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bfc] =  Ifd35529b44c957737bf422127283c08e['h017f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bfd] =  Ifd35529b44c957737bf422127283c08e['h017fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bfe] =  Ifd35529b44c957737bf422127283c08e['h017fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00bff] =  Ifd35529b44c957737bf422127283c08e['h017fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c00] =  Ifd35529b44c957737bf422127283c08e['h01800] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c01] =  Ifd35529b44c957737bf422127283c08e['h01802] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c02] =  Ifd35529b44c957737bf422127283c08e['h01804] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c03] =  Ifd35529b44c957737bf422127283c08e['h01806] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c04] =  Ifd35529b44c957737bf422127283c08e['h01808] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c05] =  Ifd35529b44c957737bf422127283c08e['h0180a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c06] =  Ifd35529b44c957737bf422127283c08e['h0180c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c07] =  Ifd35529b44c957737bf422127283c08e['h0180e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c08] =  Ifd35529b44c957737bf422127283c08e['h01810] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c09] =  Ifd35529b44c957737bf422127283c08e['h01812] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c0a] =  Ifd35529b44c957737bf422127283c08e['h01814] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c0b] =  Ifd35529b44c957737bf422127283c08e['h01816] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c0c] =  Ifd35529b44c957737bf422127283c08e['h01818] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c0d] =  Ifd35529b44c957737bf422127283c08e['h0181a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c0e] =  Ifd35529b44c957737bf422127283c08e['h0181c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c0f] =  Ifd35529b44c957737bf422127283c08e['h0181e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c10] =  Ifd35529b44c957737bf422127283c08e['h01820] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c11] =  Ifd35529b44c957737bf422127283c08e['h01822] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c12] =  Ifd35529b44c957737bf422127283c08e['h01824] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c13] =  Ifd35529b44c957737bf422127283c08e['h01826] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c14] =  Ifd35529b44c957737bf422127283c08e['h01828] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c15] =  Ifd35529b44c957737bf422127283c08e['h0182a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c16] =  Ifd35529b44c957737bf422127283c08e['h0182c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c17] =  Ifd35529b44c957737bf422127283c08e['h0182e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c18] =  Ifd35529b44c957737bf422127283c08e['h01830] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c19] =  Ifd35529b44c957737bf422127283c08e['h01832] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c1a] =  Ifd35529b44c957737bf422127283c08e['h01834] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c1b] =  Ifd35529b44c957737bf422127283c08e['h01836] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c1c] =  Ifd35529b44c957737bf422127283c08e['h01838] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c1d] =  Ifd35529b44c957737bf422127283c08e['h0183a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c1e] =  Ifd35529b44c957737bf422127283c08e['h0183c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c1f] =  Ifd35529b44c957737bf422127283c08e['h0183e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c20] =  Ifd35529b44c957737bf422127283c08e['h01840] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c21] =  Ifd35529b44c957737bf422127283c08e['h01842] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c22] =  Ifd35529b44c957737bf422127283c08e['h01844] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c23] =  Ifd35529b44c957737bf422127283c08e['h01846] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c24] =  Ifd35529b44c957737bf422127283c08e['h01848] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c25] =  Ifd35529b44c957737bf422127283c08e['h0184a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c26] =  Ifd35529b44c957737bf422127283c08e['h0184c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c27] =  Ifd35529b44c957737bf422127283c08e['h0184e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c28] =  Ifd35529b44c957737bf422127283c08e['h01850] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c29] =  Ifd35529b44c957737bf422127283c08e['h01852] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c2a] =  Ifd35529b44c957737bf422127283c08e['h01854] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c2b] =  Ifd35529b44c957737bf422127283c08e['h01856] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c2c] =  Ifd35529b44c957737bf422127283c08e['h01858] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c2d] =  Ifd35529b44c957737bf422127283c08e['h0185a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c2e] =  Ifd35529b44c957737bf422127283c08e['h0185c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c2f] =  Ifd35529b44c957737bf422127283c08e['h0185e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c30] =  Ifd35529b44c957737bf422127283c08e['h01860] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c31] =  Ifd35529b44c957737bf422127283c08e['h01862] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c32] =  Ifd35529b44c957737bf422127283c08e['h01864] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c33] =  Ifd35529b44c957737bf422127283c08e['h01866] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c34] =  Ifd35529b44c957737bf422127283c08e['h01868] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c35] =  Ifd35529b44c957737bf422127283c08e['h0186a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c36] =  Ifd35529b44c957737bf422127283c08e['h0186c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c37] =  Ifd35529b44c957737bf422127283c08e['h0186e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c38] =  Ifd35529b44c957737bf422127283c08e['h01870] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c39] =  Ifd35529b44c957737bf422127283c08e['h01872] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c3a] =  Ifd35529b44c957737bf422127283c08e['h01874] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c3b] =  Ifd35529b44c957737bf422127283c08e['h01876] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c3c] =  Ifd35529b44c957737bf422127283c08e['h01878] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c3d] =  Ifd35529b44c957737bf422127283c08e['h0187a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c3e] =  Ifd35529b44c957737bf422127283c08e['h0187c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c3f] =  Ifd35529b44c957737bf422127283c08e['h0187e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c40] =  Ifd35529b44c957737bf422127283c08e['h01880] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c41] =  Ifd35529b44c957737bf422127283c08e['h01882] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c42] =  Ifd35529b44c957737bf422127283c08e['h01884] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c43] =  Ifd35529b44c957737bf422127283c08e['h01886] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c44] =  Ifd35529b44c957737bf422127283c08e['h01888] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c45] =  Ifd35529b44c957737bf422127283c08e['h0188a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c46] =  Ifd35529b44c957737bf422127283c08e['h0188c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c47] =  Ifd35529b44c957737bf422127283c08e['h0188e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c48] =  Ifd35529b44c957737bf422127283c08e['h01890] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c49] =  Ifd35529b44c957737bf422127283c08e['h01892] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c4a] =  Ifd35529b44c957737bf422127283c08e['h01894] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c4b] =  Ifd35529b44c957737bf422127283c08e['h01896] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c4c] =  Ifd35529b44c957737bf422127283c08e['h01898] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c4d] =  Ifd35529b44c957737bf422127283c08e['h0189a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c4e] =  Ifd35529b44c957737bf422127283c08e['h0189c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c4f] =  Ifd35529b44c957737bf422127283c08e['h0189e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c50] =  Ifd35529b44c957737bf422127283c08e['h018a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c51] =  Ifd35529b44c957737bf422127283c08e['h018a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c52] =  Ifd35529b44c957737bf422127283c08e['h018a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c53] =  Ifd35529b44c957737bf422127283c08e['h018a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c54] =  Ifd35529b44c957737bf422127283c08e['h018a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c55] =  Ifd35529b44c957737bf422127283c08e['h018aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c56] =  Ifd35529b44c957737bf422127283c08e['h018ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c57] =  Ifd35529b44c957737bf422127283c08e['h018ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c58] =  Ifd35529b44c957737bf422127283c08e['h018b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c59] =  Ifd35529b44c957737bf422127283c08e['h018b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c5a] =  Ifd35529b44c957737bf422127283c08e['h018b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c5b] =  Ifd35529b44c957737bf422127283c08e['h018b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c5c] =  Ifd35529b44c957737bf422127283c08e['h018b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c5d] =  Ifd35529b44c957737bf422127283c08e['h018ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c5e] =  Ifd35529b44c957737bf422127283c08e['h018bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c5f] =  Ifd35529b44c957737bf422127283c08e['h018be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c60] =  Ifd35529b44c957737bf422127283c08e['h018c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c61] =  Ifd35529b44c957737bf422127283c08e['h018c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c62] =  Ifd35529b44c957737bf422127283c08e['h018c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c63] =  Ifd35529b44c957737bf422127283c08e['h018c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c64] =  Ifd35529b44c957737bf422127283c08e['h018c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c65] =  Ifd35529b44c957737bf422127283c08e['h018ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c66] =  Ifd35529b44c957737bf422127283c08e['h018cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c67] =  Ifd35529b44c957737bf422127283c08e['h018ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c68] =  Ifd35529b44c957737bf422127283c08e['h018d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c69] =  Ifd35529b44c957737bf422127283c08e['h018d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c6a] =  Ifd35529b44c957737bf422127283c08e['h018d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c6b] =  Ifd35529b44c957737bf422127283c08e['h018d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c6c] =  Ifd35529b44c957737bf422127283c08e['h018d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c6d] =  Ifd35529b44c957737bf422127283c08e['h018da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c6e] =  Ifd35529b44c957737bf422127283c08e['h018dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c6f] =  Ifd35529b44c957737bf422127283c08e['h018de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c70] =  Ifd35529b44c957737bf422127283c08e['h018e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c71] =  Ifd35529b44c957737bf422127283c08e['h018e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c72] =  Ifd35529b44c957737bf422127283c08e['h018e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c73] =  Ifd35529b44c957737bf422127283c08e['h018e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c74] =  Ifd35529b44c957737bf422127283c08e['h018e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c75] =  Ifd35529b44c957737bf422127283c08e['h018ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c76] =  Ifd35529b44c957737bf422127283c08e['h018ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c77] =  Ifd35529b44c957737bf422127283c08e['h018ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c78] =  Ifd35529b44c957737bf422127283c08e['h018f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c79] =  Ifd35529b44c957737bf422127283c08e['h018f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c7a] =  Ifd35529b44c957737bf422127283c08e['h018f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c7b] =  Ifd35529b44c957737bf422127283c08e['h018f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c7c] =  Ifd35529b44c957737bf422127283c08e['h018f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c7d] =  Ifd35529b44c957737bf422127283c08e['h018fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c7e] =  Ifd35529b44c957737bf422127283c08e['h018fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c7f] =  Ifd35529b44c957737bf422127283c08e['h018fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c80] =  Ifd35529b44c957737bf422127283c08e['h01900] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c81] =  Ifd35529b44c957737bf422127283c08e['h01902] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c82] =  Ifd35529b44c957737bf422127283c08e['h01904] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c83] =  Ifd35529b44c957737bf422127283c08e['h01906] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c84] =  Ifd35529b44c957737bf422127283c08e['h01908] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c85] =  Ifd35529b44c957737bf422127283c08e['h0190a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c86] =  Ifd35529b44c957737bf422127283c08e['h0190c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c87] =  Ifd35529b44c957737bf422127283c08e['h0190e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c88] =  Ifd35529b44c957737bf422127283c08e['h01910] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c89] =  Ifd35529b44c957737bf422127283c08e['h01912] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c8a] =  Ifd35529b44c957737bf422127283c08e['h01914] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c8b] =  Ifd35529b44c957737bf422127283c08e['h01916] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c8c] =  Ifd35529b44c957737bf422127283c08e['h01918] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c8d] =  Ifd35529b44c957737bf422127283c08e['h0191a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c8e] =  Ifd35529b44c957737bf422127283c08e['h0191c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c8f] =  Ifd35529b44c957737bf422127283c08e['h0191e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c90] =  Ifd35529b44c957737bf422127283c08e['h01920] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c91] =  Ifd35529b44c957737bf422127283c08e['h01922] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c92] =  Ifd35529b44c957737bf422127283c08e['h01924] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c93] =  Ifd35529b44c957737bf422127283c08e['h01926] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c94] =  Ifd35529b44c957737bf422127283c08e['h01928] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c95] =  Ifd35529b44c957737bf422127283c08e['h0192a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c96] =  Ifd35529b44c957737bf422127283c08e['h0192c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c97] =  Ifd35529b44c957737bf422127283c08e['h0192e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c98] =  Ifd35529b44c957737bf422127283c08e['h01930] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c99] =  Ifd35529b44c957737bf422127283c08e['h01932] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c9a] =  Ifd35529b44c957737bf422127283c08e['h01934] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c9b] =  Ifd35529b44c957737bf422127283c08e['h01936] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c9c] =  Ifd35529b44c957737bf422127283c08e['h01938] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c9d] =  Ifd35529b44c957737bf422127283c08e['h0193a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c9e] =  Ifd35529b44c957737bf422127283c08e['h0193c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00c9f] =  Ifd35529b44c957737bf422127283c08e['h0193e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ca0] =  Ifd35529b44c957737bf422127283c08e['h01940] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ca1] =  Ifd35529b44c957737bf422127283c08e['h01942] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ca2] =  Ifd35529b44c957737bf422127283c08e['h01944] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ca3] =  Ifd35529b44c957737bf422127283c08e['h01946] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ca4] =  Ifd35529b44c957737bf422127283c08e['h01948] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ca5] =  Ifd35529b44c957737bf422127283c08e['h0194a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ca6] =  Ifd35529b44c957737bf422127283c08e['h0194c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ca7] =  Ifd35529b44c957737bf422127283c08e['h0194e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ca8] =  Ifd35529b44c957737bf422127283c08e['h01950] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ca9] =  Ifd35529b44c957737bf422127283c08e['h01952] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00caa] =  Ifd35529b44c957737bf422127283c08e['h01954] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cab] =  Ifd35529b44c957737bf422127283c08e['h01956] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cac] =  Ifd35529b44c957737bf422127283c08e['h01958] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cad] =  Ifd35529b44c957737bf422127283c08e['h0195a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cae] =  Ifd35529b44c957737bf422127283c08e['h0195c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00caf] =  Ifd35529b44c957737bf422127283c08e['h0195e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cb0] =  Ifd35529b44c957737bf422127283c08e['h01960] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cb1] =  Ifd35529b44c957737bf422127283c08e['h01962] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cb2] =  Ifd35529b44c957737bf422127283c08e['h01964] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cb3] =  Ifd35529b44c957737bf422127283c08e['h01966] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cb4] =  Ifd35529b44c957737bf422127283c08e['h01968] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cb5] =  Ifd35529b44c957737bf422127283c08e['h0196a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cb6] =  Ifd35529b44c957737bf422127283c08e['h0196c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cb7] =  Ifd35529b44c957737bf422127283c08e['h0196e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cb8] =  Ifd35529b44c957737bf422127283c08e['h01970] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cb9] =  Ifd35529b44c957737bf422127283c08e['h01972] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cba] =  Ifd35529b44c957737bf422127283c08e['h01974] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cbb] =  Ifd35529b44c957737bf422127283c08e['h01976] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cbc] =  Ifd35529b44c957737bf422127283c08e['h01978] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cbd] =  Ifd35529b44c957737bf422127283c08e['h0197a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cbe] =  Ifd35529b44c957737bf422127283c08e['h0197c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cbf] =  Ifd35529b44c957737bf422127283c08e['h0197e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cc0] =  Ifd35529b44c957737bf422127283c08e['h01980] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cc1] =  Ifd35529b44c957737bf422127283c08e['h01982] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cc2] =  Ifd35529b44c957737bf422127283c08e['h01984] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cc3] =  Ifd35529b44c957737bf422127283c08e['h01986] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cc4] =  Ifd35529b44c957737bf422127283c08e['h01988] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cc5] =  Ifd35529b44c957737bf422127283c08e['h0198a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cc6] =  Ifd35529b44c957737bf422127283c08e['h0198c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cc7] =  Ifd35529b44c957737bf422127283c08e['h0198e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cc8] =  Ifd35529b44c957737bf422127283c08e['h01990] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cc9] =  Ifd35529b44c957737bf422127283c08e['h01992] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cca] =  Ifd35529b44c957737bf422127283c08e['h01994] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ccb] =  Ifd35529b44c957737bf422127283c08e['h01996] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ccc] =  Ifd35529b44c957737bf422127283c08e['h01998] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ccd] =  Ifd35529b44c957737bf422127283c08e['h0199a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cce] =  Ifd35529b44c957737bf422127283c08e['h0199c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ccf] =  Ifd35529b44c957737bf422127283c08e['h0199e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cd0] =  Ifd35529b44c957737bf422127283c08e['h019a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cd1] =  Ifd35529b44c957737bf422127283c08e['h019a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cd2] =  Ifd35529b44c957737bf422127283c08e['h019a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cd3] =  Ifd35529b44c957737bf422127283c08e['h019a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cd4] =  Ifd35529b44c957737bf422127283c08e['h019a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cd5] =  Ifd35529b44c957737bf422127283c08e['h019aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cd6] =  Ifd35529b44c957737bf422127283c08e['h019ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cd7] =  Ifd35529b44c957737bf422127283c08e['h019ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cd8] =  Ifd35529b44c957737bf422127283c08e['h019b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cd9] =  Ifd35529b44c957737bf422127283c08e['h019b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cda] =  Ifd35529b44c957737bf422127283c08e['h019b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cdb] =  Ifd35529b44c957737bf422127283c08e['h019b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cdc] =  Ifd35529b44c957737bf422127283c08e['h019b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cdd] =  Ifd35529b44c957737bf422127283c08e['h019ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cde] =  Ifd35529b44c957737bf422127283c08e['h019bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cdf] =  Ifd35529b44c957737bf422127283c08e['h019be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ce0] =  Ifd35529b44c957737bf422127283c08e['h019c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ce1] =  Ifd35529b44c957737bf422127283c08e['h019c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ce2] =  Ifd35529b44c957737bf422127283c08e['h019c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ce3] =  Ifd35529b44c957737bf422127283c08e['h019c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ce4] =  Ifd35529b44c957737bf422127283c08e['h019c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ce5] =  Ifd35529b44c957737bf422127283c08e['h019ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ce6] =  Ifd35529b44c957737bf422127283c08e['h019cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ce7] =  Ifd35529b44c957737bf422127283c08e['h019ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ce8] =  Ifd35529b44c957737bf422127283c08e['h019d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ce9] =  Ifd35529b44c957737bf422127283c08e['h019d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cea] =  Ifd35529b44c957737bf422127283c08e['h019d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ceb] =  Ifd35529b44c957737bf422127283c08e['h019d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cec] =  Ifd35529b44c957737bf422127283c08e['h019d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ced] =  Ifd35529b44c957737bf422127283c08e['h019da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cee] =  Ifd35529b44c957737bf422127283c08e['h019dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cef] =  Ifd35529b44c957737bf422127283c08e['h019de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cf0] =  Ifd35529b44c957737bf422127283c08e['h019e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cf1] =  Ifd35529b44c957737bf422127283c08e['h019e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cf2] =  Ifd35529b44c957737bf422127283c08e['h019e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cf3] =  Ifd35529b44c957737bf422127283c08e['h019e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cf4] =  Ifd35529b44c957737bf422127283c08e['h019e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cf5] =  Ifd35529b44c957737bf422127283c08e['h019ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cf6] =  Ifd35529b44c957737bf422127283c08e['h019ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cf7] =  Ifd35529b44c957737bf422127283c08e['h019ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cf8] =  Ifd35529b44c957737bf422127283c08e['h019f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cf9] =  Ifd35529b44c957737bf422127283c08e['h019f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cfa] =  Ifd35529b44c957737bf422127283c08e['h019f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cfb] =  Ifd35529b44c957737bf422127283c08e['h019f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cfc] =  Ifd35529b44c957737bf422127283c08e['h019f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cfd] =  Ifd35529b44c957737bf422127283c08e['h019fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cfe] =  Ifd35529b44c957737bf422127283c08e['h019fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00cff] =  Ifd35529b44c957737bf422127283c08e['h019fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d00] =  Ifd35529b44c957737bf422127283c08e['h01a00] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d01] =  Ifd35529b44c957737bf422127283c08e['h01a02] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d02] =  Ifd35529b44c957737bf422127283c08e['h01a04] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d03] =  Ifd35529b44c957737bf422127283c08e['h01a06] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d04] =  Ifd35529b44c957737bf422127283c08e['h01a08] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d05] =  Ifd35529b44c957737bf422127283c08e['h01a0a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d06] =  Ifd35529b44c957737bf422127283c08e['h01a0c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d07] =  Ifd35529b44c957737bf422127283c08e['h01a0e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d08] =  Ifd35529b44c957737bf422127283c08e['h01a10] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d09] =  Ifd35529b44c957737bf422127283c08e['h01a12] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d0a] =  Ifd35529b44c957737bf422127283c08e['h01a14] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d0b] =  Ifd35529b44c957737bf422127283c08e['h01a16] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d0c] =  Ifd35529b44c957737bf422127283c08e['h01a18] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d0d] =  Ifd35529b44c957737bf422127283c08e['h01a1a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d0e] =  Ifd35529b44c957737bf422127283c08e['h01a1c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d0f] =  Ifd35529b44c957737bf422127283c08e['h01a1e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d10] =  Ifd35529b44c957737bf422127283c08e['h01a20] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d11] =  Ifd35529b44c957737bf422127283c08e['h01a22] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d12] =  Ifd35529b44c957737bf422127283c08e['h01a24] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d13] =  Ifd35529b44c957737bf422127283c08e['h01a26] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d14] =  Ifd35529b44c957737bf422127283c08e['h01a28] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d15] =  Ifd35529b44c957737bf422127283c08e['h01a2a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d16] =  Ifd35529b44c957737bf422127283c08e['h01a2c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d17] =  Ifd35529b44c957737bf422127283c08e['h01a2e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d18] =  Ifd35529b44c957737bf422127283c08e['h01a30] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d19] =  Ifd35529b44c957737bf422127283c08e['h01a32] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d1a] =  Ifd35529b44c957737bf422127283c08e['h01a34] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d1b] =  Ifd35529b44c957737bf422127283c08e['h01a36] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d1c] =  Ifd35529b44c957737bf422127283c08e['h01a38] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d1d] =  Ifd35529b44c957737bf422127283c08e['h01a3a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d1e] =  Ifd35529b44c957737bf422127283c08e['h01a3c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d1f] =  Ifd35529b44c957737bf422127283c08e['h01a3e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d20] =  Ifd35529b44c957737bf422127283c08e['h01a40] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d21] =  Ifd35529b44c957737bf422127283c08e['h01a42] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d22] =  Ifd35529b44c957737bf422127283c08e['h01a44] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d23] =  Ifd35529b44c957737bf422127283c08e['h01a46] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d24] =  Ifd35529b44c957737bf422127283c08e['h01a48] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d25] =  Ifd35529b44c957737bf422127283c08e['h01a4a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d26] =  Ifd35529b44c957737bf422127283c08e['h01a4c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d27] =  Ifd35529b44c957737bf422127283c08e['h01a4e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d28] =  Ifd35529b44c957737bf422127283c08e['h01a50] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d29] =  Ifd35529b44c957737bf422127283c08e['h01a52] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d2a] =  Ifd35529b44c957737bf422127283c08e['h01a54] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d2b] =  Ifd35529b44c957737bf422127283c08e['h01a56] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d2c] =  Ifd35529b44c957737bf422127283c08e['h01a58] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d2d] =  Ifd35529b44c957737bf422127283c08e['h01a5a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d2e] =  Ifd35529b44c957737bf422127283c08e['h01a5c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d2f] =  Ifd35529b44c957737bf422127283c08e['h01a5e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d30] =  Ifd35529b44c957737bf422127283c08e['h01a60] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d31] =  Ifd35529b44c957737bf422127283c08e['h01a62] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d32] =  Ifd35529b44c957737bf422127283c08e['h01a64] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d33] =  Ifd35529b44c957737bf422127283c08e['h01a66] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d34] =  Ifd35529b44c957737bf422127283c08e['h01a68] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d35] =  Ifd35529b44c957737bf422127283c08e['h01a6a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d36] =  Ifd35529b44c957737bf422127283c08e['h01a6c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d37] =  Ifd35529b44c957737bf422127283c08e['h01a6e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d38] =  Ifd35529b44c957737bf422127283c08e['h01a70] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d39] =  Ifd35529b44c957737bf422127283c08e['h01a72] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d3a] =  Ifd35529b44c957737bf422127283c08e['h01a74] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d3b] =  Ifd35529b44c957737bf422127283c08e['h01a76] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d3c] =  Ifd35529b44c957737bf422127283c08e['h01a78] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d3d] =  Ifd35529b44c957737bf422127283c08e['h01a7a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d3e] =  Ifd35529b44c957737bf422127283c08e['h01a7c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d3f] =  Ifd35529b44c957737bf422127283c08e['h01a7e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d40] =  Ifd35529b44c957737bf422127283c08e['h01a80] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d41] =  Ifd35529b44c957737bf422127283c08e['h01a82] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d42] =  Ifd35529b44c957737bf422127283c08e['h01a84] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d43] =  Ifd35529b44c957737bf422127283c08e['h01a86] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d44] =  Ifd35529b44c957737bf422127283c08e['h01a88] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d45] =  Ifd35529b44c957737bf422127283c08e['h01a8a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d46] =  Ifd35529b44c957737bf422127283c08e['h01a8c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d47] =  Ifd35529b44c957737bf422127283c08e['h01a8e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d48] =  Ifd35529b44c957737bf422127283c08e['h01a90] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d49] =  Ifd35529b44c957737bf422127283c08e['h01a92] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d4a] =  Ifd35529b44c957737bf422127283c08e['h01a94] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d4b] =  Ifd35529b44c957737bf422127283c08e['h01a96] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d4c] =  Ifd35529b44c957737bf422127283c08e['h01a98] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d4d] =  Ifd35529b44c957737bf422127283c08e['h01a9a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d4e] =  Ifd35529b44c957737bf422127283c08e['h01a9c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d4f] =  Ifd35529b44c957737bf422127283c08e['h01a9e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d50] =  Ifd35529b44c957737bf422127283c08e['h01aa0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d51] =  Ifd35529b44c957737bf422127283c08e['h01aa2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d52] =  Ifd35529b44c957737bf422127283c08e['h01aa4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d53] =  Ifd35529b44c957737bf422127283c08e['h01aa6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d54] =  Ifd35529b44c957737bf422127283c08e['h01aa8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d55] =  Ifd35529b44c957737bf422127283c08e['h01aaa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d56] =  Ifd35529b44c957737bf422127283c08e['h01aac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d57] =  Ifd35529b44c957737bf422127283c08e['h01aae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d58] =  Ifd35529b44c957737bf422127283c08e['h01ab0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d59] =  Ifd35529b44c957737bf422127283c08e['h01ab2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d5a] =  Ifd35529b44c957737bf422127283c08e['h01ab4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d5b] =  Ifd35529b44c957737bf422127283c08e['h01ab6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d5c] =  Ifd35529b44c957737bf422127283c08e['h01ab8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d5d] =  Ifd35529b44c957737bf422127283c08e['h01aba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d5e] =  Ifd35529b44c957737bf422127283c08e['h01abc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d5f] =  Ifd35529b44c957737bf422127283c08e['h01abe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d60] =  Ifd35529b44c957737bf422127283c08e['h01ac0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d61] =  Ifd35529b44c957737bf422127283c08e['h01ac2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d62] =  Ifd35529b44c957737bf422127283c08e['h01ac4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d63] =  Ifd35529b44c957737bf422127283c08e['h01ac6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d64] =  Ifd35529b44c957737bf422127283c08e['h01ac8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d65] =  Ifd35529b44c957737bf422127283c08e['h01aca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d66] =  Ifd35529b44c957737bf422127283c08e['h01acc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d67] =  Ifd35529b44c957737bf422127283c08e['h01ace] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d68] =  Ifd35529b44c957737bf422127283c08e['h01ad0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d69] =  Ifd35529b44c957737bf422127283c08e['h01ad2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d6a] =  Ifd35529b44c957737bf422127283c08e['h01ad4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d6b] =  Ifd35529b44c957737bf422127283c08e['h01ad6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d6c] =  Ifd35529b44c957737bf422127283c08e['h01ad8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d6d] =  Ifd35529b44c957737bf422127283c08e['h01ada] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d6e] =  Ifd35529b44c957737bf422127283c08e['h01adc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d6f] =  Ifd35529b44c957737bf422127283c08e['h01ade] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d70] =  Ifd35529b44c957737bf422127283c08e['h01ae0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d71] =  Ifd35529b44c957737bf422127283c08e['h01ae2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d72] =  Ifd35529b44c957737bf422127283c08e['h01ae4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d73] =  Ifd35529b44c957737bf422127283c08e['h01ae6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d74] =  Ifd35529b44c957737bf422127283c08e['h01ae8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d75] =  Ifd35529b44c957737bf422127283c08e['h01aea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d76] =  Ifd35529b44c957737bf422127283c08e['h01aec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d77] =  Ifd35529b44c957737bf422127283c08e['h01aee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d78] =  Ifd35529b44c957737bf422127283c08e['h01af0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d79] =  Ifd35529b44c957737bf422127283c08e['h01af2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d7a] =  Ifd35529b44c957737bf422127283c08e['h01af4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d7b] =  Ifd35529b44c957737bf422127283c08e['h01af6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d7c] =  Ifd35529b44c957737bf422127283c08e['h01af8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d7d] =  Ifd35529b44c957737bf422127283c08e['h01afa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d7e] =  Ifd35529b44c957737bf422127283c08e['h01afc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d7f] =  Ifd35529b44c957737bf422127283c08e['h01afe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d80] =  Ifd35529b44c957737bf422127283c08e['h01b00] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d81] =  Ifd35529b44c957737bf422127283c08e['h01b02] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d82] =  Ifd35529b44c957737bf422127283c08e['h01b04] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d83] =  Ifd35529b44c957737bf422127283c08e['h01b06] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d84] =  Ifd35529b44c957737bf422127283c08e['h01b08] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d85] =  Ifd35529b44c957737bf422127283c08e['h01b0a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d86] =  Ifd35529b44c957737bf422127283c08e['h01b0c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d87] =  Ifd35529b44c957737bf422127283c08e['h01b0e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d88] =  Ifd35529b44c957737bf422127283c08e['h01b10] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d89] =  Ifd35529b44c957737bf422127283c08e['h01b12] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d8a] =  Ifd35529b44c957737bf422127283c08e['h01b14] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d8b] =  Ifd35529b44c957737bf422127283c08e['h01b16] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d8c] =  Ifd35529b44c957737bf422127283c08e['h01b18] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d8d] =  Ifd35529b44c957737bf422127283c08e['h01b1a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d8e] =  Ifd35529b44c957737bf422127283c08e['h01b1c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d8f] =  Ifd35529b44c957737bf422127283c08e['h01b1e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d90] =  Ifd35529b44c957737bf422127283c08e['h01b20] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d91] =  Ifd35529b44c957737bf422127283c08e['h01b22] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d92] =  Ifd35529b44c957737bf422127283c08e['h01b24] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d93] =  Ifd35529b44c957737bf422127283c08e['h01b26] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d94] =  Ifd35529b44c957737bf422127283c08e['h01b28] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d95] =  Ifd35529b44c957737bf422127283c08e['h01b2a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d96] =  Ifd35529b44c957737bf422127283c08e['h01b2c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d97] =  Ifd35529b44c957737bf422127283c08e['h01b2e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d98] =  Ifd35529b44c957737bf422127283c08e['h01b30] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d99] =  Ifd35529b44c957737bf422127283c08e['h01b32] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d9a] =  Ifd35529b44c957737bf422127283c08e['h01b34] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d9b] =  Ifd35529b44c957737bf422127283c08e['h01b36] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d9c] =  Ifd35529b44c957737bf422127283c08e['h01b38] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d9d] =  Ifd35529b44c957737bf422127283c08e['h01b3a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d9e] =  Ifd35529b44c957737bf422127283c08e['h01b3c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00d9f] =  Ifd35529b44c957737bf422127283c08e['h01b3e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00da0] =  Ifd35529b44c957737bf422127283c08e['h01b40] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00da1] =  Ifd35529b44c957737bf422127283c08e['h01b42] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00da2] =  Ifd35529b44c957737bf422127283c08e['h01b44] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00da3] =  Ifd35529b44c957737bf422127283c08e['h01b46] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00da4] =  Ifd35529b44c957737bf422127283c08e['h01b48] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00da5] =  Ifd35529b44c957737bf422127283c08e['h01b4a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00da6] =  Ifd35529b44c957737bf422127283c08e['h01b4c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00da7] =  Ifd35529b44c957737bf422127283c08e['h01b4e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00da8] =  Ifd35529b44c957737bf422127283c08e['h01b50] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00da9] =  Ifd35529b44c957737bf422127283c08e['h01b52] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00daa] =  Ifd35529b44c957737bf422127283c08e['h01b54] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dab] =  Ifd35529b44c957737bf422127283c08e['h01b56] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dac] =  Ifd35529b44c957737bf422127283c08e['h01b58] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dad] =  Ifd35529b44c957737bf422127283c08e['h01b5a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dae] =  Ifd35529b44c957737bf422127283c08e['h01b5c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00daf] =  Ifd35529b44c957737bf422127283c08e['h01b5e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00db0] =  Ifd35529b44c957737bf422127283c08e['h01b60] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00db1] =  Ifd35529b44c957737bf422127283c08e['h01b62] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00db2] =  Ifd35529b44c957737bf422127283c08e['h01b64] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00db3] =  Ifd35529b44c957737bf422127283c08e['h01b66] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00db4] =  Ifd35529b44c957737bf422127283c08e['h01b68] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00db5] =  Ifd35529b44c957737bf422127283c08e['h01b6a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00db6] =  Ifd35529b44c957737bf422127283c08e['h01b6c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00db7] =  Ifd35529b44c957737bf422127283c08e['h01b6e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00db8] =  Ifd35529b44c957737bf422127283c08e['h01b70] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00db9] =  Ifd35529b44c957737bf422127283c08e['h01b72] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dba] =  Ifd35529b44c957737bf422127283c08e['h01b74] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dbb] =  Ifd35529b44c957737bf422127283c08e['h01b76] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dbc] =  Ifd35529b44c957737bf422127283c08e['h01b78] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dbd] =  Ifd35529b44c957737bf422127283c08e['h01b7a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dbe] =  Ifd35529b44c957737bf422127283c08e['h01b7c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dbf] =  Ifd35529b44c957737bf422127283c08e['h01b7e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dc0] =  Ifd35529b44c957737bf422127283c08e['h01b80] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dc1] =  Ifd35529b44c957737bf422127283c08e['h01b82] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dc2] =  Ifd35529b44c957737bf422127283c08e['h01b84] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dc3] =  Ifd35529b44c957737bf422127283c08e['h01b86] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dc4] =  Ifd35529b44c957737bf422127283c08e['h01b88] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dc5] =  Ifd35529b44c957737bf422127283c08e['h01b8a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dc6] =  Ifd35529b44c957737bf422127283c08e['h01b8c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dc7] =  Ifd35529b44c957737bf422127283c08e['h01b8e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dc8] =  Ifd35529b44c957737bf422127283c08e['h01b90] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dc9] =  Ifd35529b44c957737bf422127283c08e['h01b92] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dca] =  Ifd35529b44c957737bf422127283c08e['h01b94] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dcb] =  Ifd35529b44c957737bf422127283c08e['h01b96] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dcc] =  Ifd35529b44c957737bf422127283c08e['h01b98] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dcd] =  Ifd35529b44c957737bf422127283c08e['h01b9a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dce] =  Ifd35529b44c957737bf422127283c08e['h01b9c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dcf] =  Ifd35529b44c957737bf422127283c08e['h01b9e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dd0] =  Ifd35529b44c957737bf422127283c08e['h01ba0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dd1] =  Ifd35529b44c957737bf422127283c08e['h01ba2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dd2] =  Ifd35529b44c957737bf422127283c08e['h01ba4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dd3] =  Ifd35529b44c957737bf422127283c08e['h01ba6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dd4] =  Ifd35529b44c957737bf422127283c08e['h01ba8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dd5] =  Ifd35529b44c957737bf422127283c08e['h01baa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dd6] =  Ifd35529b44c957737bf422127283c08e['h01bac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dd7] =  Ifd35529b44c957737bf422127283c08e['h01bae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dd8] =  Ifd35529b44c957737bf422127283c08e['h01bb0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dd9] =  Ifd35529b44c957737bf422127283c08e['h01bb2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dda] =  Ifd35529b44c957737bf422127283c08e['h01bb4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ddb] =  Ifd35529b44c957737bf422127283c08e['h01bb6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ddc] =  Ifd35529b44c957737bf422127283c08e['h01bb8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ddd] =  Ifd35529b44c957737bf422127283c08e['h01bba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dde] =  Ifd35529b44c957737bf422127283c08e['h01bbc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ddf] =  Ifd35529b44c957737bf422127283c08e['h01bbe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00de0] =  Ifd35529b44c957737bf422127283c08e['h01bc0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00de1] =  Ifd35529b44c957737bf422127283c08e['h01bc2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00de2] =  Ifd35529b44c957737bf422127283c08e['h01bc4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00de3] =  Ifd35529b44c957737bf422127283c08e['h01bc6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00de4] =  Ifd35529b44c957737bf422127283c08e['h01bc8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00de5] =  Ifd35529b44c957737bf422127283c08e['h01bca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00de6] =  Ifd35529b44c957737bf422127283c08e['h01bcc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00de7] =  Ifd35529b44c957737bf422127283c08e['h01bce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00de8] =  Ifd35529b44c957737bf422127283c08e['h01bd0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00de9] =  Ifd35529b44c957737bf422127283c08e['h01bd2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dea] =  Ifd35529b44c957737bf422127283c08e['h01bd4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00deb] =  Ifd35529b44c957737bf422127283c08e['h01bd6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dec] =  Ifd35529b44c957737bf422127283c08e['h01bd8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ded] =  Ifd35529b44c957737bf422127283c08e['h01bda] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dee] =  Ifd35529b44c957737bf422127283c08e['h01bdc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00def] =  Ifd35529b44c957737bf422127283c08e['h01bde] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00df0] =  Ifd35529b44c957737bf422127283c08e['h01be0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00df1] =  Ifd35529b44c957737bf422127283c08e['h01be2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00df2] =  Ifd35529b44c957737bf422127283c08e['h01be4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00df3] =  Ifd35529b44c957737bf422127283c08e['h01be6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00df4] =  Ifd35529b44c957737bf422127283c08e['h01be8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00df5] =  Ifd35529b44c957737bf422127283c08e['h01bea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00df6] =  Ifd35529b44c957737bf422127283c08e['h01bec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00df7] =  Ifd35529b44c957737bf422127283c08e['h01bee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00df8] =  Ifd35529b44c957737bf422127283c08e['h01bf0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00df9] =  Ifd35529b44c957737bf422127283c08e['h01bf2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dfa] =  Ifd35529b44c957737bf422127283c08e['h01bf4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dfb] =  Ifd35529b44c957737bf422127283c08e['h01bf6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dfc] =  Ifd35529b44c957737bf422127283c08e['h01bf8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dfd] =  Ifd35529b44c957737bf422127283c08e['h01bfa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dfe] =  Ifd35529b44c957737bf422127283c08e['h01bfc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00dff] =  Ifd35529b44c957737bf422127283c08e['h01bfe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e00] =  Ifd35529b44c957737bf422127283c08e['h01c00] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e01] =  Ifd35529b44c957737bf422127283c08e['h01c02] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e02] =  Ifd35529b44c957737bf422127283c08e['h01c04] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e03] =  Ifd35529b44c957737bf422127283c08e['h01c06] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e04] =  Ifd35529b44c957737bf422127283c08e['h01c08] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e05] =  Ifd35529b44c957737bf422127283c08e['h01c0a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e06] =  Ifd35529b44c957737bf422127283c08e['h01c0c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e07] =  Ifd35529b44c957737bf422127283c08e['h01c0e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e08] =  Ifd35529b44c957737bf422127283c08e['h01c10] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e09] =  Ifd35529b44c957737bf422127283c08e['h01c12] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e0a] =  Ifd35529b44c957737bf422127283c08e['h01c14] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e0b] =  Ifd35529b44c957737bf422127283c08e['h01c16] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e0c] =  Ifd35529b44c957737bf422127283c08e['h01c18] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e0d] =  Ifd35529b44c957737bf422127283c08e['h01c1a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e0e] =  Ifd35529b44c957737bf422127283c08e['h01c1c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e0f] =  Ifd35529b44c957737bf422127283c08e['h01c1e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e10] =  Ifd35529b44c957737bf422127283c08e['h01c20] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e11] =  Ifd35529b44c957737bf422127283c08e['h01c22] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e12] =  Ifd35529b44c957737bf422127283c08e['h01c24] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e13] =  Ifd35529b44c957737bf422127283c08e['h01c26] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e14] =  Ifd35529b44c957737bf422127283c08e['h01c28] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e15] =  Ifd35529b44c957737bf422127283c08e['h01c2a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e16] =  Ifd35529b44c957737bf422127283c08e['h01c2c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e17] =  Ifd35529b44c957737bf422127283c08e['h01c2e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e18] =  Ifd35529b44c957737bf422127283c08e['h01c30] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e19] =  Ifd35529b44c957737bf422127283c08e['h01c32] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e1a] =  Ifd35529b44c957737bf422127283c08e['h01c34] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e1b] =  Ifd35529b44c957737bf422127283c08e['h01c36] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e1c] =  Ifd35529b44c957737bf422127283c08e['h01c38] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e1d] =  Ifd35529b44c957737bf422127283c08e['h01c3a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e1e] =  Ifd35529b44c957737bf422127283c08e['h01c3c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e1f] =  Ifd35529b44c957737bf422127283c08e['h01c3e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e20] =  Ifd35529b44c957737bf422127283c08e['h01c40] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e21] =  Ifd35529b44c957737bf422127283c08e['h01c42] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e22] =  Ifd35529b44c957737bf422127283c08e['h01c44] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e23] =  Ifd35529b44c957737bf422127283c08e['h01c46] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e24] =  Ifd35529b44c957737bf422127283c08e['h01c48] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e25] =  Ifd35529b44c957737bf422127283c08e['h01c4a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e26] =  Ifd35529b44c957737bf422127283c08e['h01c4c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e27] =  Ifd35529b44c957737bf422127283c08e['h01c4e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e28] =  Ifd35529b44c957737bf422127283c08e['h01c50] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e29] =  Ifd35529b44c957737bf422127283c08e['h01c52] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e2a] =  Ifd35529b44c957737bf422127283c08e['h01c54] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e2b] =  Ifd35529b44c957737bf422127283c08e['h01c56] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e2c] =  Ifd35529b44c957737bf422127283c08e['h01c58] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e2d] =  Ifd35529b44c957737bf422127283c08e['h01c5a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e2e] =  Ifd35529b44c957737bf422127283c08e['h01c5c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e2f] =  Ifd35529b44c957737bf422127283c08e['h01c5e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e30] =  Ifd35529b44c957737bf422127283c08e['h01c60] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e31] =  Ifd35529b44c957737bf422127283c08e['h01c62] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e32] =  Ifd35529b44c957737bf422127283c08e['h01c64] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e33] =  Ifd35529b44c957737bf422127283c08e['h01c66] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e34] =  Ifd35529b44c957737bf422127283c08e['h01c68] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e35] =  Ifd35529b44c957737bf422127283c08e['h01c6a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e36] =  Ifd35529b44c957737bf422127283c08e['h01c6c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e37] =  Ifd35529b44c957737bf422127283c08e['h01c6e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e38] =  Ifd35529b44c957737bf422127283c08e['h01c70] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e39] =  Ifd35529b44c957737bf422127283c08e['h01c72] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e3a] =  Ifd35529b44c957737bf422127283c08e['h01c74] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e3b] =  Ifd35529b44c957737bf422127283c08e['h01c76] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e3c] =  Ifd35529b44c957737bf422127283c08e['h01c78] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e3d] =  Ifd35529b44c957737bf422127283c08e['h01c7a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e3e] =  Ifd35529b44c957737bf422127283c08e['h01c7c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e3f] =  Ifd35529b44c957737bf422127283c08e['h01c7e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e40] =  Ifd35529b44c957737bf422127283c08e['h01c80] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e41] =  Ifd35529b44c957737bf422127283c08e['h01c82] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e42] =  Ifd35529b44c957737bf422127283c08e['h01c84] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e43] =  Ifd35529b44c957737bf422127283c08e['h01c86] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e44] =  Ifd35529b44c957737bf422127283c08e['h01c88] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e45] =  Ifd35529b44c957737bf422127283c08e['h01c8a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e46] =  Ifd35529b44c957737bf422127283c08e['h01c8c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e47] =  Ifd35529b44c957737bf422127283c08e['h01c8e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e48] =  Ifd35529b44c957737bf422127283c08e['h01c90] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e49] =  Ifd35529b44c957737bf422127283c08e['h01c92] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e4a] =  Ifd35529b44c957737bf422127283c08e['h01c94] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e4b] =  Ifd35529b44c957737bf422127283c08e['h01c96] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e4c] =  Ifd35529b44c957737bf422127283c08e['h01c98] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e4d] =  Ifd35529b44c957737bf422127283c08e['h01c9a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e4e] =  Ifd35529b44c957737bf422127283c08e['h01c9c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e4f] =  Ifd35529b44c957737bf422127283c08e['h01c9e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e50] =  Ifd35529b44c957737bf422127283c08e['h01ca0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e51] =  Ifd35529b44c957737bf422127283c08e['h01ca2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e52] =  Ifd35529b44c957737bf422127283c08e['h01ca4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e53] =  Ifd35529b44c957737bf422127283c08e['h01ca6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e54] =  Ifd35529b44c957737bf422127283c08e['h01ca8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e55] =  Ifd35529b44c957737bf422127283c08e['h01caa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e56] =  Ifd35529b44c957737bf422127283c08e['h01cac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e57] =  Ifd35529b44c957737bf422127283c08e['h01cae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e58] =  Ifd35529b44c957737bf422127283c08e['h01cb0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e59] =  Ifd35529b44c957737bf422127283c08e['h01cb2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e5a] =  Ifd35529b44c957737bf422127283c08e['h01cb4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e5b] =  Ifd35529b44c957737bf422127283c08e['h01cb6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e5c] =  Ifd35529b44c957737bf422127283c08e['h01cb8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e5d] =  Ifd35529b44c957737bf422127283c08e['h01cba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e5e] =  Ifd35529b44c957737bf422127283c08e['h01cbc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e5f] =  Ifd35529b44c957737bf422127283c08e['h01cbe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e60] =  Ifd35529b44c957737bf422127283c08e['h01cc0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e61] =  Ifd35529b44c957737bf422127283c08e['h01cc2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e62] =  Ifd35529b44c957737bf422127283c08e['h01cc4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e63] =  Ifd35529b44c957737bf422127283c08e['h01cc6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e64] =  Ifd35529b44c957737bf422127283c08e['h01cc8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e65] =  Ifd35529b44c957737bf422127283c08e['h01cca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e66] =  Ifd35529b44c957737bf422127283c08e['h01ccc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e67] =  Ifd35529b44c957737bf422127283c08e['h01cce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e68] =  Ifd35529b44c957737bf422127283c08e['h01cd0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e69] =  Ifd35529b44c957737bf422127283c08e['h01cd2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e6a] =  Ifd35529b44c957737bf422127283c08e['h01cd4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e6b] =  Ifd35529b44c957737bf422127283c08e['h01cd6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e6c] =  Ifd35529b44c957737bf422127283c08e['h01cd8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e6d] =  Ifd35529b44c957737bf422127283c08e['h01cda] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e6e] =  Ifd35529b44c957737bf422127283c08e['h01cdc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e6f] =  Ifd35529b44c957737bf422127283c08e['h01cde] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e70] =  Ifd35529b44c957737bf422127283c08e['h01ce0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e71] =  Ifd35529b44c957737bf422127283c08e['h01ce2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e72] =  Ifd35529b44c957737bf422127283c08e['h01ce4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e73] =  Ifd35529b44c957737bf422127283c08e['h01ce6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e74] =  Ifd35529b44c957737bf422127283c08e['h01ce8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e75] =  Ifd35529b44c957737bf422127283c08e['h01cea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e76] =  Ifd35529b44c957737bf422127283c08e['h01cec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e77] =  Ifd35529b44c957737bf422127283c08e['h01cee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e78] =  Ifd35529b44c957737bf422127283c08e['h01cf0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e79] =  Ifd35529b44c957737bf422127283c08e['h01cf2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e7a] =  Ifd35529b44c957737bf422127283c08e['h01cf4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e7b] =  Ifd35529b44c957737bf422127283c08e['h01cf6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e7c] =  Ifd35529b44c957737bf422127283c08e['h01cf8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e7d] =  Ifd35529b44c957737bf422127283c08e['h01cfa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e7e] =  Ifd35529b44c957737bf422127283c08e['h01cfc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e7f] =  Ifd35529b44c957737bf422127283c08e['h01cfe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e80] =  Ifd35529b44c957737bf422127283c08e['h01d00] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e81] =  Ifd35529b44c957737bf422127283c08e['h01d02] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e82] =  Ifd35529b44c957737bf422127283c08e['h01d04] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e83] =  Ifd35529b44c957737bf422127283c08e['h01d06] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e84] =  Ifd35529b44c957737bf422127283c08e['h01d08] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e85] =  Ifd35529b44c957737bf422127283c08e['h01d0a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e86] =  Ifd35529b44c957737bf422127283c08e['h01d0c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e87] =  Ifd35529b44c957737bf422127283c08e['h01d0e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e88] =  Ifd35529b44c957737bf422127283c08e['h01d10] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e89] =  Ifd35529b44c957737bf422127283c08e['h01d12] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e8a] =  Ifd35529b44c957737bf422127283c08e['h01d14] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e8b] =  Ifd35529b44c957737bf422127283c08e['h01d16] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e8c] =  Ifd35529b44c957737bf422127283c08e['h01d18] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e8d] =  Ifd35529b44c957737bf422127283c08e['h01d1a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e8e] =  Ifd35529b44c957737bf422127283c08e['h01d1c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e8f] =  Ifd35529b44c957737bf422127283c08e['h01d1e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e90] =  Ifd35529b44c957737bf422127283c08e['h01d20] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e91] =  Ifd35529b44c957737bf422127283c08e['h01d22] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e92] =  Ifd35529b44c957737bf422127283c08e['h01d24] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e93] =  Ifd35529b44c957737bf422127283c08e['h01d26] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e94] =  Ifd35529b44c957737bf422127283c08e['h01d28] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e95] =  Ifd35529b44c957737bf422127283c08e['h01d2a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e96] =  Ifd35529b44c957737bf422127283c08e['h01d2c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e97] =  Ifd35529b44c957737bf422127283c08e['h01d2e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e98] =  Ifd35529b44c957737bf422127283c08e['h01d30] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e99] =  Ifd35529b44c957737bf422127283c08e['h01d32] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e9a] =  Ifd35529b44c957737bf422127283c08e['h01d34] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e9b] =  Ifd35529b44c957737bf422127283c08e['h01d36] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e9c] =  Ifd35529b44c957737bf422127283c08e['h01d38] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e9d] =  Ifd35529b44c957737bf422127283c08e['h01d3a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e9e] =  Ifd35529b44c957737bf422127283c08e['h01d3c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00e9f] =  Ifd35529b44c957737bf422127283c08e['h01d3e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ea0] =  Ifd35529b44c957737bf422127283c08e['h01d40] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ea1] =  Ifd35529b44c957737bf422127283c08e['h01d42] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ea2] =  Ifd35529b44c957737bf422127283c08e['h01d44] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ea3] =  Ifd35529b44c957737bf422127283c08e['h01d46] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ea4] =  Ifd35529b44c957737bf422127283c08e['h01d48] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ea5] =  Ifd35529b44c957737bf422127283c08e['h01d4a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ea6] =  Ifd35529b44c957737bf422127283c08e['h01d4c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ea7] =  Ifd35529b44c957737bf422127283c08e['h01d4e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ea8] =  Ifd35529b44c957737bf422127283c08e['h01d50] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ea9] =  Ifd35529b44c957737bf422127283c08e['h01d52] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00eaa] =  Ifd35529b44c957737bf422127283c08e['h01d54] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00eab] =  Ifd35529b44c957737bf422127283c08e['h01d56] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00eac] =  Ifd35529b44c957737bf422127283c08e['h01d58] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ead] =  Ifd35529b44c957737bf422127283c08e['h01d5a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00eae] =  Ifd35529b44c957737bf422127283c08e['h01d5c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00eaf] =  Ifd35529b44c957737bf422127283c08e['h01d5e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00eb0] =  Ifd35529b44c957737bf422127283c08e['h01d60] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00eb1] =  Ifd35529b44c957737bf422127283c08e['h01d62] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00eb2] =  Ifd35529b44c957737bf422127283c08e['h01d64] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00eb3] =  Ifd35529b44c957737bf422127283c08e['h01d66] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00eb4] =  Ifd35529b44c957737bf422127283c08e['h01d68] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00eb5] =  Ifd35529b44c957737bf422127283c08e['h01d6a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00eb6] =  Ifd35529b44c957737bf422127283c08e['h01d6c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00eb7] =  Ifd35529b44c957737bf422127283c08e['h01d6e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00eb8] =  Ifd35529b44c957737bf422127283c08e['h01d70] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00eb9] =  Ifd35529b44c957737bf422127283c08e['h01d72] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00eba] =  Ifd35529b44c957737bf422127283c08e['h01d74] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ebb] =  Ifd35529b44c957737bf422127283c08e['h01d76] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ebc] =  Ifd35529b44c957737bf422127283c08e['h01d78] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ebd] =  Ifd35529b44c957737bf422127283c08e['h01d7a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ebe] =  Ifd35529b44c957737bf422127283c08e['h01d7c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ebf] =  Ifd35529b44c957737bf422127283c08e['h01d7e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ec0] =  Ifd35529b44c957737bf422127283c08e['h01d80] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ec1] =  Ifd35529b44c957737bf422127283c08e['h01d82] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ec2] =  Ifd35529b44c957737bf422127283c08e['h01d84] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ec3] =  Ifd35529b44c957737bf422127283c08e['h01d86] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ec4] =  Ifd35529b44c957737bf422127283c08e['h01d88] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ec5] =  Ifd35529b44c957737bf422127283c08e['h01d8a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ec6] =  Ifd35529b44c957737bf422127283c08e['h01d8c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ec7] =  Ifd35529b44c957737bf422127283c08e['h01d8e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ec8] =  Ifd35529b44c957737bf422127283c08e['h01d90] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ec9] =  Ifd35529b44c957737bf422127283c08e['h01d92] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00eca] =  Ifd35529b44c957737bf422127283c08e['h01d94] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ecb] =  Ifd35529b44c957737bf422127283c08e['h01d96] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ecc] =  Ifd35529b44c957737bf422127283c08e['h01d98] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ecd] =  Ifd35529b44c957737bf422127283c08e['h01d9a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ece] =  Ifd35529b44c957737bf422127283c08e['h01d9c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ecf] =  Ifd35529b44c957737bf422127283c08e['h01d9e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ed0] =  Ifd35529b44c957737bf422127283c08e['h01da0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ed1] =  Ifd35529b44c957737bf422127283c08e['h01da2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ed2] =  Ifd35529b44c957737bf422127283c08e['h01da4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ed3] =  Ifd35529b44c957737bf422127283c08e['h01da6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ed4] =  Ifd35529b44c957737bf422127283c08e['h01da8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ed5] =  Ifd35529b44c957737bf422127283c08e['h01daa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ed6] =  Ifd35529b44c957737bf422127283c08e['h01dac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ed7] =  Ifd35529b44c957737bf422127283c08e['h01dae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ed8] =  Ifd35529b44c957737bf422127283c08e['h01db0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ed9] =  Ifd35529b44c957737bf422127283c08e['h01db2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00eda] =  Ifd35529b44c957737bf422127283c08e['h01db4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00edb] =  Ifd35529b44c957737bf422127283c08e['h01db6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00edc] =  Ifd35529b44c957737bf422127283c08e['h01db8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00edd] =  Ifd35529b44c957737bf422127283c08e['h01dba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ede] =  Ifd35529b44c957737bf422127283c08e['h01dbc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00edf] =  Ifd35529b44c957737bf422127283c08e['h01dbe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ee0] =  Ifd35529b44c957737bf422127283c08e['h01dc0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ee1] =  Ifd35529b44c957737bf422127283c08e['h01dc2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ee2] =  Ifd35529b44c957737bf422127283c08e['h01dc4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ee3] =  Ifd35529b44c957737bf422127283c08e['h01dc6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ee4] =  Ifd35529b44c957737bf422127283c08e['h01dc8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ee5] =  Ifd35529b44c957737bf422127283c08e['h01dca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ee6] =  Ifd35529b44c957737bf422127283c08e['h01dcc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ee7] =  Ifd35529b44c957737bf422127283c08e['h01dce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ee8] =  Ifd35529b44c957737bf422127283c08e['h01dd0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ee9] =  Ifd35529b44c957737bf422127283c08e['h01dd2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00eea] =  Ifd35529b44c957737bf422127283c08e['h01dd4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00eeb] =  Ifd35529b44c957737bf422127283c08e['h01dd6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00eec] =  Ifd35529b44c957737bf422127283c08e['h01dd8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00eed] =  Ifd35529b44c957737bf422127283c08e['h01dda] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00eee] =  Ifd35529b44c957737bf422127283c08e['h01ddc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00eef] =  Ifd35529b44c957737bf422127283c08e['h01dde] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ef0] =  Ifd35529b44c957737bf422127283c08e['h01de0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ef1] =  Ifd35529b44c957737bf422127283c08e['h01de2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ef2] =  Ifd35529b44c957737bf422127283c08e['h01de4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ef3] =  Ifd35529b44c957737bf422127283c08e['h01de6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ef4] =  Ifd35529b44c957737bf422127283c08e['h01de8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ef5] =  Ifd35529b44c957737bf422127283c08e['h01dea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ef6] =  Ifd35529b44c957737bf422127283c08e['h01dec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ef7] =  Ifd35529b44c957737bf422127283c08e['h01dee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ef8] =  Ifd35529b44c957737bf422127283c08e['h01df0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ef9] =  Ifd35529b44c957737bf422127283c08e['h01df2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00efa] =  Ifd35529b44c957737bf422127283c08e['h01df4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00efb] =  Ifd35529b44c957737bf422127283c08e['h01df6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00efc] =  Ifd35529b44c957737bf422127283c08e['h01df8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00efd] =  Ifd35529b44c957737bf422127283c08e['h01dfa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00efe] =  Ifd35529b44c957737bf422127283c08e['h01dfc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00eff] =  Ifd35529b44c957737bf422127283c08e['h01dfe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f00] =  Ifd35529b44c957737bf422127283c08e['h01e00] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f01] =  Ifd35529b44c957737bf422127283c08e['h01e02] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f02] =  Ifd35529b44c957737bf422127283c08e['h01e04] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f03] =  Ifd35529b44c957737bf422127283c08e['h01e06] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f04] =  Ifd35529b44c957737bf422127283c08e['h01e08] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f05] =  Ifd35529b44c957737bf422127283c08e['h01e0a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f06] =  Ifd35529b44c957737bf422127283c08e['h01e0c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f07] =  Ifd35529b44c957737bf422127283c08e['h01e0e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f08] =  Ifd35529b44c957737bf422127283c08e['h01e10] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f09] =  Ifd35529b44c957737bf422127283c08e['h01e12] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f0a] =  Ifd35529b44c957737bf422127283c08e['h01e14] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f0b] =  Ifd35529b44c957737bf422127283c08e['h01e16] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f0c] =  Ifd35529b44c957737bf422127283c08e['h01e18] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f0d] =  Ifd35529b44c957737bf422127283c08e['h01e1a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f0e] =  Ifd35529b44c957737bf422127283c08e['h01e1c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f0f] =  Ifd35529b44c957737bf422127283c08e['h01e1e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f10] =  Ifd35529b44c957737bf422127283c08e['h01e20] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f11] =  Ifd35529b44c957737bf422127283c08e['h01e22] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f12] =  Ifd35529b44c957737bf422127283c08e['h01e24] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f13] =  Ifd35529b44c957737bf422127283c08e['h01e26] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f14] =  Ifd35529b44c957737bf422127283c08e['h01e28] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f15] =  Ifd35529b44c957737bf422127283c08e['h01e2a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f16] =  Ifd35529b44c957737bf422127283c08e['h01e2c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f17] =  Ifd35529b44c957737bf422127283c08e['h01e2e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f18] =  Ifd35529b44c957737bf422127283c08e['h01e30] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f19] =  Ifd35529b44c957737bf422127283c08e['h01e32] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f1a] =  Ifd35529b44c957737bf422127283c08e['h01e34] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f1b] =  Ifd35529b44c957737bf422127283c08e['h01e36] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f1c] =  Ifd35529b44c957737bf422127283c08e['h01e38] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f1d] =  Ifd35529b44c957737bf422127283c08e['h01e3a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f1e] =  Ifd35529b44c957737bf422127283c08e['h01e3c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f1f] =  Ifd35529b44c957737bf422127283c08e['h01e3e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f20] =  Ifd35529b44c957737bf422127283c08e['h01e40] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f21] =  Ifd35529b44c957737bf422127283c08e['h01e42] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f22] =  Ifd35529b44c957737bf422127283c08e['h01e44] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f23] =  Ifd35529b44c957737bf422127283c08e['h01e46] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f24] =  Ifd35529b44c957737bf422127283c08e['h01e48] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f25] =  Ifd35529b44c957737bf422127283c08e['h01e4a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f26] =  Ifd35529b44c957737bf422127283c08e['h01e4c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f27] =  Ifd35529b44c957737bf422127283c08e['h01e4e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f28] =  Ifd35529b44c957737bf422127283c08e['h01e50] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f29] =  Ifd35529b44c957737bf422127283c08e['h01e52] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f2a] =  Ifd35529b44c957737bf422127283c08e['h01e54] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f2b] =  Ifd35529b44c957737bf422127283c08e['h01e56] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f2c] =  Ifd35529b44c957737bf422127283c08e['h01e58] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f2d] =  Ifd35529b44c957737bf422127283c08e['h01e5a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f2e] =  Ifd35529b44c957737bf422127283c08e['h01e5c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f2f] =  Ifd35529b44c957737bf422127283c08e['h01e5e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f30] =  Ifd35529b44c957737bf422127283c08e['h01e60] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f31] =  Ifd35529b44c957737bf422127283c08e['h01e62] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f32] =  Ifd35529b44c957737bf422127283c08e['h01e64] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f33] =  Ifd35529b44c957737bf422127283c08e['h01e66] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f34] =  Ifd35529b44c957737bf422127283c08e['h01e68] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f35] =  Ifd35529b44c957737bf422127283c08e['h01e6a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f36] =  Ifd35529b44c957737bf422127283c08e['h01e6c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f37] =  Ifd35529b44c957737bf422127283c08e['h01e6e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f38] =  Ifd35529b44c957737bf422127283c08e['h01e70] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f39] =  Ifd35529b44c957737bf422127283c08e['h01e72] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f3a] =  Ifd35529b44c957737bf422127283c08e['h01e74] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f3b] =  Ifd35529b44c957737bf422127283c08e['h01e76] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f3c] =  Ifd35529b44c957737bf422127283c08e['h01e78] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f3d] =  Ifd35529b44c957737bf422127283c08e['h01e7a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f3e] =  Ifd35529b44c957737bf422127283c08e['h01e7c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f3f] =  Ifd35529b44c957737bf422127283c08e['h01e7e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f40] =  Ifd35529b44c957737bf422127283c08e['h01e80] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f41] =  Ifd35529b44c957737bf422127283c08e['h01e82] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f42] =  Ifd35529b44c957737bf422127283c08e['h01e84] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f43] =  Ifd35529b44c957737bf422127283c08e['h01e86] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f44] =  Ifd35529b44c957737bf422127283c08e['h01e88] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f45] =  Ifd35529b44c957737bf422127283c08e['h01e8a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f46] =  Ifd35529b44c957737bf422127283c08e['h01e8c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f47] =  Ifd35529b44c957737bf422127283c08e['h01e8e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f48] =  Ifd35529b44c957737bf422127283c08e['h01e90] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f49] =  Ifd35529b44c957737bf422127283c08e['h01e92] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f4a] =  Ifd35529b44c957737bf422127283c08e['h01e94] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f4b] =  Ifd35529b44c957737bf422127283c08e['h01e96] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f4c] =  Ifd35529b44c957737bf422127283c08e['h01e98] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f4d] =  Ifd35529b44c957737bf422127283c08e['h01e9a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f4e] =  Ifd35529b44c957737bf422127283c08e['h01e9c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f4f] =  Ifd35529b44c957737bf422127283c08e['h01e9e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f50] =  Ifd35529b44c957737bf422127283c08e['h01ea0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f51] =  Ifd35529b44c957737bf422127283c08e['h01ea2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f52] =  Ifd35529b44c957737bf422127283c08e['h01ea4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f53] =  Ifd35529b44c957737bf422127283c08e['h01ea6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f54] =  Ifd35529b44c957737bf422127283c08e['h01ea8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f55] =  Ifd35529b44c957737bf422127283c08e['h01eaa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f56] =  Ifd35529b44c957737bf422127283c08e['h01eac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f57] =  Ifd35529b44c957737bf422127283c08e['h01eae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f58] =  Ifd35529b44c957737bf422127283c08e['h01eb0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f59] =  Ifd35529b44c957737bf422127283c08e['h01eb2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f5a] =  Ifd35529b44c957737bf422127283c08e['h01eb4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f5b] =  Ifd35529b44c957737bf422127283c08e['h01eb6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f5c] =  Ifd35529b44c957737bf422127283c08e['h01eb8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f5d] =  Ifd35529b44c957737bf422127283c08e['h01eba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f5e] =  Ifd35529b44c957737bf422127283c08e['h01ebc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f5f] =  Ifd35529b44c957737bf422127283c08e['h01ebe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f60] =  Ifd35529b44c957737bf422127283c08e['h01ec0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f61] =  Ifd35529b44c957737bf422127283c08e['h01ec2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f62] =  Ifd35529b44c957737bf422127283c08e['h01ec4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f63] =  Ifd35529b44c957737bf422127283c08e['h01ec6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f64] =  Ifd35529b44c957737bf422127283c08e['h01ec8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f65] =  Ifd35529b44c957737bf422127283c08e['h01eca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f66] =  Ifd35529b44c957737bf422127283c08e['h01ecc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f67] =  Ifd35529b44c957737bf422127283c08e['h01ece] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f68] =  Ifd35529b44c957737bf422127283c08e['h01ed0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f69] =  Ifd35529b44c957737bf422127283c08e['h01ed2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f6a] =  Ifd35529b44c957737bf422127283c08e['h01ed4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f6b] =  Ifd35529b44c957737bf422127283c08e['h01ed6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f6c] =  Ifd35529b44c957737bf422127283c08e['h01ed8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f6d] =  Ifd35529b44c957737bf422127283c08e['h01eda] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f6e] =  Ifd35529b44c957737bf422127283c08e['h01edc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f6f] =  Ifd35529b44c957737bf422127283c08e['h01ede] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f70] =  Ifd35529b44c957737bf422127283c08e['h01ee0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f71] =  Ifd35529b44c957737bf422127283c08e['h01ee2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f72] =  Ifd35529b44c957737bf422127283c08e['h01ee4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f73] =  Ifd35529b44c957737bf422127283c08e['h01ee6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f74] =  Ifd35529b44c957737bf422127283c08e['h01ee8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f75] =  Ifd35529b44c957737bf422127283c08e['h01eea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f76] =  Ifd35529b44c957737bf422127283c08e['h01eec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f77] =  Ifd35529b44c957737bf422127283c08e['h01eee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f78] =  Ifd35529b44c957737bf422127283c08e['h01ef0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f79] =  Ifd35529b44c957737bf422127283c08e['h01ef2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f7a] =  Ifd35529b44c957737bf422127283c08e['h01ef4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f7b] =  Ifd35529b44c957737bf422127283c08e['h01ef6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f7c] =  Ifd35529b44c957737bf422127283c08e['h01ef8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f7d] =  Ifd35529b44c957737bf422127283c08e['h01efa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f7e] =  Ifd35529b44c957737bf422127283c08e['h01efc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f7f] =  Ifd35529b44c957737bf422127283c08e['h01efe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f80] =  Ifd35529b44c957737bf422127283c08e['h01f00] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f81] =  Ifd35529b44c957737bf422127283c08e['h01f02] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f82] =  Ifd35529b44c957737bf422127283c08e['h01f04] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f83] =  Ifd35529b44c957737bf422127283c08e['h01f06] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f84] =  Ifd35529b44c957737bf422127283c08e['h01f08] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f85] =  Ifd35529b44c957737bf422127283c08e['h01f0a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f86] =  Ifd35529b44c957737bf422127283c08e['h01f0c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f87] =  Ifd35529b44c957737bf422127283c08e['h01f0e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f88] =  Ifd35529b44c957737bf422127283c08e['h01f10] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f89] =  Ifd35529b44c957737bf422127283c08e['h01f12] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f8a] =  Ifd35529b44c957737bf422127283c08e['h01f14] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f8b] =  Ifd35529b44c957737bf422127283c08e['h01f16] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f8c] =  Ifd35529b44c957737bf422127283c08e['h01f18] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f8d] =  Ifd35529b44c957737bf422127283c08e['h01f1a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f8e] =  Ifd35529b44c957737bf422127283c08e['h01f1c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f8f] =  Ifd35529b44c957737bf422127283c08e['h01f1e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f90] =  Ifd35529b44c957737bf422127283c08e['h01f20] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f91] =  Ifd35529b44c957737bf422127283c08e['h01f22] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f92] =  Ifd35529b44c957737bf422127283c08e['h01f24] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f93] =  Ifd35529b44c957737bf422127283c08e['h01f26] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f94] =  Ifd35529b44c957737bf422127283c08e['h01f28] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f95] =  Ifd35529b44c957737bf422127283c08e['h01f2a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f96] =  Ifd35529b44c957737bf422127283c08e['h01f2c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f97] =  Ifd35529b44c957737bf422127283c08e['h01f2e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f98] =  Ifd35529b44c957737bf422127283c08e['h01f30] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f99] =  Ifd35529b44c957737bf422127283c08e['h01f32] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f9a] =  Ifd35529b44c957737bf422127283c08e['h01f34] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f9b] =  Ifd35529b44c957737bf422127283c08e['h01f36] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f9c] =  Ifd35529b44c957737bf422127283c08e['h01f38] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f9d] =  Ifd35529b44c957737bf422127283c08e['h01f3a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f9e] =  Ifd35529b44c957737bf422127283c08e['h01f3c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00f9f] =  Ifd35529b44c957737bf422127283c08e['h01f3e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fa0] =  Ifd35529b44c957737bf422127283c08e['h01f40] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fa1] =  Ifd35529b44c957737bf422127283c08e['h01f42] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fa2] =  Ifd35529b44c957737bf422127283c08e['h01f44] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fa3] =  Ifd35529b44c957737bf422127283c08e['h01f46] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fa4] =  Ifd35529b44c957737bf422127283c08e['h01f48] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fa5] =  Ifd35529b44c957737bf422127283c08e['h01f4a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fa6] =  Ifd35529b44c957737bf422127283c08e['h01f4c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fa7] =  Ifd35529b44c957737bf422127283c08e['h01f4e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fa8] =  Ifd35529b44c957737bf422127283c08e['h01f50] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fa9] =  Ifd35529b44c957737bf422127283c08e['h01f52] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00faa] =  Ifd35529b44c957737bf422127283c08e['h01f54] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fab] =  Ifd35529b44c957737bf422127283c08e['h01f56] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fac] =  Ifd35529b44c957737bf422127283c08e['h01f58] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fad] =  Ifd35529b44c957737bf422127283c08e['h01f5a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fae] =  Ifd35529b44c957737bf422127283c08e['h01f5c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00faf] =  Ifd35529b44c957737bf422127283c08e['h01f5e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fb0] =  Ifd35529b44c957737bf422127283c08e['h01f60] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fb1] =  Ifd35529b44c957737bf422127283c08e['h01f62] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fb2] =  Ifd35529b44c957737bf422127283c08e['h01f64] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fb3] =  Ifd35529b44c957737bf422127283c08e['h01f66] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fb4] =  Ifd35529b44c957737bf422127283c08e['h01f68] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fb5] =  Ifd35529b44c957737bf422127283c08e['h01f6a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fb6] =  Ifd35529b44c957737bf422127283c08e['h01f6c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fb7] =  Ifd35529b44c957737bf422127283c08e['h01f6e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fb8] =  Ifd35529b44c957737bf422127283c08e['h01f70] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fb9] =  Ifd35529b44c957737bf422127283c08e['h01f72] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fba] =  Ifd35529b44c957737bf422127283c08e['h01f74] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fbb] =  Ifd35529b44c957737bf422127283c08e['h01f76] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fbc] =  Ifd35529b44c957737bf422127283c08e['h01f78] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fbd] =  Ifd35529b44c957737bf422127283c08e['h01f7a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fbe] =  Ifd35529b44c957737bf422127283c08e['h01f7c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fbf] =  Ifd35529b44c957737bf422127283c08e['h01f7e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fc0] =  Ifd35529b44c957737bf422127283c08e['h01f80] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fc1] =  Ifd35529b44c957737bf422127283c08e['h01f82] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fc2] =  Ifd35529b44c957737bf422127283c08e['h01f84] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fc3] =  Ifd35529b44c957737bf422127283c08e['h01f86] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fc4] =  Ifd35529b44c957737bf422127283c08e['h01f88] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fc5] =  Ifd35529b44c957737bf422127283c08e['h01f8a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fc6] =  Ifd35529b44c957737bf422127283c08e['h01f8c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fc7] =  Ifd35529b44c957737bf422127283c08e['h01f8e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fc8] =  Ifd35529b44c957737bf422127283c08e['h01f90] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fc9] =  Ifd35529b44c957737bf422127283c08e['h01f92] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fca] =  Ifd35529b44c957737bf422127283c08e['h01f94] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fcb] =  Ifd35529b44c957737bf422127283c08e['h01f96] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fcc] =  Ifd35529b44c957737bf422127283c08e['h01f98] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fcd] =  Ifd35529b44c957737bf422127283c08e['h01f9a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fce] =  Ifd35529b44c957737bf422127283c08e['h01f9c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fcf] =  Ifd35529b44c957737bf422127283c08e['h01f9e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fd0] =  Ifd35529b44c957737bf422127283c08e['h01fa0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fd1] =  Ifd35529b44c957737bf422127283c08e['h01fa2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fd2] =  Ifd35529b44c957737bf422127283c08e['h01fa4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fd3] =  Ifd35529b44c957737bf422127283c08e['h01fa6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fd4] =  Ifd35529b44c957737bf422127283c08e['h01fa8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fd5] =  Ifd35529b44c957737bf422127283c08e['h01faa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fd6] =  Ifd35529b44c957737bf422127283c08e['h01fac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fd7] =  Ifd35529b44c957737bf422127283c08e['h01fae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fd8] =  Ifd35529b44c957737bf422127283c08e['h01fb0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fd9] =  Ifd35529b44c957737bf422127283c08e['h01fb2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fda] =  Ifd35529b44c957737bf422127283c08e['h01fb4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fdb] =  Ifd35529b44c957737bf422127283c08e['h01fb6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fdc] =  Ifd35529b44c957737bf422127283c08e['h01fb8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fdd] =  Ifd35529b44c957737bf422127283c08e['h01fba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fde] =  Ifd35529b44c957737bf422127283c08e['h01fbc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fdf] =  Ifd35529b44c957737bf422127283c08e['h01fbe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fe0] =  Ifd35529b44c957737bf422127283c08e['h01fc0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fe1] =  Ifd35529b44c957737bf422127283c08e['h01fc2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fe2] =  Ifd35529b44c957737bf422127283c08e['h01fc4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fe3] =  Ifd35529b44c957737bf422127283c08e['h01fc6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fe4] =  Ifd35529b44c957737bf422127283c08e['h01fc8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fe5] =  Ifd35529b44c957737bf422127283c08e['h01fca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fe6] =  Ifd35529b44c957737bf422127283c08e['h01fcc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fe7] =  Ifd35529b44c957737bf422127283c08e['h01fce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fe8] =  Ifd35529b44c957737bf422127283c08e['h01fd0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fe9] =  Ifd35529b44c957737bf422127283c08e['h01fd2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fea] =  Ifd35529b44c957737bf422127283c08e['h01fd4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00feb] =  Ifd35529b44c957737bf422127283c08e['h01fd6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fec] =  Ifd35529b44c957737bf422127283c08e['h01fd8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fed] =  Ifd35529b44c957737bf422127283c08e['h01fda] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fee] =  Ifd35529b44c957737bf422127283c08e['h01fdc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fef] =  Ifd35529b44c957737bf422127283c08e['h01fde] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ff0] =  Ifd35529b44c957737bf422127283c08e['h01fe0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ff1] =  Ifd35529b44c957737bf422127283c08e['h01fe2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ff2] =  Ifd35529b44c957737bf422127283c08e['h01fe4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ff3] =  Ifd35529b44c957737bf422127283c08e['h01fe6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ff4] =  Ifd35529b44c957737bf422127283c08e['h01fe8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ff5] =  Ifd35529b44c957737bf422127283c08e['h01fea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ff6] =  Ifd35529b44c957737bf422127283c08e['h01fec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ff7] =  Ifd35529b44c957737bf422127283c08e['h01fee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ff8] =  Ifd35529b44c957737bf422127283c08e['h01ff0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ff9] =  Ifd35529b44c957737bf422127283c08e['h01ff2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ffa] =  Ifd35529b44c957737bf422127283c08e['h01ff4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ffb] =  Ifd35529b44c957737bf422127283c08e['h01ff6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ffc] =  Ifd35529b44c957737bf422127283c08e['h01ff8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ffd] =  Ifd35529b44c957737bf422127283c08e['h01ffa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00ffe] =  Ifd35529b44c957737bf422127283c08e['h01ffc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h00fff] =  Ifd35529b44c957737bf422127283c08e['h01ffe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01000] =  Ifd35529b44c957737bf422127283c08e['h02000] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01001] =  Ifd35529b44c957737bf422127283c08e['h02002] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01002] =  Ifd35529b44c957737bf422127283c08e['h02004] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01003] =  Ifd35529b44c957737bf422127283c08e['h02006] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01004] =  Ifd35529b44c957737bf422127283c08e['h02008] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01005] =  Ifd35529b44c957737bf422127283c08e['h0200a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01006] =  Ifd35529b44c957737bf422127283c08e['h0200c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01007] =  Ifd35529b44c957737bf422127283c08e['h0200e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01008] =  Ifd35529b44c957737bf422127283c08e['h02010] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01009] =  Ifd35529b44c957737bf422127283c08e['h02012] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0100a] =  Ifd35529b44c957737bf422127283c08e['h02014] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0100b] =  Ifd35529b44c957737bf422127283c08e['h02016] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0100c] =  Ifd35529b44c957737bf422127283c08e['h02018] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0100d] =  Ifd35529b44c957737bf422127283c08e['h0201a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0100e] =  Ifd35529b44c957737bf422127283c08e['h0201c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0100f] =  Ifd35529b44c957737bf422127283c08e['h0201e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01010] =  Ifd35529b44c957737bf422127283c08e['h02020] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01011] =  Ifd35529b44c957737bf422127283c08e['h02022] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01012] =  Ifd35529b44c957737bf422127283c08e['h02024] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01013] =  Ifd35529b44c957737bf422127283c08e['h02026] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01014] =  Ifd35529b44c957737bf422127283c08e['h02028] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01015] =  Ifd35529b44c957737bf422127283c08e['h0202a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01016] =  Ifd35529b44c957737bf422127283c08e['h0202c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01017] =  Ifd35529b44c957737bf422127283c08e['h0202e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01018] =  Ifd35529b44c957737bf422127283c08e['h02030] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01019] =  Ifd35529b44c957737bf422127283c08e['h02032] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0101a] =  Ifd35529b44c957737bf422127283c08e['h02034] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0101b] =  Ifd35529b44c957737bf422127283c08e['h02036] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0101c] =  Ifd35529b44c957737bf422127283c08e['h02038] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0101d] =  Ifd35529b44c957737bf422127283c08e['h0203a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0101e] =  Ifd35529b44c957737bf422127283c08e['h0203c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0101f] =  Ifd35529b44c957737bf422127283c08e['h0203e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01020] =  Ifd35529b44c957737bf422127283c08e['h02040] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01021] =  Ifd35529b44c957737bf422127283c08e['h02042] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01022] =  Ifd35529b44c957737bf422127283c08e['h02044] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01023] =  Ifd35529b44c957737bf422127283c08e['h02046] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01024] =  Ifd35529b44c957737bf422127283c08e['h02048] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01025] =  Ifd35529b44c957737bf422127283c08e['h0204a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01026] =  Ifd35529b44c957737bf422127283c08e['h0204c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01027] =  Ifd35529b44c957737bf422127283c08e['h0204e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01028] =  Ifd35529b44c957737bf422127283c08e['h02050] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01029] =  Ifd35529b44c957737bf422127283c08e['h02052] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0102a] =  Ifd35529b44c957737bf422127283c08e['h02054] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0102b] =  Ifd35529b44c957737bf422127283c08e['h02056] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0102c] =  Ifd35529b44c957737bf422127283c08e['h02058] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0102d] =  Ifd35529b44c957737bf422127283c08e['h0205a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0102e] =  Ifd35529b44c957737bf422127283c08e['h0205c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0102f] =  Ifd35529b44c957737bf422127283c08e['h0205e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01030] =  Ifd35529b44c957737bf422127283c08e['h02060] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01031] =  Ifd35529b44c957737bf422127283c08e['h02062] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01032] =  Ifd35529b44c957737bf422127283c08e['h02064] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01033] =  Ifd35529b44c957737bf422127283c08e['h02066] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01034] =  Ifd35529b44c957737bf422127283c08e['h02068] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01035] =  Ifd35529b44c957737bf422127283c08e['h0206a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01036] =  Ifd35529b44c957737bf422127283c08e['h0206c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01037] =  Ifd35529b44c957737bf422127283c08e['h0206e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01038] =  Ifd35529b44c957737bf422127283c08e['h02070] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01039] =  Ifd35529b44c957737bf422127283c08e['h02072] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0103a] =  Ifd35529b44c957737bf422127283c08e['h02074] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0103b] =  Ifd35529b44c957737bf422127283c08e['h02076] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0103c] =  Ifd35529b44c957737bf422127283c08e['h02078] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0103d] =  Ifd35529b44c957737bf422127283c08e['h0207a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0103e] =  Ifd35529b44c957737bf422127283c08e['h0207c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0103f] =  Ifd35529b44c957737bf422127283c08e['h0207e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01040] =  Ifd35529b44c957737bf422127283c08e['h02080] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01041] =  Ifd35529b44c957737bf422127283c08e['h02082] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01042] =  Ifd35529b44c957737bf422127283c08e['h02084] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01043] =  Ifd35529b44c957737bf422127283c08e['h02086] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01044] =  Ifd35529b44c957737bf422127283c08e['h02088] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01045] =  Ifd35529b44c957737bf422127283c08e['h0208a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01046] =  Ifd35529b44c957737bf422127283c08e['h0208c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01047] =  Ifd35529b44c957737bf422127283c08e['h0208e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01048] =  Ifd35529b44c957737bf422127283c08e['h02090] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01049] =  Ifd35529b44c957737bf422127283c08e['h02092] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0104a] =  Ifd35529b44c957737bf422127283c08e['h02094] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0104b] =  Ifd35529b44c957737bf422127283c08e['h02096] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0104c] =  Ifd35529b44c957737bf422127283c08e['h02098] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0104d] =  Ifd35529b44c957737bf422127283c08e['h0209a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0104e] =  Ifd35529b44c957737bf422127283c08e['h0209c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0104f] =  Ifd35529b44c957737bf422127283c08e['h0209e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01050] =  Ifd35529b44c957737bf422127283c08e['h020a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01051] =  Ifd35529b44c957737bf422127283c08e['h020a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01052] =  Ifd35529b44c957737bf422127283c08e['h020a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01053] =  Ifd35529b44c957737bf422127283c08e['h020a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01054] =  Ifd35529b44c957737bf422127283c08e['h020a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01055] =  Ifd35529b44c957737bf422127283c08e['h020aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01056] =  Ifd35529b44c957737bf422127283c08e['h020ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01057] =  Ifd35529b44c957737bf422127283c08e['h020ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01058] =  Ifd35529b44c957737bf422127283c08e['h020b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01059] =  Ifd35529b44c957737bf422127283c08e['h020b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0105a] =  Ifd35529b44c957737bf422127283c08e['h020b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0105b] =  Ifd35529b44c957737bf422127283c08e['h020b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0105c] =  Ifd35529b44c957737bf422127283c08e['h020b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0105d] =  Ifd35529b44c957737bf422127283c08e['h020ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0105e] =  Ifd35529b44c957737bf422127283c08e['h020bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0105f] =  Ifd35529b44c957737bf422127283c08e['h020be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01060] =  Ifd35529b44c957737bf422127283c08e['h020c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01061] =  Ifd35529b44c957737bf422127283c08e['h020c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01062] =  Ifd35529b44c957737bf422127283c08e['h020c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01063] =  Ifd35529b44c957737bf422127283c08e['h020c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01064] =  Ifd35529b44c957737bf422127283c08e['h020c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01065] =  Ifd35529b44c957737bf422127283c08e['h020ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01066] =  Ifd35529b44c957737bf422127283c08e['h020cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01067] =  Ifd35529b44c957737bf422127283c08e['h020ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01068] =  Ifd35529b44c957737bf422127283c08e['h020d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01069] =  Ifd35529b44c957737bf422127283c08e['h020d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0106a] =  Ifd35529b44c957737bf422127283c08e['h020d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0106b] =  Ifd35529b44c957737bf422127283c08e['h020d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0106c] =  Ifd35529b44c957737bf422127283c08e['h020d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0106d] =  Ifd35529b44c957737bf422127283c08e['h020da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0106e] =  Ifd35529b44c957737bf422127283c08e['h020dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0106f] =  Ifd35529b44c957737bf422127283c08e['h020de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01070] =  Ifd35529b44c957737bf422127283c08e['h020e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01071] =  Ifd35529b44c957737bf422127283c08e['h020e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01072] =  Ifd35529b44c957737bf422127283c08e['h020e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01073] =  Ifd35529b44c957737bf422127283c08e['h020e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01074] =  Ifd35529b44c957737bf422127283c08e['h020e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01075] =  Ifd35529b44c957737bf422127283c08e['h020ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01076] =  Ifd35529b44c957737bf422127283c08e['h020ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01077] =  Ifd35529b44c957737bf422127283c08e['h020ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01078] =  Ifd35529b44c957737bf422127283c08e['h020f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01079] =  Ifd35529b44c957737bf422127283c08e['h020f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0107a] =  Ifd35529b44c957737bf422127283c08e['h020f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0107b] =  Ifd35529b44c957737bf422127283c08e['h020f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0107c] =  Ifd35529b44c957737bf422127283c08e['h020f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0107d] =  Ifd35529b44c957737bf422127283c08e['h020fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0107e] =  Ifd35529b44c957737bf422127283c08e['h020fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0107f] =  Ifd35529b44c957737bf422127283c08e['h020fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01080] =  Ifd35529b44c957737bf422127283c08e['h02100] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01081] =  Ifd35529b44c957737bf422127283c08e['h02102] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01082] =  Ifd35529b44c957737bf422127283c08e['h02104] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01083] =  Ifd35529b44c957737bf422127283c08e['h02106] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01084] =  Ifd35529b44c957737bf422127283c08e['h02108] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01085] =  Ifd35529b44c957737bf422127283c08e['h0210a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01086] =  Ifd35529b44c957737bf422127283c08e['h0210c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01087] =  Ifd35529b44c957737bf422127283c08e['h0210e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01088] =  Ifd35529b44c957737bf422127283c08e['h02110] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01089] =  Ifd35529b44c957737bf422127283c08e['h02112] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0108a] =  Ifd35529b44c957737bf422127283c08e['h02114] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0108b] =  Ifd35529b44c957737bf422127283c08e['h02116] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0108c] =  Ifd35529b44c957737bf422127283c08e['h02118] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0108d] =  Ifd35529b44c957737bf422127283c08e['h0211a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0108e] =  Ifd35529b44c957737bf422127283c08e['h0211c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0108f] =  Ifd35529b44c957737bf422127283c08e['h0211e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01090] =  Ifd35529b44c957737bf422127283c08e['h02120] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01091] =  Ifd35529b44c957737bf422127283c08e['h02122] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01092] =  Ifd35529b44c957737bf422127283c08e['h02124] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01093] =  Ifd35529b44c957737bf422127283c08e['h02126] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01094] =  Ifd35529b44c957737bf422127283c08e['h02128] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01095] =  Ifd35529b44c957737bf422127283c08e['h0212a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01096] =  Ifd35529b44c957737bf422127283c08e['h0212c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01097] =  Ifd35529b44c957737bf422127283c08e['h0212e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01098] =  Ifd35529b44c957737bf422127283c08e['h02130] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01099] =  Ifd35529b44c957737bf422127283c08e['h02132] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0109a] =  Ifd35529b44c957737bf422127283c08e['h02134] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0109b] =  Ifd35529b44c957737bf422127283c08e['h02136] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0109c] =  Ifd35529b44c957737bf422127283c08e['h02138] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0109d] =  Ifd35529b44c957737bf422127283c08e['h0213a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0109e] =  Ifd35529b44c957737bf422127283c08e['h0213c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0109f] =  Ifd35529b44c957737bf422127283c08e['h0213e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010a0] =  Ifd35529b44c957737bf422127283c08e['h02140] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010a1] =  Ifd35529b44c957737bf422127283c08e['h02142] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010a2] =  Ifd35529b44c957737bf422127283c08e['h02144] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010a3] =  Ifd35529b44c957737bf422127283c08e['h02146] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010a4] =  Ifd35529b44c957737bf422127283c08e['h02148] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010a5] =  Ifd35529b44c957737bf422127283c08e['h0214a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010a6] =  Ifd35529b44c957737bf422127283c08e['h0214c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010a7] =  Ifd35529b44c957737bf422127283c08e['h0214e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010a8] =  Ifd35529b44c957737bf422127283c08e['h02150] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010a9] =  Ifd35529b44c957737bf422127283c08e['h02152] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010aa] =  Ifd35529b44c957737bf422127283c08e['h02154] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010ab] =  Ifd35529b44c957737bf422127283c08e['h02156] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010ac] =  Ifd35529b44c957737bf422127283c08e['h02158] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010ad] =  Ifd35529b44c957737bf422127283c08e['h0215a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010ae] =  Ifd35529b44c957737bf422127283c08e['h0215c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010af] =  Ifd35529b44c957737bf422127283c08e['h0215e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010b0] =  Ifd35529b44c957737bf422127283c08e['h02160] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010b1] =  Ifd35529b44c957737bf422127283c08e['h02162] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010b2] =  Ifd35529b44c957737bf422127283c08e['h02164] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010b3] =  Ifd35529b44c957737bf422127283c08e['h02166] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010b4] =  Ifd35529b44c957737bf422127283c08e['h02168] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010b5] =  Ifd35529b44c957737bf422127283c08e['h0216a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010b6] =  Ifd35529b44c957737bf422127283c08e['h0216c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010b7] =  Ifd35529b44c957737bf422127283c08e['h0216e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010b8] =  Ifd35529b44c957737bf422127283c08e['h02170] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010b9] =  Ifd35529b44c957737bf422127283c08e['h02172] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010ba] =  Ifd35529b44c957737bf422127283c08e['h02174] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010bb] =  Ifd35529b44c957737bf422127283c08e['h02176] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010bc] =  Ifd35529b44c957737bf422127283c08e['h02178] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010bd] =  Ifd35529b44c957737bf422127283c08e['h0217a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010be] =  Ifd35529b44c957737bf422127283c08e['h0217c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010bf] =  Ifd35529b44c957737bf422127283c08e['h0217e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010c0] =  Ifd35529b44c957737bf422127283c08e['h02180] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010c1] =  Ifd35529b44c957737bf422127283c08e['h02182] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010c2] =  Ifd35529b44c957737bf422127283c08e['h02184] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010c3] =  Ifd35529b44c957737bf422127283c08e['h02186] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010c4] =  Ifd35529b44c957737bf422127283c08e['h02188] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010c5] =  Ifd35529b44c957737bf422127283c08e['h0218a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010c6] =  Ifd35529b44c957737bf422127283c08e['h0218c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010c7] =  Ifd35529b44c957737bf422127283c08e['h0218e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010c8] =  Ifd35529b44c957737bf422127283c08e['h02190] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010c9] =  Ifd35529b44c957737bf422127283c08e['h02192] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010ca] =  Ifd35529b44c957737bf422127283c08e['h02194] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010cb] =  Ifd35529b44c957737bf422127283c08e['h02196] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010cc] =  Ifd35529b44c957737bf422127283c08e['h02198] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010cd] =  Ifd35529b44c957737bf422127283c08e['h0219a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010ce] =  Ifd35529b44c957737bf422127283c08e['h0219c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010cf] =  Ifd35529b44c957737bf422127283c08e['h0219e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010d0] =  Ifd35529b44c957737bf422127283c08e['h021a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010d1] =  Ifd35529b44c957737bf422127283c08e['h021a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010d2] =  Ifd35529b44c957737bf422127283c08e['h021a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010d3] =  Ifd35529b44c957737bf422127283c08e['h021a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010d4] =  Ifd35529b44c957737bf422127283c08e['h021a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010d5] =  Ifd35529b44c957737bf422127283c08e['h021aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010d6] =  Ifd35529b44c957737bf422127283c08e['h021ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010d7] =  Ifd35529b44c957737bf422127283c08e['h021ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010d8] =  Ifd35529b44c957737bf422127283c08e['h021b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010d9] =  Ifd35529b44c957737bf422127283c08e['h021b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010da] =  Ifd35529b44c957737bf422127283c08e['h021b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010db] =  Ifd35529b44c957737bf422127283c08e['h021b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010dc] =  Ifd35529b44c957737bf422127283c08e['h021b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010dd] =  Ifd35529b44c957737bf422127283c08e['h021ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010de] =  Ifd35529b44c957737bf422127283c08e['h021bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010df] =  Ifd35529b44c957737bf422127283c08e['h021be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010e0] =  Ifd35529b44c957737bf422127283c08e['h021c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010e1] =  Ifd35529b44c957737bf422127283c08e['h021c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010e2] =  Ifd35529b44c957737bf422127283c08e['h021c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010e3] =  Ifd35529b44c957737bf422127283c08e['h021c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010e4] =  Ifd35529b44c957737bf422127283c08e['h021c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010e5] =  Ifd35529b44c957737bf422127283c08e['h021ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010e6] =  Ifd35529b44c957737bf422127283c08e['h021cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010e7] =  Ifd35529b44c957737bf422127283c08e['h021ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010e8] =  Ifd35529b44c957737bf422127283c08e['h021d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010e9] =  Ifd35529b44c957737bf422127283c08e['h021d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010ea] =  Ifd35529b44c957737bf422127283c08e['h021d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010eb] =  Ifd35529b44c957737bf422127283c08e['h021d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010ec] =  Ifd35529b44c957737bf422127283c08e['h021d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010ed] =  Ifd35529b44c957737bf422127283c08e['h021da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010ee] =  Ifd35529b44c957737bf422127283c08e['h021dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010ef] =  Ifd35529b44c957737bf422127283c08e['h021de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010f0] =  Ifd35529b44c957737bf422127283c08e['h021e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010f1] =  Ifd35529b44c957737bf422127283c08e['h021e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010f2] =  Ifd35529b44c957737bf422127283c08e['h021e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010f3] =  Ifd35529b44c957737bf422127283c08e['h021e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010f4] =  Ifd35529b44c957737bf422127283c08e['h021e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010f5] =  Ifd35529b44c957737bf422127283c08e['h021ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010f6] =  Ifd35529b44c957737bf422127283c08e['h021ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010f7] =  Ifd35529b44c957737bf422127283c08e['h021ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010f8] =  Ifd35529b44c957737bf422127283c08e['h021f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010f9] =  Ifd35529b44c957737bf422127283c08e['h021f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010fa] =  Ifd35529b44c957737bf422127283c08e['h021f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010fb] =  Ifd35529b44c957737bf422127283c08e['h021f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010fc] =  Ifd35529b44c957737bf422127283c08e['h021f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010fd] =  Ifd35529b44c957737bf422127283c08e['h021fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010fe] =  Ifd35529b44c957737bf422127283c08e['h021fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h010ff] =  Ifd35529b44c957737bf422127283c08e['h021fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01100] =  Ifd35529b44c957737bf422127283c08e['h02200] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01101] =  Ifd35529b44c957737bf422127283c08e['h02202] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01102] =  Ifd35529b44c957737bf422127283c08e['h02204] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01103] =  Ifd35529b44c957737bf422127283c08e['h02206] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01104] =  Ifd35529b44c957737bf422127283c08e['h02208] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01105] =  Ifd35529b44c957737bf422127283c08e['h0220a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01106] =  Ifd35529b44c957737bf422127283c08e['h0220c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01107] =  Ifd35529b44c957737bf422127283c08e['h0220e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01108] =  Ifd35529b44c957737bf422127283c08e['h02210] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01109] =  Ifd35529b44c957737bf422127283c08e['h02212] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0110a] =  Ifd35529b44c957737bf422127283c08e['h02214] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0110b] =  Ifd35529b44c957737bf422127283c08e['h02216] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0110c] =  Ifd35529b44c957737bf422127283c08e['h02218] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0110d] =  Ifd35529b44c957737bf422127283c08e['h0221a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0110e] =  Ifd35529b44c957737bf422127283c08e['h0221c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0110f] =  Ifd35529b44c957737bf422127283c08e['h0221e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01110] =  Ifd35529b44c957737bf422127283c08e['h02220] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01111] =  Ifd35529b44c957737bf422127283c08e['h02222] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01112] =  Ifd35529b44c957737bf422127283c08e['h02224] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01113] =  Ifd35529b44c957737bf422127283c08e['h02226] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01114] =  Ifd35529b44c957737bf422127283c08e['h02228] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01115] =  Ifd35529b44c957737bf422127283c08e['h0222a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01116] =  Ifd35529b44c957737bf422127283c08e['h0222c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01117] =  Ifd35529b44c957737bf422127283c08e['h0222e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01118] =  Ifd35529b44c957737bf422127283c08e['h02230] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01119] =  Ifd35529b44c957737bf422127283c08e['h02232] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0111a] =  Ifd35529b44c957737bf422127283c08e['h02234] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0111b] =  Ifd35529b44c957737bf422127283c08e['h02236] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0111c] =  Ifd35529b44c957737bf422127283c08e['h02238] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0111d] =  Ifd35529b44c957737bf422127283c08e['h0223a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0111e] =  Ifd35529b44c957737bf422127283c08e['h0223c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0111f] =  Ifd35529b44c957737bf422127283c08e['h0223e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01120] =  Ifd35529b44c957737bf422127283c08e['h02240] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01121] =  Ifd35529b44c957737bf422127283c08e['h02242] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01122] =  Ifd35529b44c957737bf422127283c08e['h02244] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01123] =  Ifd35529b44c957737bf422127283c08e['h02246] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01124] =  Ifd35529b44c957737bf422127283c08e['h02248] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01125] =  Ifd35529b44c957737bf422127283c08e['h0224a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01126] =  Ifd35529b44c957737bf422127283c08e['h0224c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01127] =  Ifd35529b44c957737bf422127283c08e['h0224e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01128] =  Ifd35529b44c957737bf422127283c08e['h02250] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01129] =  Ifd35529b44c957737bf422127283c08e['h02252] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0112a] =  Ifd35529b44c957737bf422127283c08e['h02254] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0112b] =  Ifd35529b44c957737bf422127283c08e['h02256] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0112c] =  Ifd35529b44c957737bf422127283c08e['h02258] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0112d] =  Ifd35529b44c957737bf422127283c08e['h0225a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0112e] =  Ifd35529b44c957737bf422127283c08e['h0225c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0112f] =  Ifd35529b44c957737bf422127283c08e['h0225e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01130] =  Ifd35529b44c957737bf422127283c08e['h02260] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01131] =  Ifd35529b44c957737bf422127283c08e['h02262] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01132] =  Ifd35529b44c957737bf422127283c08e['h02264] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01133] =  Ifd35529b44c957737bf422127283c08e['h02266] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01134] =  Ifd35529b44c957737bf422127283c08e['h02268] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01135] =  Ifd35529b44c957737bf422127283c08e['h0226a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01136] =  Ifd35529b44c957737bf422127283c08e['h0226c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01137] =  Ifd35529b44c957737bf422127283c08e['h0226e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01138] =  Ifd35529b44c957737bf422127283c08e['h02270] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01139] =  Ifd35529b44c957737bf422127283c08e['h02272] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0113a] =  Ifd35529b44c957737bf422127283c08e['h02274] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0113b] =  Ifd35529b44c957737bf422127283c08e['h02276] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0113c] =  Ifd35529b44c957737bf422127283c08e['h02278] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0113d] =  Ifd35529b44c957737bf422127283c08e['h0227a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0113e] =  Ifd35529b44c957737bf422127283c08e['h0227c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0113f] =  Ifd35529b44c957737bf422127283c08e['h0227e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01140] =  Ifd35529b44c957737bf422127283c08e['h02280] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01141] =  Ifd35529b44c957737bf422127283c08e['h02282] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01142] =  Ifd35529b44c957737bf422127283c08e['h02284] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01143] =  Ifd35529b44c957737bf422127283c08e['h02286] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01144] =  Ifd35529b44c957737bf422127283c08e['h02288] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01145] =  Ifd35529b44c957737bf422127283c08e['h0228a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01146] =  Ifd35529b44c957737bf422127283c08e['h0228c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01147] =  Ifd35529b44c957737bf422127283c08e['h0228e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01148] =  Ifd35529b44c957737bf422127283c08e['h02290] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01149] =  Ifd35529b44c957737bf422127283c08e['h02292] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0114a] =  Ifd35529b44c957737bf422127283c08e['h02294] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0114b] =  Ifd35529b44c957737bf422127283c08e['h02296] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0114c] =  Ifd35529b44c957737bf422127283c08e['h02298] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0114d] =  Ifd35529b44c957737bf422127283c08e['h0229a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0114e] =  Ifd35529b44c957737bf422127283c08e['h0229c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0114f] =  Ifd35529b44c957737bf422127283c08e['h0229e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01150] =  Ifd35529b44c957737bf422127283c08e['h022a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01151] =  Ifd35529b44c957737bf422127283c08e['h022a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01152] =  Ifd35529b44c957737bf422127283c08e['h022a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01153] =  Ifd35529b44c957737bf422127283c08e['h022a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01154] =  Ifd35529b44c957737bf422127283c08e['h022a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01155] =  Ifd35529b44c957737bf422127283c08e['h022aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01156] =  Ifd35529b44c957737bf422127283c08e['h022ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01157] =  Ifd35529b44c957737bf422127283c08e['h022ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01158] =  Ifd35529b44c957737bf422127283c08e['h022b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01159] =  Ifd35529b44c957737bf422127283c08e['h022b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0115a] =  Ifd35529b44c957737bf422127283c08e['h022b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0115b] =  Ifd35529b44c957737bf422127283c08e['h022b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0115c] =  Ifd35529b44c957737bf422127283c08e['h022b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0115d] =  Ifd35529b44c957737bf422127283c08e['h022ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0115e] =  Ifd35529b44c957737bf422127283c08e['h022bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0115f] =  Ifd35529b44c957737bf422127283c08e['h022be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01160] =  Ifd35529b44c957737bf422127283c08e['h022c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01161] =  Ifd35529b44c957737bf422127283c08e['h022c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01162] =  Ifd35529b44c957737bf422127283c08e['h022c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01163] =  Ifd35529b44c957737bf422127283c08e['h022c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01164] =  Ifd35529b44c957737bf422127283c08e['h022c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01165] =  Ifd35529b44c957737bf422127283c08e['h022ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01166] =  Ifd35529b44c957737bf422127283c08e['h022cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01167] =  Ifd35529b44c957737bf422127283c08e['h022ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01168] =  Ifd35529b44c957737bf422127283c08e['h022d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01169] =  Ifd35529b44c957737bf422127283c08e['h022d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0116a] =  Ifd35529b44c957737bf422127283c08e['h022d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0116b] =  Ifd35529b44c957737bf422127283c08e['h022d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0116c] =  Ifd35529b44c957737bf422127283c08e['h022d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0116d] =  Ifd35529b44c957737bf422127283c08e['h022da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0116e] =  Ifd35529b44c957737bf422127283c08e['h022dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0116f] =  Ifd35529b44c957737bf422127283c08e['h022de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01170] =  Ifd35529b44c957737bf422127283c08e['h022e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01171] =  Ifd35529b44c957737bf422127283c08e['h022e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01172] =  Ifd35529b44c957737bf422127283c08e['h022e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01173] =  Ifd35529b44c957737bf422127283c08e['h022e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01174] =  Ifd35529b44c957737bf422127283c08e['h022e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01175] =  Ifd35529b44c957737bf422127283c08e['h022ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01176] =  Ifd35529b44c957737bf422127283c08e['h022ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01177] =  Ifd35529b44c957737bf422127283c08e['h022ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01178] =  Ifd35529b44c957737bf422127283c08e['h022f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01179] =  Ifd35529b44c957737bf422127283c08e['h022f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0117a] =  Ifd35529b44c957737bf422127283c08e['h022f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0117b] =  Ifd35529b44c957737bf422127283c08e['h022f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0117c] =  Ifd35529b44c957737bf422127283c08e['h022f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0117d] =  Ifd35529b44c957737bf422127283c08e['h022fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0117e] =  Ifd35529b44c957737bf422127283c08e['h022fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0117f] =  Ifd35529b44c957737bf422127283c08e['h022fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01180] =  Ifd35529b44c957737bf422127283c08e['h02300] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01181] =  Ifd35529b44c957737bf422127283c08e['h02302] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01182] =  Ifd35529b44c957737bf422127283c08e['h02304] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01183] =  Ifd35529b44c957737bf422127283c08e['h02306] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01184] =  Ifd35529b44c957737bf422127283c08e['h02308] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01185] =  Ifd35529b44c957737bf422127283c08e['h0230a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01186] =  Ifd35529b44c957737bf422127283c08e['h0230c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01187] =  Ifd35529b44c957737bf422127283c08e['h0230e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01188] =  Ifd35529b44c957737bf422127283c08e['h02310] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01189] =  Ifd35529b44c957737bf422127283c08e['h02312] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0118a] =  Ifd35529b44c957737bf422127283c08e['h02314] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0118b] =  Ifd35529b44c957737bf422127283c08e['h02316] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0118c] =  Ifd35529b44c957737bf422127283c08e['h02318] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0118d] =  Ifd35529b44c957737bf422127283c08e['h0231a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0118e] =  Ifd35529b44c957737bf422127283c08e['h0231c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0118f] =  Ifd35529b44c957737bf422127283c08e['h0231e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01190] =  Ifd35529b44c957737bf422127283c08e['h02320] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01191] =  Ifd35529b44c957737bf422127283c08e['h02322] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01192] =  Ifd35529b44c957737bf422127283c08e['h02324] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01193] =  Ifd35529b44c957737bf422127283c08e['h02326] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01194] =  Ifd35529b44c957737bf422127283c08e['h02328] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01195] =  Ifd35529b44c957737bf422127283c08e['h0232a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01196] =  Ifd35529b44c957737bf422127283c08e['h0232c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01197] =  Ifd35529b44c957737bf422127283c08e['h0232e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01198] =  Ifd35529b44c957737bf422127283c08e['h02330] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01199] =  Ifd35529b44c957737bf422127283c08e['h02332] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0119a] =  Ifd35529b44c957737bf422127283c08e['h02334] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0119b] =  Ifd35529b44c957737bf422127283c08e['h02336] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0119c] =  Ifd35529b44c957737bf422127283c08e['h02338] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0119d] =  Ifd35529b44c957737bf422127283c08e['h0233a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0119e] =  Ifd35529b44c957737bf422127283c08e['h0233c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0119f] =  Ifd35529b44c957737bf422127283c08e['h0233e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011a0] =  Ifd35529b44c957737bf422127283c08e['h02340] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011a1] =  Ifd35529b44c957737bf422127283c08e['h02342] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011a2] =  Ifd35529b44c957737bf422127283c08e['h02344] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011a3] =  Ifd35529b44c957737bf422127283c08e['h02346] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011a4] =  Ifd35529b44c957737bf422127283c08e['h02348] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011a5] =  Ifd35529b44c957737bf422127283c08e['h0234a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011a6] =  Ifd35529b44c957737bf422127283c08e['h0234c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011a7] =  Ifd35529b44c957737bf422127283c08e['h0234e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011a8] =  Ifd35529b44c957737bf422127283c08e['h02350] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011a9] =  Ifd35529b44c957737bf422127283c08e['h02352] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011aa] =  Ifd35529b44c957737bf422127283c08e['h02354] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011ab] =  Ifd35529b44c957737bf422127283c08e['h02356] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011ac] =  Ifd35529b44c957737bf422127283c08e['h02358] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011ad] =  Ifd35529b44c957737bf422127283c08e['h0235a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011ae] =  Ifd35529b44c957737bf422127283c08e['h0235c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011af] =  Ifd35529b44c957737bf422127283c08e['h0235e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011b0] =  Ifd35529b44c957737bf422127283c08e['h02360] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011b1] =  Ifd35529b44c957737bf422127283c08e['h02362] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011b2] =  Ifd35529b44c957737bf422127283c08e['h02364] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011b3] =  Ifd35529b44c957737bf422127283c08e['h02366] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011b4] =  Ifd35529b44c957737bf422127283c08e['h02368] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011b5] =  Ifd35529b44c957737bf422127283c08e['h0236a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011b6] =  Ifd35529b44c957737bf422127283c08e['h0236c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011b7] =  Ifd35529b44c957737bf422127283c08e['h0236e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011b8] =  Ifd35529b44c957737bf422127283c08e['h02370] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011b9] =  Ifd35529b44c957737bf422127283c08e['h02372] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011ba] =  Ifd35529b44c957737bf422127283c08e['h02374] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011bb] =  Ifd35529b44c957737bf422127283c08e['h02376] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011bc] =  Ifd35529b44c957737bf422127283c08e['h02378] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011bd] =  Ifd35529b44c957737bf422127283c08e['h0237a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011be] =  Ifd35529b44c957737bf422127283c08e['h0237c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011bf] =  Ifd35529b44c957737bf422127283c08e['h0237e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011c0] =  Ifd35529b44c957737bf422127283c08e['h02380] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011c1] =  Ifd35529b44c957737bf422127283c08e['h02382] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011c2] =  Ifd35529b44c957737bf422127283c08e['h02384] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011c3] =  Ifd35529b44c957737bf422127283c08e['h02386] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011c4] =  Ifd35529b44c957737bf422127283c08e['h02388] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011c5] =  Ifd35529b44c957737bf422127283c08e['h0238a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011c6] =  Ifd35529b44c957737bf422127283c08e['h0238c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011c7] =  Ifd35529b44c957737bf422127283c08e['h0238e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011c8] =  Ifd35529b44c957737bf422127283c08e['h02390] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011c9] =  Ifd35529b44c957737bf422127283c08e['h02392] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011ca] =  Ifd35529b44c957737bf422127283c08e['h02394] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011cb] =  Ifd35529b44c957737bf422127283c08e['h02396] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011cc] =  Ifd35529b44c957737bf422127283c08e['h02398] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011cd] =  Ifd35529b44c957737bf422127283c08e['h0239a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011ce] =  Ifd35529b44c957737bf422127283c08e['h0239c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011cf] =  Ifd35529b44c957737bf422127283c08e['h0239e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011d0] =  Ifd35529b44c957737bf422127283c08e['h023a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011d1] =  Ifd35529b44c957737bf422127283c08e['h023a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011d2] =  Ifd35529b44c957737bf422127283c08e['h023a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011d3] =  Ifd35529b44c957737bf422127283c08e['h023a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011d4] =  Ifd35529b44c957737bf422127283c08e['h023a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011d5] =  Ifd35529b44c957737bf422127283c08e['h023aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011d6] =  Ifd35529b44c957737bf422127283c08e['h023ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011d7] =  Ifd35529b44c957737bf422127283c08e['h023ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011d8] =  Ifd35529b44c957737bf422127283c08e['h023b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011d9] =  Ifd35529b44c957737bf422127283c08e['h023b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011da] =  Ifd35529b44c957737bf422127283c08e['h023b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011db] =  Ifd35529b44c957737bf422127283c08e['h023b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011dc] =  Ifd35529b44c957737bf422127283c08e['h023b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011dd] =  Ifd35529b44c957737bf422127283c08e['h023ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011de] =  Ifd35529b44c957737bf422127283c08e['h023bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011df] =  Ifd35529b44c957737bf422127283c08e['h023be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011e0] =  Ifd35529b44c957737bf422127283c08e['h023c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011e1] =  Ifd35529b44c957737bf422127283c08e['h023c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011e2] =  Ifd35529b44c957737bf422127283c08e['h023c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011e3] =  Ifd35529b44c957737bf422127283c08e['h023c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011e4] =  Ifd35529b44c957737bf422127283c08e['h023c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011e5] =  Ifd35529b44c957737bf422127283c08e['h023ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011e6] =  Ifd35529b44c957737bf422127283c08e['h023cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011e7] =  Ifd35529b44c957737bf422127283c08e['h023ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011e8] =  Ifd35529b44c957737bf422127283c08e['h023d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011e9] =  Ifd35529b44c957737bf422127283c08e['h023d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011ea] =  Ifd35529b44c957737bf422127283c08e['h023d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011eb] =  Ifd35529b44c957737bf422127283c08e['h023d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011ec] =  Ifd35529b44c957737bf422127283c08e['h023d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011ed] =  Ifd35529b44c957737bf422127283c08e['h023da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011ee] =  Ifd35529b44c957737bf422127283c08e['h023dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011ef] =  Ifd35529b44c957737bf422127283c08e['h023de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011f0] =  Ifd35529b44c957737bf422127283c08e['h023e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011f1] =  Ifd35529b44c957737bf422127283c08e['h023e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011f2] =  Ifd35529b44c957737bf422127283c08e['h023e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011f3] =  Ifd35529b44c957737bf422127283c08e['h023e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011f4] =  Ifd35529b44c957737bf422127283c08e['h023e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011f5] =  Ifd35529b44c957737bf422127283c08e['h023ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011f6] =  Ifd35529b44c957737bf422127283c08e['h023ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011f7] =  Ifd35529b44c957737bf422127283c08e['h023ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011f8] =  Ifd35529b44c957737bf422127283c08e['h023f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011f9] =  Ifd35529b44c957737bf422127283c08e['h023f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011fa] =  Ifd35529b44c957737bf422127283c08e['h023f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011fb] =  Ifd35529b44c957737bf422127283c08e['h023f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011fc] =  Ifd35529b44c957737bf422127283c08e['h023f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011fd] =  Ifd35529b44c957737bf422127283c08e['h023fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011fe] =  Ifd35529b44c957737bf422127283c08e['h023fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h011ff] =  Ifd35529b44c957737bf422127283c08e['h023fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01200] =  Ifd35529b44c957737bf422127283c08e['h02400] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01201] =  Ifd35529b44c957737bf422127283c08e['h02402] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01202] =  Ifd35529b44c957737bf422127283c08e['h02404] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01203] =  Ifd35529b44c957737bf422127283c08e['h02406] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01204] =  Ifd35529b44c957737bf422127283c08e['h02408] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01205] =  Ifd35529b44c957737bf422127283c08e['h0240a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01206] =  Ifd35529b44c957737bf422127283c08e['h0240c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01207] =  Ifd35529b44c957737bf422127283c08e['h0240e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01208] =  Ifd35529b44c957737bf422127283c08e['h02410] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01209] =  Ifd35529b44c957737bf422127283c08e['h02412] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0120a] =  Ifd35529b44c957737bf422127283c08e['h02414] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0120b] =  Ifd35529b44c957737bf422127283c08e['h02416] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0120c] =  Ifd35529b44c957737bf422127283c08e['h02418] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0120d] =  Ifd35529b44c957737bf422127283c08e['h0241a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0120e] =  Ifd35529b44c957737bf422127283c08e['h0241c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0120f] =  Ifd35529b44c957737bf422127283c08e['h0241e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01210] =  Ifd35529b44c957737bf422127283c08e['h02420] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01211] =  Ifd35529b44c957737bf422127283c08e['h02422] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01212] =  Ifd35529b44c957737bf422127283c08e['h02424] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01213] =  Ifd35529b44c957737bf422127283c08e['h02426] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01214] =  Ifd35529b44c957737bf422127283c08e['h02428] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01215] =  Ifd35529b44c957737bf422127283c08e['h0242a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01216] =  Ifd35529b44c957737bf422127283c08e['h0242c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01217] =  Ifd35529b44c957737bf422127283c08e['h0242e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01218] =  Ifd35529b44c957737bf422127283c08e['h02430] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01219] =  Ifd35529b44c957737bf422127283c08e['h02432] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0121a] =  Ifd35529b44c957737bf422127283c08e['h02434] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0121b] =  Ifd35529b44c957737bf422127283c08e['h02436] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0121c] =  Ifd35529b44c957737bf422127283c08e['h02438] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0121d] =  Ifd35529b44c957737bf422127283c08e['h0243a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0121e] =  Ifd35529b44c957737bf422127283c08e['h0243c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0121f] =  Ifd35529b44c957737bf422127283c08e['h0243e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01220] =  Ifd35529b44c957737bf422127283c08e['h02440] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01221] =  Ifd35529b44c957737bf422127283c08e['h02442] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01222] =  Ifd35529b44c957737bf422127283c08e['h02444] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01223] =  Ifd35529b44c957737bf422127283c08e['h02446] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01224] =  Ifd35529b44c957737bf422127283c08e['h02448] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01225] =  Ifd35529b44c957737bf422127283c08e['h0244a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01226] =  Ifd35529b44c957737bf422127283c08e['h0244c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01227] =  Ifd35529b44c957737bf422127283c08e['h0244e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01228] =  Ifd35529b44c957737bf422127283c08e['h02450] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01229] =  Ifd35529b44c957737bf422127283c08e['h02452] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0122a] =  Ifd35529b44c957737bf422127283c08e['h02454] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0122b] =  Ifd35529b44c957737bf422127283c08e['h02456] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0122c] =  Ifd35529b44c957737bf422127283c08e['h02458] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0122d] =  Ifd35529b44c957737bf422127283c08e['h0245a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0122e] =  Ifd35529b44c957737bf422127283c08e['h0245c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0122f] =  Ifd35529b44c957737bf422127283c08e['h0245e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01230] =  Ifd35529b44c957737bf422127283c08e['h02460] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01231] =  Ifd35529b44c957737bf422127283c08e['h02462] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01232] =  Ifd35529b44c957737bf422127283c08e['h02464] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01233] =  Ifd35529b44c957737bf422127283c08e['h02466] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01234] =  Ifd35529b44c957737bf422127283c08e['h02468] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01235] =  Ifd35529b44c957737bf422127283c08e['h0246a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01236] =  Ifd35529b44c957737bf422127283c08e['h0246c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01237] =  Ifd35529b44c957737bf422127283c08e['h0246e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01238] =  Ifd35529b44c957737bf422127283c08e['h02470] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01239] =  Ifd35529b44c957737bf422127283c08e['h02472] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0123a] =  Ifd35529b44c957737bf422127283c08e['h02474] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0123b] =  Ifd35529b44c957737bf422127283c08e['h02476] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0123c] =  Ifd35529b44c957737bf422127283c08e['h02478] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0123d] =  Ifd35529b44c957737bf422127283c08e['h0247a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0123e] =  Ifd35529b44c957737bf422127283c08e['h0247c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0123f] =  Ifd35529b44c957737bf422127283c08e['h0247e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01240] =  Ifd35529b44c957737bf422127283c08e['h02480] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01241] =  Ifd35529b44c957737bf422127283c08e['h02482] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01242] =  Ifd35529b44c957737bf422127283c08e['h02484] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01243] =  Ifd35529b44c957737bf422127283c08e['h02486] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01244] =  Ifd35529b44c957737bf422127283c08e['h02488] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01245] =  Ifd35529b44c957737bf422127283c08e['h0248a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01246] =  Ifd35529b44c957737bf422127283c08e['h0248c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01247] =  Ifd35529b44c957737bf422127283c08e['h0248e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01248] =  Ifd35529b44c957737bf422127283c08e['h02490] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01249] =  Ifd35529b44c957737bf422127283c08e['h02492] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0124a] =  Ifd35529b44c957737bf422127283c08e['h02494] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0124b] =  Ifd35529b44c957737bf422127283c08e['h02496] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0124c] =  Ifd35529b44c957737bf422127283c08e['h02498] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0124d] =  Ifd35529b44c957737bf422127283c08e['h0249a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0124e] =  Ifd35529b44c957737bf422127283c08e['h0249c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0124f] =  Ifd35529b44c957737bf422127283c08e['h0249e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01250] =  Ifd35529b44c957737bf422127283c08e['h024a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01251] =  Ifd35529b44c957737bf422127283c08e['h024a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01252] =  Ifd35529b44c957737bf422127283c08e['h024a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01253] =  Ifd35529b44c957737bf422127283c08e['h024a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01254] =  Ifd35529b44c957737bf422127283c08e['h024a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01255] =  Ifd35529b44c957737bf422127283c08e['h024aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01256] =  Ifd35529b44c957737bf422127283c08e['h024ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01257] =  Ifd35529b44c957737bf422127283c08e['h024ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01258] =  Ifd35529b44c957737bf422127283c08e['h024b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01259] =  Ifd35529b44c957737bf422127283c08e['h024b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0125a] =  Ifd35529b44c957737bf422127283c08e['h024b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0125b] =  Ifd35529b44c957737bf422127283c08e['h024b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0125c] =  Ifd35529b44c957737bf422127283c08e['h024b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0125d] =  Ifd35529b44c957737bf422127283c08e['h024ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0125e] =  Ifd35529b44c957737bf422127283c08e['h024bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0125f] =  Ifd35529b44c957737bf422127283c08e['h024be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01260] =  Ifd35529b44c957737bf422127283c08e['h024c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01261] =  Ifd35529b44c957737bf422127283c08e['h024c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01262] =  Ifd35529b44c957737bf422127283c08e['h024c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01263] =  Ifd35529b44c957737bf422127283c08e['h024c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01264] =  Ifd35529b44c957737bf422127283c08e['h024c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01265] =  Ifd35529b44c957737bf422127283c08e['h024ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01266] =  Ifd35529b44c957737bf422127283c08e['h024cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01267] =  Ifd35529b44c957737bf422127283c08e['h024ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01268] =  Ifd35529b44c957737bf422127283c08e['h024d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01269] =  Ifd35529b44c957737bf422127283c08e['h024d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0126a] =  Ifd35529b44c957737bf422127283c08e['h024d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0126b] =  Ifd35529b44c957737bf422127283c08e['h024d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0126c] =  Ifd35529b44c957737bf422127283c08e['h024d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0126d] =  Ifd35529b44c957737bf422127283c08e['h024da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0126e] =  Ifd35529b44c957737bf422127283c08e['h024dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0126f] =  Ifd35529b44c957737bf422127283c08e['h024de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01270] =  Ifd35529b44c957737bf422127283c08e['h024e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01271] =  Ifd35529b44c957737bf422127283c08e['h024e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01272] =  Ifd35529b44c957737bf422127283c08e['h024e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01273] =  Ifd35529b44c957737bf422127283c08e['h024e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01274] =  Ifd35529b44c957737bf422127283c08e['h024e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01275] =  Ifd35529b44c957737bf422127283c08e['h024ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01276] =  Ifd35529b44c957737bf422127283c08e['h024ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01277] =  Ifd35529b44c957737bf422127283c08e['h024ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01278] =  Ifd35529b44c957737bf422127283c08e['h024f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01279] =  Ifd35529b44c957737bf422127283c08e['h024f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0127a] =  Ifd35529b44c957737bf422127283c08e['h024f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0127b] =  Ifd35529b44c957737bf422127283c08e['h024f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0127c] =  Ifd35529b44c957737bf422127283c08e['h024f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0127d] =  Ifd35529b44c957737bf422127283c08e['h024fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0127e] =  Ifd35529b44c957737bf422127283c08e['h024fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0127f] =  Ifd35529b44c957737bf422127283c08e['h024fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01280] =  Ifd35529b44c957737bf422127283c08e['h02500] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01281] =  Ifd35529b44c957737bf422127283c08e['h02502] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01282] =  Ifd35529b44c957737bf422127283c08e['h02504] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01283] =  Ifd35529b44c957737bf422127283c08e['h02506] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01284] =  Ifd35529b44c957737bf422127283c08e['h02508] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01285] =  Ifd35529b44c957737bf422127283c08e['h0250a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01286] =  Ifd35529b44c957737bf422127283c08e['h0250c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01287] =  Ifd35529b44c957737bf422127283c08e['h0250e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01288] =  Ifd35529b44c957737bf422127283c08e['h02510] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01289] =  Ifd35529b44c957737bf422127283c08e['h02512] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0128a] =  Ifd35529b44c957737bf422127283c08e['h02514] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0128b] =  Ifd35529b44c957737bf422127283c08e['h02516] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0128c] =  Ifd35529b44c957737bf422127283c08e['h02518] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0128d] =  Ifd35529b44c957737bf422127283c08e['h0251a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0128e] =  Ifd35529b44c957737bf422127283c08e['h0251c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0128f] =  Ifd35529b44c957737bf422127283c08e['h0251e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01290] =  Ifd35529b44c957737bf422127283c08e['h02520] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01291] =  Ifd35529b44c957737bf422127283c08e['h02522] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01292] =  Ifd35529b44c957737bf422127283c08e['h02524] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01293] =  Ifd35529b44c957737bf422127283c08e['h02526] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01294] =  Ifd35529b44c957737bf422127283c08e['h02528] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01295] =  Ifd35529b44c957737bf422127283c08e['h0252a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01296] =  Ifd35529b44c957737bf422127283c08e['h0252c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01297] =  Ifd35529b44c957737bf422127283c08e['h0252e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01298] =  Ifd35529b44c957737bf422127283c08e['h02530] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01299] =  Ifd35529b44c957737bf422127283c08e['h02532] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0129a] =  Ifd35529b44c957737bf422127283c08e['h02534] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0129b] =  Ifd35529b44c957737bf422127283c08e['h02536] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0129c] =  Ifd35529b44c957737bf422127283c08e['h02538] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0129d] =  Ifd35529b44c957737bf422127283c08e['h0253a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0129e] =  Ifd35529b44c957737bf422127283c08e['h0253c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0129f] =  Ifd35529b44c957737bf422127283c08e['h0253e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012a0] =  Ifd35529b44c957737bf422127283c08e['h02540] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012a1] =  Ifd35529b44c957737bf422127283c08e['h02542] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012a2] =  Ifd35529b44c957737bf422127283c08e['h02544] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012a3] =  Ifd35529b44c957737bf422127283c08e['h02546] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012a4] =  Ifd35529b44c957737bf422127283c08e['h02548] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012a5] =  Ifd35529b44c957737bf422127283c08e['h0254a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012a6] =  Ifd35529b44c957737bf422127283c08e['h0254c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012a7] =  Ifd35529b44c957737bf422127283c08e['h0254e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012a8] =  Ifd35529b44c957737bf422127283c08e['h02550] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012a9] =  Ifd35529b44c957737bf422127283c08e['h02552] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012aa] =  Ifd35529b44c957737bf422127283c08e['h02554] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012ab] =  Ifd35529b44c957737bf422127283c08e['h02556] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012ac] =  Ifd35529b44c957737bf422127283c08e['h02558] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012ad] =  Ifd35529b44c957737bf422127283c08e['h0255a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012ae] =  Ifd35529b44c957737bf422127283c08e['h0255c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012af] =  Ifd35529b44c957737bf422127283c08e['h0255e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012b0] =  Ifd35529b44c957737bf422127283c08e['h02560] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012b1] =  Ifd35529b44c957737bf422127283c08e['h02562] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012b2] =  Ifd35529b44c957737bf422127283c08e['h02564] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012b3] =  Ifd35529b44c957737bf422127283c08e['h02566] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012b4] =  Ifd35529b44c957737bf422127283c08e['h02568] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012b5] =  Ifd35529b44c957737bf422127283c08e['h0256a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012b6] =  Ifd35529b44c957737bf422127283c08e['h0256c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012b7] =  Ifd35529b44c957737bf422127283c08e['h0256e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012b8] =  Ifd35529b44c957737bf422127283c08e['h02570] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012b9] =  Ifd35529b44c957737bf422127283c08e['h02572] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012ba] =  Ifd35529b44c957737bf422127283c08e['h02574] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012bb] =  Ifd35529b44c957737bf422127283c08e['h02576] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012bc] =  Ifd35529b44c957737bf422127283c08e['h02578] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012bd] =  Ifd35529b44c957737bf422127283c08e['h0257a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012be] =  Ifd35529b44c957737bf422127283c08e['h0257c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012bf] =  Ifd35529b44c957737bf422127283c08e['h0257e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012c0] =  Ifd35529b44c957737bf422127283c08e['h02580] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012c1] =  Ifd35529b44c957737bf422127283c08e['h02582] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012c2] =  Ifd35529b44c957737bf422127283c08e['h02584] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012c3] =  Ifd35529b44c957737bf422127283c08e['h02586] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012c4] =  Ifd35529b44c957737bf422127283c08e['h02588] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012c5] =  Ifd35529b44c957737bf422127283c08e['h0258a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012c6] =  Ifd35529b44c957737bf422127283c08e['h0258c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012c7] =  Ifd35529b44c957737bf422127283c08e['h0258e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012c8] =  Ifd35529b44c957737bf422127283c08e['h02590] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012c9] =  Ifd35529b44c957737bf422127283c08e['h02592] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012ca] =  Ifd35529b44c957737bf422127283c08e['h02594] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012cb] =  Ifd35529b44c957737bf422127283c08e['h02596] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012cc] =  Ifd35529b44c957737bf422127283c08e['h02598] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012cd] =  Ifd35529b44c957737bf422127283c08e['h0259a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012ce] =  Ifd35529b44c957737bf422127283c08e['h0259c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012cf] =  Ifd35529b44c957737bf422127283c08e['h0259e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012d0] =  Ifd35529b44c957737bf422127283c08e['h025a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012d1] =  Ifd35529b44c957737bf422127283c08e['h025a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012d2] =  Ifd35529b44c957737bf422127283c08e['h025a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012d3] =  Ifd35529b44c957737bf422127283c08e['h025a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012d4] =  Ifd35529b44c957737bf422127283c08e['h025a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012d5] =  Ifd35529b44c957737bf422127283c08e['h025aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012d6] =  Ifd35529b44c957737bf422127283c08e['h025ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012d7] =  Ifd35529b44c957737bf422127283c08e['h025ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012d8] =  Ifd35529b44c957737bf422127283c08e['h025b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012d9] =  Ifd35529b44c957737bf422127283c08e['h025b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012da] =  Ifd35529b44c957737bf422127283c08e['h025b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012db] =  Ifd35529b44c957737bf422127283c08e['h025b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012dc] =  Ifd35529b44c957737bf422127283c08e['h025b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012dd] =  Ifd35529b44c957737bf422127283c08e['h025ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012de] =  Ifd35529b44c957737bf422127283c08e['h025bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012df] =  Ifd35529b44c957737bf422127283c08e['h025be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012e0] =  Ifd35529b44c957737bf422127283c08e['h025c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012e1] =  Ifd35529b44c957737bf422127283c08e['h025c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012e2] =  Ifd35529b44c957737bf422127283c08e['h025c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012e3] =  Ifd35529b44c957737bf422127283c08e['h025c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012e4] =  Ifd35529b44c957737bf422127283c08e['h025c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012e5] =  Ifd35529b44c957737bf422127283c08e['h025ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012e6] =  Ifd35529b44c957737bf422127283c08e['h025cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012e7] =  Ifd35529b44c957737bf422127283c08e['h025ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012e8] =  Ifd35529b44c957737bf422127283c08e['h025d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012e9] =  Ifd35529b44c957737bf422127283c08e['h025d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012ea] =  Ifd35529b44c957737bf422127283c08e['h025d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012eb] =  Ifd35529b44c957737bf422127283c08e['h025d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012ec] =  Ifd35529b44c957737bf422127283c08e['h025d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012ed] =  Ifd35529b44c957737bf422127283c08e['h025da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012ee] =  Ifd35529b44c957737bf422127283c08e['h025dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012ef] =  Ifd35529b44c957737bf422127283c08e['h025de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012f0] =  Ifd35529b44c957737bf422127283c08e['h025e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012f1] =  Ifd35529b44c957737bf422127283c08e['h025e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012f2] =  Ifd35529b44c957737bf422127283c08e['h025e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012f3] =  Ifd35529b44c957737bf422127283c08e['h025e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012f4] =  Ifd35529b44c957737bf422127283c08e['h025e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012f5] =  Ifd35529b44c957737bf422127283c08e['h025ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012f6] =  Ifd35529b44c957737bf422127283c08e['h025ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012f7] =  Ifd35529b44c957737bf422127283c08e['h025ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012f8] =  Ifd35529b44c957737bf422127283c08e['h025f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012f9] =  Ifd35529b44c957737bf422127283c08e['h025f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012fa] =  Ifd35529b44c957737bf422127283c08e['h025f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012fb] =  Ifd35529b44c957737bf422127283c08e['h025f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012fc] =  Ifd35529b44c957737bf422127283c08e['h025f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012fd] =  Ifd35529b44c957737bf422127283c08e['h025fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012fe] =  Ifd35529b44c957737bf422127283c08e['h025fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h012ff] =  Ifd35529b44c957737bf422127283c08e['h025fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01300] =  Ifd35529b44c957737bf422127283c08e['h02600] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01301] =  Ifd35529b44c957737bf422127283c08e['h02602] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01302] =  Ifd35529b44c957737bf422127283c08e['h02604] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01303] =  Ifd35529b44c957737bf422127283c08e['h02606] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01304] =  Ifd35529b44c957737bf422127283c08e['h02608] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01305] =  Ifd35529b44c957737bf422127283c08e['h0260a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01306] =  Ifd35529b44c957737bf422127283c08e['h0260c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01307] =  Ifd35529b44c957737bf422127283c08e['h0260e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01308] =  Ifd35529b44c957737bf422127283c08e['h02610] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01309] =  Ifd35529b44c957737bf422127283c08e['h02612] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0130a] =  Ifd35529b44c957737bf422127283c08e['h02614] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0130b] =  Ifd35529b44c957737bf422127283c08e['h02616] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0130c] =  Ifd35529b44c957737bf422127283c08e['h02618] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0130d] =  Ifd35529b44c957737bf422127283c08e['h0261a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0130e] =  Ifd35529b44c957737bf422127283c08e['h0261c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0130f] =  Ifd35529b44c957737bf422127283c08e['h0261e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01310] =  Ifd35529b44c957737bf422127283c08e['h02620] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01311] =  Ifd35529b44c957737bf422127283c08e['h02622] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01312] =  Ifd35529b44c957737bf422127283c08e['h02624] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01313] =  Ifd35529b44c957737bf422127283c08e['h02626] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01314] =  Ifd35529b44c957737bf422127283c08e['h02628] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01315] =  Ifd35529b44c957737bf422127283c08e['h0262a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01316] =  Ifd35529b44c957737bf422127283c08e['h0262c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01317] =  Ifd35529b44c957737bf422127283c08e['h0262e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01318] =  Ifd35529b44c957737bf422127283c08e['h02630] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01319] =  Ifd35529b44c957737bf422127283c08e['h02632] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0131a] =  Ifd35529b44c957737bf422127283c08e['h02634] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0131b] =  Ifd35529b44c957737bf422127283c08e['h02636] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0131c] =  Ifd35529b44c957737bf422127283c08e['h02638] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0131d] =  Ifd35529b44c957737bf422127283c08e['h0263a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0131e] =  Ifd35529b44c957737bf422127283c08e['h0263c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0131f] =  Ifd35529b44c957737bf422127283c08e['h0263e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01320] =  Ifd35529b44c957737bf422127283c08e['h02640] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01321] =  Ifd35529b44c957737bf422127283c08e['h02642] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01322] =  Ifd35529b44c957737bf422127283c08e['h02644] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01323] =  Ifd35529b44c957737bf422127283c08e['h02646] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01324] =  Ifd35529b44c957737bf422127283c08e['h02648] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01325] =  Ifd35529b44c957737bf422127283c08e['h0264a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01326] =  Ifd35529b44c957737bf422127283c08e['h0264c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01327] =  Ifd35529b44c957737bf422127283c08e['h0264e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01328] =  Ifd35529b44c957737bf422127283c08e['h02650] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01329] =  Ifd35529b44c957737bf422127283c08e['h02652] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0132a] =  Ifd35529b44c957737bf422127283c08e['h02654] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0132b] =  Ifd35529b44c957737bf422127283c08e['h02656] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0132c] =  Ifd35529b44c957737bf422127283c08e['h02658] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0132d] =  Ifd35529b44c957737bf422127283c08e['h0265a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0132e] =  Ifd35529b44c957737bf422127283c08e['h0265c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0132f] =  Ifd35529b44c957737bf422127283c08e['h0265e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01330] =  Ifd35529b44c957737bf422127283c08e['h02660] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01331] =  Ifd35529b44c957737bf422127283c08e['h02662] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01332] =  Ifd35529b44c957737bf422127283c08e['h02664] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01333] =  Ifd35529b44c957737bf422127283c08e['h02666] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01334] =  Ifd35529b44c957737bf422127283c08e['h02668] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01335] =  Ifd35529b44c957737bf422127283c08e['h0266a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01336] =  Ifd35529b44c957737bf422127283c08e['h0266c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01337] =  Ifd35529b44c957737bf422127283c08e['h0266e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01338] =  Ifd35529b44c957737bf422127283c08e['h02670] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01339] =  Ifd35529b44c957737bf422127283c08e['h02672] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0133a] =  Ifd35529b44c957737bf422127283c08e['h02674] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0133b] =  Ifd35529b44c957737bf422127283c08e['h02676] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0133c] =  Ifd35529b44c957737bf422127283c08e['h02678] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0133d] =  Ifd35529b44c957737bf422127283c08e['h0267a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0133e] =  Ifd35529b44c957737bf422127283c08e['h0267c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0133f] =  Ifd35529b44c957737bf422127283c08e['h0267e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01340] =  Ifd35529b44c957737bf422127283c08e['h02680] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01341] =  Ifd35529b44c957737bf422127283c08e['h02682] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01342] =  Ifd35529b44c957737bf422127283c08e['h02684] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01343] =  Ifd35529b44c957737bf422127283c08e['h02686] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01344] =  Ifd35529b44c957737bf422127283c08e['h02688] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01345] =  Ifd35529b44c957737bf422127283c08e['h0268a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01346] =  Ifd35529b44c957737bf422127283c08e['h0268c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01347] =  Ifd35529b44c957737bf422127283c08e['h0268e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01348] =  Ifd35529b44c957737bf422127283c08e['h02690] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01349] =  Ifd35529b44c957737bf422127283c08e['h02692] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0134a] =  Ifd35529b44c957737bf422127283c08e['h02694] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0134b] =  Ifd35529b44c957737bf422127283c08e['h02696] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0134c] =  Ifd35529b44c957737bf422127283c08e['h02698] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0134d] =  Ifd35529b44c957737bf422127283c08e['h0269a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0134e] =  Ifd35529b44c957737bf422127283c08e['h0269c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0134f] =  Ifd35529b44c957737bf422127283c08e['h0269e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01350] =  Ifd35529b44c957737bf422127283c08e['h026a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01351] =  Ifd35529b44c957737bf422127283c08e['h026a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01352] =  Ifd35529b44c957737bf422127283c08e['h026a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01353] =  Ifd35529b44c957737bf422127283c08e['h026a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01354] =  Ifd35529b44c957737bf422127283c08e['h026a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01355] =  Ifd35529b44c957737bf422127283c08e['h026aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01356] =  Ifd35529b44c957737bf422127283c08e['h026ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01357] =  Ifd35529b44c957737bf422127283c08e['h026ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01358] =  Ifd35529b44c957737bf422127283c08e['h026b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01359] =  Ifd35529b44c957737bf422127283c08e['h026b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0135a] =  Ifd35529b44c957737bf422127283c08e['h026b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0135b] =  Ifd35529b44c957737bf422127283c08e['h026b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0135c] =  Ifd35529b44c957737bf422127283c08e['h026b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0135d] =  Ifd35529b44c957737bf422127283c08e['h026ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0135e] =  Ifd35529b44c957737bf422127283c08e['h026bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0135f] =  Ifd35529b44c957737bf422127283c08e['h026be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01360] =  Ifd35529b44c957737bf422127283c08e['h026c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01361] =  Ifd35529b44c957737bf422127283c08e['h026c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01362] =  Ifd35529b44c957737bf422127283c08e['h026c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01363] =  Ifd35529b44c957737bf422127283c08e['h026c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01364] =  Ifd35529b44c957737bf422127283c08e['h026c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01365] =  Ifd35529b44c957737bf422127283c08e['h026ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01366] =  Ifd35529b44c957737bf422127283c08e['h026cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01367] =  Ifd35529b44c957737bf422127283c08e['h026ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01368] =  Ifd35529b44c957737bf422127283c08e['h026d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01369] =  Ifd35529b44c957737bf422127283c08e['h026d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0136a] =  Ifd35529b44c957737bf422127283c08e['h026d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0136b] =  Ifd35529b44c957737bf422127283c08e['h026d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0136c] =  Ifd35529b44c957737bf422127283c08e['h026d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0136d] =  Ifd35529b44c957737bf422127283c08e['h026da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0136e] =  Ifd35529b44c957737bf422127283c08e['h026dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0136f] =  Ifd35529b44c957737bf422127283c08e['h026de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01370] =  Ifd35529b44c957737bf422127283c08e['h026e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01371] =  Ifd35529b44c957737bf422127283c08e['h026e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01372] =  Ifd35529b44c957737bf422127283c08e['h026e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01373] =  Ifd35529b44c957737bf422127283c08e['h026e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01374] =  Ifd35529b44c957737bf422127283c08e['h026e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01375] =  Ifd35529b44c957737bf422127283c08e['h026ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01376] =  Ifd35529b44c957737bf422127283c08e['h026ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01377] =  Ifd35529b44c957737bf422127283c08e['h026ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01378] =  Ifd35529b44c957737bf422127283c08e['h026f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01379] =  Ifd35529b44c957737bf422127283c08e['h026f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0137a] =  Ifd35529b44c957737bf422127283c08e['h026f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0137b] =  Ifd35529b44c957737bf422127283c08e['h026f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0137c] =  Ifd35529b44c957737bf422127283c08e['h026f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0137d] =  Ifd35529b44c957737bf422127283c08e['h026fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0137e] =  Ifd35529b44c957737bf422127283c08e['h026fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0137f] =  Ifd35529b44c957737bf422127283c08e['h026fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01380] =  Ifd35529b44c957737bf422127283c08e['h02700] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01381] =  Ifd35529b44c957737bf422127283c08e['h02702] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01382] =  Ifd35529b44c957737bf422127283c08e['h02704] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01383] =  Ifd35529b44c957737bf422127283c08e['h02706] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01384] =  Ifd35529b44c957737bf422127283c08e['h02708] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01385] =  Ifd35529b44c957737bf422127283c08e['h0270a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01386] =  Ifd35529b44c957737bf422127283c08e['h0270c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01387] =  Ifd35529b44c957737bf422127283c08e['h0270e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01388] =  Ifd35529b44c957737bf422127283c08e['h02710] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01389] =  Ifd35529b44c957737bf422127283c08e['h02712] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0138a] =  Ifd35529b44c957737bf422127283c08e['h02714] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0138b] =  Ifd35529b44c957737bf422127283c08e['h02716] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0138c] =  Ifd35529b44c957737bf422127283c08e['h02718] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0138d] =  Ifd35529b44c957737bf422127283c08e['h0271a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0138e] =  Ifd35529b44c957737bf422127283c08e['h0271c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0138f] =  Ifd35529b44c957737bf422127283c08e['h0271e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01390] =  Ifd35529b44c957737bf422127283c08e['h02720] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01391] =  Ifd35529b44c957737bf422127283c08e['h02722] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01392] =  Ifd35529b44c957737bf422127283c08e['h02724] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01393] =  Ifd35529b44c957737bf422127283c08e['h02726] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01394] =  Ifd35529b44c957737bf422127283c08e['h02728] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01395] =  Ifd35529b44c957737bf422127283c08e['h0272a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01396] =  Ifd35529b44c957737bf422127283c08e['h0272c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01397] =  Ifd35529b44c957737bf422127283c08e['h0272e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01398] =  Ifd35529b44c957737bf422127283c08e['h02730] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01399] =  Ifd35529b44c957737bf422127283c08e['h02732] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0139a] =  Ifd35529b44c957737bf422127283c08e['h02734] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0139b] =  Ifd35529b44c957737bf422127283c08e['h02736] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0139c] =  Ifd35529b44c957737bf422127283c08e['h02738] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0139d] =  Ifd35529b44c957737bf422127283c08e['h0273a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0139e] =  Ifd35529b44c957737bf422127283c08e['h0273c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0139f] =  Ifd35529b44c957737bf422127283c08e['h0273e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013a0] =  Ifd35529b44c957737bf422127283c08e['h02740] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013a1] =  Ifd35529b44c957737bf422127283c08e['h02742] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013a2] =  Ifd35529b44c957737bf422127283c08e['h02744] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013a3] =  Ifd35529b44c957737bf422127283c08e['h02746] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013a4] =  Ifd35529b44c957737bf422127283c08e['h02748] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013a5] =  Ifd35529b44c957737bf422127283c08e['h0274a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013a6] =  Ifd35529b44c957737bf422127283c08e['h0274c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013a7] =  Ifd35529b44c957737bf422127283c08e['h0274e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013a8] =  Ifd35529b44c957737bf422127283c08e['h02750] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013a9] =  Ifd35529b44c957737bf422127283c08e['h02752] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013aa] =  Ifd35529b44c957737bf422127283c08e['h02754] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013ab] =  Ifd35529b44c957737bf422127283c08e['h02756] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013ac] =  Ifd35529b44c957737bf422127283c08e['h02758] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013ad] =  Ifd35529b44c957737bf422127283c08e['h0275a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013ae] =  Ifd35529b44c957737bf422127283c08e['h0275c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013af] =  Ifd35529b44c957737bf422127283c08e['h0275e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013b0] =  Ifd35529b44c957737bf422127283c08e['h02760] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013b1] =  Ifd35529b44c957737bf422127283c08e['h02762] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013b2] =  Ifd35529b44c957737bf422127283c08e['h02764] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013b3] =  Ifd35529b44c957737bf422127283c08e['h02766] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013b4] =  Ifd35529b44c957737bf422127283c08e['h02768] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013b5] =  Ifd35529b44c957737bf422127283c08e['h0276a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013b6] =  Ifd35529b44c957737bf422127283c08e['h0276c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013b7] =  Ifd35529b44c957737bf422127283c08e['h0276e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013b8] =  Ifd35529b44c957737bf422127283c08e['h02770] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013b9] =  Ifd35529b44c957737bf422127283c08e['h02772] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013ba] =  Ifd35529b44c957737bf422127283c08e['h02774] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013bb] =  Ifd35529b44c957737bf422127283c08e['h02776] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013bc] =  Ifd35529b44c957737bf422127283c08e['h02778] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013bd] =  Ifd35529b44c957737bf422127283c08e['h0277a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013be] =  Ifd35529b44c957737bf422127283c08e['h0277c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013bf] =  Ifd35529b44c957737bf422127283c08e['h0277e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013c0] =  Ifd35529b44c957737bf422127283c08e['h02780] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013c1] =  Ifd35529b44c957737bf422127283c08e['h02782] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013c2] =  Ifd35529b44c957737bf422127283c08e['h02784] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013c3] =  Ifd35529b44c957737bf422127283c08e['h02786] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013c4] =  Ifd35529b44c957737bf422127283c08e['h02788] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013c5] =  Ifd35529b44c957737bf422127283c08e['h0278a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013c6] =  Ifd35529b44c957737bf422127283c08e['h0278c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013c7] =  Ifd35529b44c957737bf422127283c08e['h0278e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013c8] =  Ifd35529b44c957737bf422127283c08e['h02790] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013c9] =  Ifd35529b44c957737bf422127283c08e['h02792] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013ca] =  Ifd35529b44c957737bf422127283c08e['h02794] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013cb] =  Ifd35529b44c957737bf422127283c08e['h02796] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013cc] =  Ifd35529b44c957737bf422127283c08e['h02798] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013cd] =  Ifd35529b44c957737bf422127283c08e['h0279a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013ce] =  Ifd35529b44c957737bf422127283c08e['h0279c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013cf] =  Ifd35529b44c957737bf422127283c08e['h0279e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013d0] =  Ifd35529b44c957737bf422127283c08e['h027a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013d1] =  Ifd35529b44c957737bf422127283c08e['h027a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013d2] =  Ifd35529b44c957737bf422127283c08e['h027a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013d3] =  Ifd35529b44c957737bf422127283c08e['h027a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013d4] =  Ifd35529b44c957737bf422127283c08e['h027a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013d5] =  Ifd35529b44c957737bf422127283c08e['h027aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013d6] =  Ifd35529b44c957737bf422127283c08e['h027ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013d7] =  Ifd35529b44c957737bf422127283c08e['h027ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013d8] =  Ifd35529b44c957737bf422127283c08e['h027b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013d9] =  Ifd35529b44c957737bf422127283c08e['h027b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013da] =  Ifd35529b44c957737bf422127283c08e['h027b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013db] =  Ifd35529b44c957737bf422127283c08e['h027b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013dc] =  Ifd35529b44c957737bf422127283c08e['h027b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013dd] =  Ifd35529b44c957737bf422127283c08e['h027ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013de] =  Ifd35529b44c957737bf422127283c08e['h027bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013df] =  Ifd35529b44c957737bf422127283c08e['h027be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013e0] =  Ifd35529b44c957737bf422127283c08e['h027c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013e1] =  Ifd35529b44c957737bf422127283c08e['h027c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013e2] =  Ifd35529b44c957737bf422127283c08e['h027c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013e3] =  Ifd35529b44c957737bf422127283c08e['h027c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013e4] =  Ifd35529b44c957737bf422127283c08e['h027c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013e5] =  Ifd35529b44c957737bf422127283c08e['h027ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013e6] =  Ifd35529b44c957737bf422127283c08e['h027cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013e7] =  Ifd35529b44c957737bf422127283c08e['h027ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013e8] =  Ifd35529b44c957737bf422127283c08e['h027d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013e9] =  Ifd35529b44c957737bf422127283c08e['h027d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013ea] =  Ifd35529b44c957737bf422127283c08e['h027d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013eb] =  Ifd35529b44c957737bf422127283c08e['h027d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013ec] =  Ifd35529b44c957737bf422127283c08e['h027d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013ed] =  Ifd35529b44c957737bf422127283c08e['h027da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013ee] =  Ifd35529b44c957737bf422127283c08e['h027dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013ef] =  Ifd35529b44c957737bf422127283c08e['h027de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013f0] =  Ifd35529b44c957737bf422127283c08e['h027e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013f1] =  Ifd35529b44c957737bf422127283c08e['h027e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013f2] =  Ifd35529b44c957737bf422127283c08e['h027e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013f3] =  Ifd35529b44c957737bf422127283c08e['h027e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013f4] =  Ifd35529b44c957737bf422127283c08e['h027e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013f5] =  Ifd35529b44c957737bf422127283c08e['h027ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013f6] =  Ifd35529b44c957737bf422127283c08e['h027ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013f7] =  Ifd35529b44c957737bf422127283c08e['h027ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013f8] =  Ifd35529b44c957737bf422127283c08e['h027f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013f9] =  Ifd35529b44c957737bf422127283c08e['h027f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013fa] =  Ifd35529b44c957737bf422127283c08e['h027f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013fb] =  Ifd35529b44c957737bf422127283c08e['h027f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013fc] =  Ifd35529b44c957737bf422127283c08e['h027f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013fd] =  Ifd35529b44c957737bf422127283c08e['h027fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013fe] =  Ifd35529b44c957737bf422127283c08e['h027fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h013ff] =  Ifd35529b44c957737bf422127283c08e['h027fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01400] =  Ifd35529b44c957737bf422127283c08e['h02800] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01401] =  Ifd35529b44c957737bf422127283c08e['h02802] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01402] =  Ifd35529b44c957737bf422127283c08e['h02804] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01403] =  Ifd35529b44c957737bf422127283c08e['h02806] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01404] =  Ifd35529b44c957737bf422127283c08e['h02808] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01405] =  Ifd35529b44c957737bf422127283c08e['h0280a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01406] =  Ifd35529b44c957737bf422127283c08e['h0280c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01407] =  Ifd35529b44c957737bf422127283c08e['h0280e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01408] =  Ifd35529b44c957737bf422127283c08e['h02810] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01409] =  Ifd35529b44c957737bf422127283c08e['h02812] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0140a] =  Ifd35529b44c957737bf422127283c08e['h02814] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0140b] =  Ifd35529b44c957737bf422127283c08e['h02816] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0140c] =  Ifd35529b44c957737bf422127283c08e['h02818] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0140d] =  Ifd35529b44c957737bf422127283c08e['h0281a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0140e] =  Ifd35529b44c957737bf422127283c08e['h0281c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0140f] =  Ifd35529b44c957737bf422127283c08e['h0281e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01410] =  Ifd35529b44c957737bf422127283c08e['h02820] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01411] =  Ifd35529b44c957737bf422127283c08e['h02822] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01412] =  Ifd35529b44c957737bf422127283c08e['h02824] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01413] =  Ifd35529b44c957737bf422127283c08e['h02826] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01414] =  Ifd35529b44c957737bf422127283c08e['h02828] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01415] =  Ifd35529b44c957737bf422127283c08e['h0282a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01416] =  Ifd35529b44c957737bf422127283c08e['h0282c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01417] =  Ifd35529b44c957737bf422127283c08e['h0282e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01418] =  Ifd35529b44c957737bf422127283c08e['h02830] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01419] =  Ifd35529b44c957737bf422127283c08e['h02832] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0141a] =  Ifd35529b44c957737bf422127283c08e['h02834] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0141b] =  Ifd35529b44c957737bf422127283c08e['h02836] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0141c] =  Ifd35529b44c957737bf422127283c08e['h02838] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0141d] =  Ifd35529b44c957737bf422127283c08e['h0283a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0141e] =  Ifd35529b44c957737bf422127283c08e['h0283c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0141f] =  Ifd35529b44c957737bf422127283c08e['h0283e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01420] =  Ifd35529b44c957737bf422127283c08e['h02840] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01421] =  Ifd35529b44c957737bf422127283c08e['h02842] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01422] =  Ifd35529b44c957737bf422127283c08e['h02844] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01423] =  Ifd35529b44c957737bf422127283c08e['h02846] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01424] =  Ifd35529b44c957737bf422127283c08e['h02848] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01425] =  Ifd35529b44c957737bf422127283c08e['h0284a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01426] =  Ifd35529b44c957737bf422127283c08e['h0284c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01427] =  Ifd35529b44c957737bf422127283c08e['h0284e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01428] =  Ifd35529b44c957737bf422127283c08e['h02850] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01429] =  Ifd35529b44c957737bf422127283c08e['h02852] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0142a] =  Ifd35529b44c957737bf422127283c08e['h02854] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0142b] =  Ifd35529b44c957737bf422127283c08e['h02856] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0142c] =  Ifd35529b44c957737bf422127283c08e['h02858] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0142d] =  Ifd35529b44c957737bf422127283c08e['h0285a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0142e] =  Ifd35529b44c957737bf422127283c08e['h0285c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0142f] =  Ifd35529b44c957737bf422127283c08e['h0285e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01430] =  Ifd35529b44c957737bf422127283c08e['h02860] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01431] =  Ifd35529b44c957737bf422127283c08e['h02862] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01432] =  Ifd35529b44c957737bf422127283c08e['h02864] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01433] =  Ifd35529b44c957737bf422127283c08e['h02866] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01434] =  Ifd35529b44c957737bf422127283c08e['h02868] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01435] =  Ifd35529b44c957737bf422127283c08e['h0286a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01436] =  Ifd35529b44c957737bf422127283c08e['h0286c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01437] =  Ifd35529b44c957737bf422127283c08e['h0286e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01438] =  Ifd35529b44c957737bf422127283c08e['h02870] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01439] =  Ifd35529b44c957737bf422127283c08e['h02872] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0143a] =  Ifd35529b44c957737bf422127283c08e['h02874] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0143b] =  Ifd35529b44c957737bf422127283c08e['h02876] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0143c] =  Ifd35529b44c957737bf422127283c08e['h02878] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0143d] =  Ifd35529b44c957737bf422127283c08e['h0287a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0143e] =  Ifd35529b44c957737bf422127283c08e['h0287c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0143f] =  Ifd35529b44c957737bf422127283c08e['h0287e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01440] =  Ifd35529b44c957737bf422127283c08e['h02880] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01441] =  Ifd35529b44c957737bf422127283c08e['h02882] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01442] =  Ifd35529b44c957737bf422127283c08e['h02884] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01443] =  Ifd35529b44c957737bf422127283c08e['h02886] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01444] =  Ifd35529b44c957737bf422127283c08e['h02888] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01445] =  Ifd35529b44c957737bf422127283c08e['h0288a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01446] =  Ifd35529b44c957737bf422127283c08e['h0288c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01447] =  Ifd35529b44c957737bf422127283c08e['h0288e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01448] =  Ifd35529b44c957737bf422127283c08e['h02890] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01449] =  Ifd35529b44c957737bf422127283c08e['h02892] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0144a] =  Ifd35529b44c957737bf422127283c08e['h02894] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0144b] =  Ifd35529b44c957737bf422127283c08e['h02896] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0144c] =  Ifd35529b44c957737bf422127283c08e['h02898] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0144d] =  Ifd35529b44c957737bf422127283c08e['h0289a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0144e] =  Ifd35529b44c957737bf422127283c08e['h0289c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0144f] =  Ifd35529b44c957737bf422127283c08e['h0289e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01450] =  Ifd35529b44c957737bf422127283c08e['h028a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01451] =  Ifd35529b44c957737bf422127283c08e['h028a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01452] =  Ifd35529b44c957737bf422127283c08e['h028a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01453] =  Ifd35529b44c957737bf422127283c08e['h028a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01454] =  Ifd35529b44c957737bf422127283c08e['h028a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01455] =  Ifd35529b44c957737bf422127283c08e['h028aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01456] =  Ifd35529b44c957737bf422127283c08e['h028ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01457] =  Ifd35529b44c957737bf422127283c08e['h028ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01458] =  Ifd35529b44c957737bf422127283c08e['h028b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01459] =  Ifd35529b44c957737bf422127283c08e['h028b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0145a] =  Ifd35529b44c957737bf422127283c08e['h028b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0145b] =  Ifd35529b44c957737bf422127283c08e['h028b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0145c] =  Ifd35529b44c957737bf422127283c08e['h028b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0145d] =  Ifd35529b44c957737bf422127283c08e['h028ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0145e] =  Ifd35529b44c957737bf422127283c08e['h028bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0145f] =  Ifd35529b44c957737bf422127283c08e['h028be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01460] =  Ifd35529b44c957737bf422127283c08e['h028c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01461] =  Ifd35529b44c957737bf422127283c08e['h028c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01462] =  Ifd35529b44c957737bf422127283c08e['h028c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01463] =  Ifd35529b44c957737bf422127283c08e['h028c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01464] =  Ifd35529b44c957737bf422127283c08e['h028c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01465] =  Ifd35529b44c957737bf422127283c08e['h028ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01466] =  Ifd35529b44c957737bf422127283c08e['h028cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01467] =  Ifd35529b44c957737bf422127283c08e['h028ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01468] =  Ifd35529b44c957737bf422127283c08e['h028d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01469] =  Ifd35529b44c957737bf422127283c08e['h028d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0146a] =  Ifd35529b44c957737bf422127283c08e['h028d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0146b] =  Ifd35529b44c957737bf422127283c08e['h028d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0146c] =  Ifd35529b44c957737bf422127283c08e['h028d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0146d] =  Ifd35529b44c957737bf422127283c08e['h028da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0146e] =  Ifd35529b44c957737bf422127283c08e['h028dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0146f] =  Ifd35529b44c957737bf422127283c08e['h028de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01470] =  Ifd35529b44c957737bf422127283c08e['h028e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01471] =  Ifd35529b44c957737bf422127283c08e['h028e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01472] =  Ifd35529b44c957737bf422127283c08e['h028e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01473] =  Ifd35529b44c957737bf422127283c08e['h028e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01474] =  Ifd35529b44c957737bf422127283c08e['h028e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01475] =  Ifd35529b44c957737bf422127283c08e['h028ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01476] =  Ifd35529b44c957737bf422127283c08e['h028ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01477] =  Ifd35529b44c957737bf422127283c08e['h028ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01478] =  Ifd35529b44c957737bf422127283c08e['h028f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01479] =  Ifd35529b44c957737bf422127283c08e['h028f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0147a] =  Ifd35529b44c957737bf422127283c08e['h028f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0147b] =  Ifd35529b44c957737bf422127283c08e['h028f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0147c] =  Ifd35529b44c957737bf422127283c08e['h028f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0147d] =  Ifd35529b44c957737bf422127283c08e['h028fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0147e] =  Ifd35529b44c957737bf422127283c08e['h028fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0147f] =  Ifd35529b44c957737bf422127283c08e['h028fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01480] =  Ifd35529b44c957737bf422127283c08e['h02900] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01481] =  Ifd35529b44c957737bf422127283c08e['h02902] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01482] =  Ifd35529b44c957737bf422127283c08e['h02904] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01483] =  Ifd35529b44c957737bf422127283c08e['h02906] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01484] =  Ifd35529b44c957737bf422127283c08e['h02908] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01485] =  Ifd35529b44c957737bf422127283c08e['h0290a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01486] =  Ifd35529b44c957737bf422127283c08e['h0290c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01487] =  Ifd35529b44c957737bf422127283c08e['h0290e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01488] =  Ifd35529b44c957737bf422127283c08e['h02910] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01489] =  Ifd35529b44c957737bf422127283c08e['h02912] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0148a] =  Ifd35529b44c957737bf422127283c08e['h02914] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0148b] =  Ifd35529b44c957737bf422127283c08e['h02916] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0148c] =  Ifd35529b44c957737bf422127283c08e['h02918] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0148d] =  Ifd35529b44c957737bf422127283c08e['h0291a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0148e] =  Ifd35529b44c957737bf422127283c08e['h0291c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0148f] =  Ifd35529b44c957737bf422127283c08e['h0291e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01490] =  Ifd35529b44c957737bf422127283c08e['h02920] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01491] =  Ifd35529b44c957737bf422127283c08e['h02922] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01492] =  Ifd35529b44c957737bf422127283c08e['h02924] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01493] =  Ifd35529b44c957737bf422127283c08e['h02926] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01494] =  Ifd35529b44c957737bf422127283c08e['h02928] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01495] =  Ifd35529b44c957737bf422127283c08e['h0292a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01496] =  Ifd35529b44c957737bf422127283c08e['h0292c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01497] =  Ifd35529b44c957737bf422127283c08e['h0292e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01498] =  Ifd35529b44c957737bf422127283c08e['h02930] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01499] =  Ifd35529b44c957737bf422127283c08e['h02932] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0149a] =  Ifd35529b44c957737bf422127283c08e['h02934] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0149b] =  Ifd35529b44c957737bf422127283c08e['h02936] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0149c] =  Ifd35529b44c957737bf422127283c08e['h02938] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0149d] =  Ifd35529b44c957737bf422127283c08e['h0293a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0149e] =  Ifd35529b44c957737bf422127283c08e['h0293c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0149f] =  Ifd35529b44c957737bf422127283c08e['h0293e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014a0] =  Ifd35529b44c957737bf422127283c08e['h02940] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014a1] =  Ifd35529b44c957737bf422127283c08e['h02942] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014a2] =  Ifd35529b44c957737bf422127283c08e['h02944] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014a3] =  Ifd35529b44c957737bf422127283c08e['h02946] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014a4] =  Ifd35529b44c957737bf422127283c08e['h02948] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014a5] =  Ifd35529b44c957737bf422127283c08e['h0294a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014a6] =  Ifd35529b44c957737bf422127283c08e['h0294c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014a7] =  Ifd35529b44c957737bf422127283c08e['h0294e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014a8] =  Ifd35529b44c957737bf422127283c08e['h02950] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014a9] =  Ifd35529b44c957737bf422127283c08e['h02952] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014aa] =  Ifd35529b44c957737bf422127283c08e['h02954] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014ab] =  Ifd35529b44c957737bf422127283c08e['h02956] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014ac] =  Ifd35529b44c957737bf422127283c08e['h02958] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014ad] =  Ifd35529b44c957737bf422127283c08e['h0295a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014ae] =  Ifd35529b44c957737bf422127283c08e['h0295c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014af] =  Ifd35529b44c957737bf422127283c08e['h0295e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014b0] =  Ifd35529b44c957737bf422127283c08e['h02960] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014b1] =  Ifd35529b44c957737bf422127283c08e['h02962] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014b2] =  Ifd35529b44c957737bf422127283c08e['h02964] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014b3] =  Ifd35529b44c957737bf422127283c08e['h02966] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014b4] =  Ifd35529b44c957737bf422127283c08e['h02968] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014b5] =  Ifd35529b44c957737bf422127283c08e['h0296a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014b6] =  Ifd35529b44c957737bf422127283c08e['h0296c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014b7] =  Ifd35529b44c957737bf422127283c08e['h0296e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014b8] =  Ifd35529b44c957737bf422127283c08e['h02970] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014b9] =  Ifd35529b44c957737bf422127283c08e['h02972] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014ba] =  Ifd35529b44c957737bf422127283c08e['h02974] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014bb] =  Ifd35529b44c957737bf422127283c08e['h02976] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014bc] =  Ifd35529b44c957737bf422127283c08e['h02978] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014bd] =  Ifd35529b44c957737bf422127283c08e['h0297a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014be] =  Ifd35529b44c957737bf422127283c08e['h0297c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014bf] =  Ifd35529b44c957737bf422127283c08e['h0297e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014c0] =  Ifd35529b44c957737bf422127283c08e['h02980] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014c1] =  Ifd35529b44c957737bf422127283c08e['h02982] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014c2] =  Ifd35529b44c957737bf422127283c08e['h02984] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014c3] =  Ifd35529b44c957737bf422127283c08e['h02986] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014c4] =  Ifd35529b44c957737bf422127283c08e['h02988] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014c5] =  Ifd35529b44c957737bf422127283c08e['h0298a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014c6] =  Ifd35529b44c957737bf422127283c08e['h0298c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014c7] =  Ifd35529b44c957737bf422127283c08e['h0298e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014c8] =  Ifd35529b44c957737bf422127283c08e['h02990] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014c9] =  Ifd35529b44c957737bf422127283c08e['h02992] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014ca] =  Ifd35529b44c957737bf422127283c08e['h02994] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014cb] =  Ifd35529b44c957737bf422127283c08e['h02996] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014cc] =  Ifd35529b44c957737bf422127283c08e['h02998] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014cd] =  Ifd35529b44c957737bf422127283c08e['h0299a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014ce] =  Ifd35529b44c957737bf422127283c08e['h0299c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014cf] =  Ifd35529b44c957737bf422127283c08e['h0299e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014d0] =  Ifd35529b44c957737bf422127283c08e['h029a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014d1] =  Ifd35529b44c957737bf422127283c08e['h029a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014d2] =  Ifd35529b44c957737bf422127283c08e['h029a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014d3] =  Ifd35529b44c957737bf422127283c08e['h029a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014d4] =  Ifd35529b44c957737bf422127283c08e['h029a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014d5] =  Ifd35529b44c957737bf422127283c08e['h029aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014d6] =  Ifd35529b44c957737bf422127283c08e['h029ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014d7] =  Ifd35529b44c957737bf422127283c08e['h029ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014d8] =  Ifd35529b44c957737bf422127283c08e['h029b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014d9] =  Ifd35529b44c957737bf422127283c08e['h029b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014da] =  Ifd35529b44c957737bf422127283c08e['h029b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014db] =  Ifd35529b44c957737bf422127283c08e['h029b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014dc] =  Ifd35529b44c957737bf422127283c08e['h029b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014dd] =  Ifd35529b44c957737bf422127283c08e['h029ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014de] =  Ifd35529b44c957737bf422127283c08e['h029bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014df] =  Ifd35529b44c957737bf422127283c08e['h029be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014e0] =  Ifd35529b44c957737bf422127283c08e['h029c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014e1] =  Ifd35529b44c957737bf422127283c08e['h029c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014e2] =  Ifd35529b44c957737bf422127283c08e['h029c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014e3] =  Ifd35529b44c957737bf422127283c08e['h029c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014e4] =  Ifd35529b44c957737bf422127283c08e['h029c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014e5] =  Ifd35529b44c957737bf422127283c08e['h029ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014e6] =  Ifd35529b44c957737bf422127283c08e['h029cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014e7] =  Ifd35529b44c957737bf422127283c08e['h029ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014e8] =  Ifd35529b44c957737bf422127283c08e['h029d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014e9] =  Ifd35529b44c957737bf422127283c08e['h029d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014ea] =  Ifd35529b44c957737bf422127283c08e['h029d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014eb] =  Ifd35529b44c957737bf422127283c08e['h029d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014ec] =  Ifd35529b44c957737bf422127283c08e['h029d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014ed] =  Ifd35529b44c957737bf422127283c08e['h029da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014ee] =  Ifd35529b44c957737bf422127283c08e['h029dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014ef] =  Ifd35529b44c957737bf422127283c08e['h029de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014f0] =  Ifd35529b44c957737bf422127283c08e['h029e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014f1] =  Ifd35529b44c957737bf422127283c08e['h029e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014f2] =  Ifd35529b44c957737bf422127283c08e['h029e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014f3] =  Ifd35529b44c957737bf422127283c08e['h029e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014f4] =  Ifd35529b44c957737bf422127283c08e['h029e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014f5] =  Ifd35529b44c957737bf422127283c08e['h029ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014f6] =  Ifd35529b44c957737bf422127283c08e['h029ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014f7] =  Ifd35529b44c957737bf422127283c08e['h029ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014f8] =  Ifd35529b44c957737bf422127283c08e['h029f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014f9] =  Ifd35529b44c957737bf422127283c08e['h029f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014fa] =  Ifd35529b44c957737bf422127283c08e['h029f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014fb] =  Ifd35529b44c957737bf422127283c08e['h029f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014fc] =  Ifd35529b44c957737bf422127283c08e['h029f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014fd] =  Ifd35529b44c957737bf422127283c08e['h029fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014fe] =  Ifd35529b44c957737bf422127283c08e['h029fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h014ff] =  Ifd35529b44c957737bf422127283c08e['h029fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01500] =  Ifd35529b44c957737bf422127283c08e['h02a00] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01501] =  Ifd35529b44c957737bf422127283c08e['h02a02] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01502] =  Ifd35529b44c957737bf422127283c08e['h02a04] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01503] =  Ifd35529b44c957737bf422127283c08e['h02a06] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01504] =  Ifd35529b44c957737bf422127283c08e['h02a08] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01505] =  Ifd35529b44c957737bf422127283c08e['h02a0a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01506] =  Ifd35529b44c957737bf422127283c08e['h02a0c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01507] =  Ifd35529b44c957737bf422127283c08e['h02a0e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01508] =  Ifd35529b44c957737bf422127283c08e['h02a10] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01509] =  Ifd35529b44c957737bf422127283c08e['h02a12] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0150a] =  Ifd35529b44c957737bf422127283c08e['h02a14] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0150b] =  Ifd35529b44c957737bf422127283c08e['h02a16] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0150c] =  Ifd35529b44c957737bf422127283c08e['h02a18] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0150d] =  Ifd35529b44c957737bf422127283c08e['h02a1a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0150e] =  Ifd35529b44c957737bf422127283c08e['h02a1c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0150f] =  Ifd35529b44c957737bf422127283c08e['h02a1e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01510] =  Ifd35529b44c957737bf422127283c08e['h02a20] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01511] =  Ifd35529b44c957737bf422127283c08e['h02a22] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01512] =  Ifd35529b44c957737bf422127283c08e['h02a24] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01513] =  Ifd35529b44c957737bf422127283c08e['h02a26] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01514] =  Ifd35529b44c957737bf422127283c08e['h02a28] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01515] =  Ifd35529b44c957737bf422127283c08e['h02a2a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01516] =  Ifd35529b44c957737bf422127283c08e['h02a2c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01517] =  Ifd35529b44c957737bf422127283c08e['h02a2e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01518] =  Ifd35529b44c957737bf422127283c08e['h02a30] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01519] =  Ifd35529b44c957737bf422127283c08e['h02a32] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0151a] =  Ifd35529b44c957737bf422127283c08e['h02a34] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0151b] =  Ifd35529b44c957737bf422127283c08e['h02a36] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0151c] =  Ifd35529b44c957737bf422127283c08e['h02a38] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0151d] =  Ifd35529b44c957737bf422127283c08e['h02a3a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0151e] =  Ifd35529b44c957737bf422127283c08e['h02a3c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0151f] =  Ifd35529b44c957737bf422127283c08e['h02a3e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01520] =  Ifd35529b44c957737bf422127283c08e['h02a40] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01521] =  Ifd35529b44c957737bf422127283c08e['h02a42] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01522] =  Ifd35529b44c957737bf422127283c08e['h02a44] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01523] =  Ifd35529b44c957737bf422127283c08e['h02a46] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01524] =  Ifd35529b44c957737bf422127283c08e['h02a48] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01525] =  Ifd35529b44c957737bf422127283c08e['h02a4a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01526] =  Ifd35529b44c957737bf422127283c08e['h02a4c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01527] =  Ifd35529b44c957737bf422127283c08e['h02a4e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01528] =  Ifd35529b44c957737bf422127283c08e['h02a50] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01529] =  Ifd35529b44c957737bf422127283c08e['h02a52] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0152a] =  Ifd35529b44c957737bf422127283c08e['h02a54] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0152b] =  Ifd35529b44c957737bf422127283c08e['h02a56] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0152c] =  Ifd35529b44c957737bf422127283c08e['h02a58] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0152d] =  Ifd35529b44c957737bf422127283c08e['h02a5a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0152e] =  Ifd35529b44c957737bf422127283c08e['h02a5c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0152f] =  Ifd35529b44c957737bf422127283c08e['h02a5e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01530] =  Ifd35529b44c957737bf422127283c08e['h02a60] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01531] =  Ifd35529b44c957737bf422127283c08e['h02a62] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01532] =  Ifd35529b44c957737bf422127283c08e['h02a64] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01533] =  Ifd35529b44c957737bf422127283c08e['h02a66] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01534] =  Ifd35529b44c957737bf422127283c08e['h02a68] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01535] =  Ifd35529b44c957737bf422127283c08e['h02a6a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01536] =  Ifd35529b44c957737bf422127283c08e['h02a6c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01537] =  Ifd35529b44c957737bf422127283c08e['h02a6e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01538] =  Ifd35529b44c957737bf422127283c08e['h02a70] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01539] =  Ifd35529b44c957737bf422127283c08e['h02a72] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0153a] =  Ifd35529b44c957737bf422127283c08e['h02a74] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0153b] =  Ifd35529b44c957737bf422127283c08e['h02a76] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0153c] =  Ifd35529b44c957737bf422127283c08e['h02a78] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0153d] =  Ifd35529b44c957737bf422127283c08e['h02a7a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0153e] =  Ifd35529b44c957737bf422127283c08e['h02a7c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0153f] =  Ifd35529b44c957737bf422127283c08e['h02a7e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01540] =  Ifd35529b44c957737bf422127283c08e['h02a80] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01541] =  Ifd35529b44c957737bf422127283c08e['h02a82] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01542] =  Ifd35529b44c957737bf422127283c08e['h02a84] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01543] =  Ifd35529b44c957737bf422127283c08e['h02a86] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01544] =  Ifd35529b44c957737bf422127283c08e['h02a88] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01545] =  Ifd35529b44c957737bf422127283c08e['h02a8a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01546] =  Ifd35529b44c957737bf422127283c08e['h02a8c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01547] =  Ifd35529b44c957737bf422127283c08e['h02a8e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01548] =  Ifd35529b44c957737bf422127283c08e['h02a90] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01549] =  Ifd35529b44c957737bf422127283c08e['h02a92] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0154a] =  Ifd35529b44c957737bf422127283c08e['h02a94] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0154b] =  Ifd35529b44c957737bf422127283c08e['h02a96] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0154c] =  Ifd35529b44c957737bf422127283c08e['h02a98] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0154d] =  Ifd35529b44c957737bf422127283c08e['h02a9a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0154e] =  Ifd35529b44c957737bf422127283c08e['h02a9c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0154f] =  Ifd35529b44c957737bf422127283c08e['h02a9e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01550] =  Ifd35529b44c957737bf422127283c08e['h02aa0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01551] =  Ifd35529b44c957737bf422127283c08e['h02aa2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01552] =  Ifd35529b44c957737bf422127283c08e['h02aa4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01553] =  Ifd35529b44c957737bf422127283c08e['h02aa6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01554] =  Ifd35529b44c957737bf422127283c08e['h02aa8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01555] =  Ifd35529b44c957737bf422127283c08e['h02aaa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01556] =  Ifd35529b44c957737bf422127283c08e['h02aac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01557] =  Ifd35529b44c957737bf422127283c08e['h02aae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01558] =  Ifd35529b44c957737bf422127283c08e['h02ab0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01559] =  Ifd35529b44c957737bf422127283c08e['h02ab2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0155a] =  Ifd35529b44c957737bf422127283c08e['h02ab4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0155b] =  Ifd35529b44c957737bf422127283c08e['h02ab6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0155c] =  Ifd35529b44c957737bf422127283c08e['h02ab8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0155d] =  Ifd35529b44c957737bf422127283c08e['h02aba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0155e] =  Ifd35529b44c957737bf422127283c08e['h02abc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0155f] =  Ifd35529b44c957737bf422127283c08e['h02abe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01560] =  Ifd35529b44c957737bf422127283c08e['h02ac0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01561] =  Ifd35529b44c957737bf422127283c08e['h02ac2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01562] =  Ifd35529b44c957737bf422127283c08e['h02ac4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01563] =  Ifd35529b44c957737bf422127283c08e['h02ac6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01564] =  Ifd35529b44c957737bf422127283c08e['h02ac8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01565] =  Ifd35529b44c957737bf422127283c08e['h02aca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01566] =  Ifd35529b44c957737bf422127283c08e['h02acc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01567] =  Ifd35529b44c957737bf422127283c08e['h02ace] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01568] =  Ifd35529b44c957737bf422127283c08e['h02ad0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01569] =  Ifd35529b44c957737bf422127283c08e['h02ad2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0156a] =  Ifd35529b44c957737bf422127283c08e['h02ad4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0156b] =  Ifd35529b44c957737bf422127283c08e['h02ad6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0156c] =  Ifd35529b44c957737bf422127283c08e['h02ad8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0156d] =  Ifd35529b44c957737bf422127283c08e['h02ada] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0156e] =  Ifd35529b44c957737bf422127283c08e['h02adc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0156f] =  Ifd35529b44c957737bf422127283c08e['h02ade] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01570] =  Ifd35529b44c957737bf422127283c08e['h02ae0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01571] =  Ifd35529b44c957737bf422127283c08e['h02ae2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01572] =  Ifd35529b44c957737bf422127283c08e['h02ae4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01573] =  Ifd35529b44c957737bf422127283c08e['h02ae6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01574] =  Ifd35529b44c957737bf422127283c08e['h02ae8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01575] =  Ifd35529b44c957737bf422127283c08e['h02aea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01576] =  Ifd35529b44c957737bf422127283c08e['h02aec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01577] =  Ifd35529b44c957737bf422127283c08e['h02aee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01578] =  Ifd35529b44c957737bf422127283c08e['h02af0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01579] =  Ifd35529b44c957737bf422127283c08e['h02af2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0157a] =  Ifd35529b44c957737bf422127283c08e['h02af4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0157b] =  Ifd35529b44c957737bf422127283c08e['h02af6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0157c] =  Ifd35529b44c957737bf422127283c08e['h02af8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0157d] =  Ifd35529b44c957737bf422127283c08e['h02afa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0157e] =  Ifd35529b44c957737bf422127283c08e['h02afc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0157f] =  Ifd35529b44c957737bf422127283c08e['h02afe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01580] =  Ifd35529b44c957737bf422127283c08e['h02b00] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01581] =  Ifd35529b44c957737bf422127283c08e['h02b02] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01582] =  Ifd35529b44c957737bf422127283c08e['h02b04] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01583] =  Ifd35529b44c957737bf422127283c08e['h02b06] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01584] =  Ifd35529b44c957737bf422127283c08e['h02b08] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01585] =  Ifd35529b44c957737bf422127283c08e['h02b0a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01586] =  Ifd35529b44c957737bf422127283c08e['h02b0c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01587] =  Ifd35529b44c957737bf422127283c08e['h02b0e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01588] =  Ifd35529b44c957737bf422127283c08e['h02b10] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01589] =  Ifd35529b44c957737bf422127283c08e['h02b12] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0158a] =  Ifd35529b44c957737bf422127283c08e['h02b14] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0158b] =  Ifd35529b44c957737bf422127283c08e['h02b16] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0158c] =  Ifd35529b44c957737bf422127283c08e['h02b18] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0158d] =  Ifd35529b44c957737bf422127283c08e['h02b1a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0158e] =  Ifd35529b44c957737bf422127283c08e['h02b1c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0158f] =  Ifd35529b44c957737bf422127283c08e['h02b1e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01590] =  Ifd35529b44c957737bf422127283c08e['h02b20] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01591] =  Ifd35529b44c957737bf422127283c08e['h02b22] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01592] =  Ifd35529b44c957737bf422127283c08e['h02b24] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01593] =  Ifd35529b44c957737bf422127283c08e['h02b26] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01594] =  Ifd35529b44c957737bf422127283c08e['h02b28] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01595] =  Ifd35529b44c957737bf422127283c08e['h02b2a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01596] =  Ifd35529b44c957737bf422127283c08e['h02b2c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01597] =  Ifd35529b44c957737bf422127283c08e['h02b2e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01598] =  Ifd35529b44c957737bf422127283c08e['h02b30] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01599] =  Ifd35529b44c957737bf422127283c08e['h02b32] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0159a] =  Ifd35529b44c957737bf422127283c08e['h02b34] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0159b] =  Ifd35529b44c957737bf422127283c08e['h02b36] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0159c] =  Ifd35529b44c957737bf422127283c08e['h02b38] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0159d] =  Ifd35529b44c957737bf422127283c08e['h02b3a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0159e] =  Ifd35529b44c957737bf422127283c08e['h02b3c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0159f] =  Ifd35529b44c957737bf422127283c08e['h02b3e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015a0] =  Ifd35529b44c957737bf422127283c08e['h02b40] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015a1] =  Ifd35529b44c957737bf422127283c08e['h02b42] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015a2] =  Ifd35529b44c957737bf422127283c08e['h02b44] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015a3] =  Ifd35529b44c957737bf422127283c08e['h02b46] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015a4] =  Ifd35529b44c957737bf422127283c08e['h02b48] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015a5] =  Ifd35529b44c957737bf422127283c08e['h02b4a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015a6] =  Ifd35529b44c957737bf422127283c08e['h02b4c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015a7] =  Ifd35529b44c957737bf422127283c08e['h02b4e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015a8] =  Ifd35529b44c957737bf422127283c08e['h02b50] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015a9] =  Ifd35529b44c957737bf422127283c08e['h02b52] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015aa] =  Ifd35529b44c957737bf422127283c08e['h02b54] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015ab] =  Ifd35529b44c957737bf422127283c08e['h02b56] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015ac] =  Ifd35529b44c957737bf422127283c08e['h02b58] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015ad] =  Ifd35529b44c957737bf422127283c08e['h02b5a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015ae] =  Ifd35529b44c957737bf422127283c08e['h02b5c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015af] =  Ifd35529b44c957737bf422127283c08e['h02b5e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015b0] =  Ifd35529b44c957737bf422127283c08e['h02b60] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015b1] =  Ifd35529b44c957737bf422127283c08e['h02b62] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015b2] =  Ifd35529b44c957737bf422127283c08e['h02b64] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015b3] =  Ifd35529b44c957737bf422127283c08e['h02b66] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015b4] =  Ifd35529b44c957737bf422127283c08e['h02b68] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015b5] =  Ifd35529b44c957737bf422127283c08e['h02b6a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015b6] =  Ifd35529b44c957737bf422127283c08e['h02b6c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015b7] =  Ifd35529b44c957737bf422127283c08e['h02b6e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015b8] =  Ifd35529b44c957737bf422127283c08e['h02b70] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015b9] =  Ifd35529b44c957737bf422127283c08e['h02b72] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015ba] =  Ifd35529b44c957737bf422127283c08e['h02b74] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015bb] =  Ifd35529b44c957737bf422127283c08e['h02b76] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015bc] =  Ifd35529b44c957737bf422127283c08e['h02b78] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015bd] =  Ifd35529b44c957737bf422127283c08e['h02b7a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015be] =  Ifd35529b44c957737bf422127283c08e['h02b7c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015bf] =  Ifd35529b44c957737bf422127283c08e['h02b7e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015c0] =  Ifd35529b44c957737bf422127283c08e['h02b80] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015c1] =  Ifd35529b44c957737bf422127283c08e['h02b82] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015c2] =  Ifd35529b44c957737bf422127283c08e['h02b84] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015c3] =  Ifd35529b44c957737bf422127283c08e['h02b86] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015c4] =  Ifd35529b44c957737bf422127283c08e['h02b88] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015c5] =  Ifd35529b44c957737bf422127283c08e['h02b8a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015c6] =  Ifd35529b44c957737bf422127283c08e['h02b8c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015c7] =  Ifd35529b44c957737bf422127283c08e['h02b8e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015c8] =  Ifd35529b44c957737bf422127283c08e['h02b90] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015c9] =  Ifd35529b44c957737bf422127283c08e['h02b92] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015ca] =  Ifd35529b44c957737bf422127283c08e['h02b94] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015cb] =  Ifd35529b44c957737bf422127283c08e['h02b96] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015cc] =  Ifd35529b44c957737bf422127283c08e['h02b98] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015cd] =  Ifd35529b44c957737bf422127283c08e['h02b9a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015ce] =  Ifd35529b44c957737bf422127283c08e['h02b9c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015cf] =  Ifd35529b44c957737bf422127283c08e['h02b9e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015d0] =  Ifd35529b44c957737bf422127283c08e['h02ba0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015d1] =  Ifd35529b44c957737bf422127283c08e['h02ba2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015d2] =  Ifd35529b44c957737bf422127283c08e['h02ba4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015d3] =  Ifd35529b44c957737bf422127283c08e['h02ba6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015d4] =  Ifd35529b44c957737bf422127283c08e['h02ba8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015d5] =  Ifd35529b44c957737bf422127283c08e['h02baa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015d6] =  Ifd35529b44c957737bf422127283c08e['h02bac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015d7] =  Ifd35529b44c957737bf422127283c08e['h02bae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015d8] =  Ifd35529b44c957737bf422127283c08e['h02bb0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015d9] =  Ifd35529b44c957737bf422127283c08e['h02bb2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015da] =  Ifd35529b44c957737bf422127283c08e['h02bb4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015db] =  Ifd35529b44c957737bf422127283c08e['h02bb6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015dc] =  Ifd35529b44c957737bf422127283c08e['h02bb8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015dd] =  Ifd35529b44c957737bf422127283c08e['h02bba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015de] =  Ifd35529b44c957737bf422127283c08e['h02bbc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015df] =  Ifd35529b44c957737bf422127283c08e['h02bbe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015e0] =  Ifd35529b44c957737bf422127283c08e['h02bc0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015e1] =  Ifd35529b44c957737bf422127283c08e['h02bc2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015e2] =  Ifd35529b44c957737bf422127283c08e['h02bc4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015e3] =  Ifd35529b44c957737bf422127283c08e['h02bc6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015e4] =  Ifd35529b44c957737bf422127283c08e['h02bc8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015e5] =  Ifd35529b44c957737bf422127283c08e['h02bca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015e6] =  Ifd35529b44c957737bf422127283c08e['h02bcc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015e7] =  Ifd35529b44c957737bf422127283c08e['h02bce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015e8] =  Ifd35529b44c957737bf422127283c08e['h02bd0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015e9] =  Ifd35529b44c957737bf422127283c08e['h02bd2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015ea] =  Ifd35529b44c957737bf422127283c08e['h02bd4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015eb] =  Ifd35529b44c957737bf422127283c08e['h02bd6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015ec] =  Ifd35529b44c957737bf422127283c08e['h02bd8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015ed] =  Ifd35529b44c957737bf422127283c08e['h02bda] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015ee] =  Ifd35529b44c957737bf422127283c08e['h02bdc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015ef] =  Ifd35529b44c957737bf422127283c08e['h02bde] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015f0] =  Ifd35529b44c957737bf422127283c08e['h02be0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015f1] =  Ifd35529b44c957737bf422127283c08e['h02be2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015f2] =  Ifd35529b44c957737bf422127283c08e['h02be4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015f3] =  Ifd35529b44c957737bf422127283c08e['h02be6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015f4] =  Ifd35529b44c957737bf422127283c08e['h02be8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015f5] =  Ifd35529b44c957737bf422127283c08e['h02bea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015f6] =  Ifd35529b44c957737bf422127283c08e['h02bec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015f7] =  Ifd35529b44c957737bf422127283c08e['h02bee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015f8] =  Ifd35529b44c957737bf422127283c08e['h02bf0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015f9] =  Ifd35529b44c957737bf422127283c08e['h02bf2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015fa] =  Ifd35529b44c957737bf422127283c08e['h02bf4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015fb] =  Ifd35529b44c957737bf422127283c08e['h02bf6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015fc] =  Ifd35529b44c957737bf422127283c08e['h02bf8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015fd] =  Ifd35529b44c957737bf422127283c08e['h02bfa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015fe] =  Ifd35529b44c957737bf422127283c08e['h02bfc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h015ff] =  Ifd35529b44c957737bf422127283c08e['h02bfe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01600] =  Ifd35529b44c957737bf422127283c08e['h02c00] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01601] =  Ifd35529b44c957737bf422127283c08e['h02c02] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01602] =  Ifd35529b44c957737bf422127283c08e['h02c04] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01603] =  Ifd35529b44c957737bf422127283c08e['h02c06] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01604] =  Ifd35529b44c957737bf422127283c08e['h02c08] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01605] =  Ifd35529b44c957737bf422127283c08e['h02c0a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01606] =  Ifd35529b44c957737bf422127283c08e['h02c0c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01607] =  Ifd35529b44c957737bf422127283c08e['h02c0e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01608] =  Ifd35529b44c957737bf422127283c08e['h02c10] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01609] =  Ifd35529b44c957737bf422127283c08e['h02c12] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0160a] =  Ifd35529b44c957737bf422127283c08e['h02c14] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0160b] =  Ifd35529b44c957737bf422127283c08e['h02c16] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0160c] =  Ifd35529b44c957737bf422127283c08e['h02c18] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0160d] =  Ifd35529b44c957737bf422127283c08e['h02c1a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0160e] =  Ifd35529b44c957737bf422127283c08e['h02c1c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0160f] =  Ifd35529b44c957737bf422127283c08e['h02c1e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01610] =  Ifd35529b44c957737bf422127283c08e['h02c20] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01611] =  Ifd35529b44c957737bf422127283c08e['h02c22] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01612] =  Ifd35529b44c957737bf422127283c08e['h02c24] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01613] =  Ifd35529b44c957737bf422127283c08e['h02c26] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01614] =  Ifd35529b44c957737bf422127283c08e['h02c28] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01615] =  Ifd35529b44c957737bf422127283c08e['h02c2a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01616] =  Ifd35529b44c957737bf422127283c08e['h02c2c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01617] =  Ifd35529b44c957737bf422127283c08e['h02c2e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01618] =  Ifd35529b44c957737bf422127283c08e['h02c30] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01619] =  Ifd35529b44c957737bf422127283c08e['h02c32] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0161a] =  Ifd35529b44c957737bf422127283c08e['h02c34] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0161b] =  Ifd35529b44c957737bf422127283c08e['h02c36] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0161c] =  Ifd35529b44c957737bf422127283c08e['h02c38] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0161d] =  Ifd35529b44c957737bf422127283c08e['h02c3a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0161e] =  Ifd35529b44c957737bf422127283c08e['h02c3c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0161f] =  Ifd35529b44c957737bf422127283c08e['h02c3e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01620] =  Ifd35529b44c957737bf422127283c08e['h02c40] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01621] =  Ifd35529b44c957737bf422127283c08e['h02c42] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01622] =  Ifd35529b44c957737bf422127283c08e['h02c44] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01623] =  Ifd35529b44c957737bf422127283c08e['h02c46] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01624] =  Ifd35529b44c957737bf422127283c08e['h02c48] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01625] =  Ifd35529b44c957737bf422127283c08e['h02c4a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01626] =  Ifd35529b44c957737bf422127283c08e['h02c4c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01627] =  Ifd35529b44c957737bf422127283c08e['h02c4e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01628] =  Ifd35529b44c957737bf422127283c08e['h02c50] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01629] =  Ifd35529b44c957737bf422127283c08e['h02c52] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0162a] =  Ifd35529b44c957737bf422127283c08e['h02c54] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0162b] =  Ifd35529b44c957737bf422127283c08e['h02c56] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0162c] =  Ifd35529b44c957737bf422127283c08e['h02c58] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0162d] =  Ifd35529b44c957737bf422127283c08e['h02c5a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0162e] =  Ifd35529b44c957737bf422127283c08e['h02c5c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0162f] =  Ifd35529b44c957737bf422127283c08e['h02c5e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01630] =  Ifd35529b44c957737bf422127283c08e['h02c60] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01631] =  Ifd35529b44c957737bf422127283c08e['h02c62] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01632] =  Ifd35529b44c957737bf422127283c08e['h02c64] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01633] =  Ifd35529b44c957737bf422127283c08e['h02c66] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01634] =  Ifd35529b44c957737bf422127283c08e['h02c68] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01635] =  Ifd35529b44c957737bf422127283c08e['h02c6a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01636] =  Ifd35529b44c957737bf422127283c08e['h02c6c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01637] =  Ifd35529b44c957737bf422127283c08e['h02c6e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01638] =  Ifd35529b44c957737bf422127283c08e['h02c70] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01639] =  Ifd35529b44c957737bf422127283c08e['h02c72] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0163a] =  Ifd35529b44c957737bf422127283c08e['h02c74] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0163b] =  Ifd35529b44c957737bf422127283c08e['h02c76] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0163c] =  Ifd35529b44c957737bf422127283c08e['h02c78] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0163d] =  Ifd35529b44c957737bf422127283c08e['h02c7a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0163e] =  Ifd35529b44c957737bf422127283c08e['h02c7c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0163f] =  Ifd35529b44c957737bf422127283c08e['h02c7e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01640] =  Ifd35529b44c957737bf422127283c08e['h02c80] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01641] =  Ifd35529b44c957737bf422127283c08e['h02c82] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01642] =  Ifd35529b44c957737bf422127283c08e['h02c84] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01643] =  Ifd35529b44c957737bf422127283c08e['h02c86] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01644] =  Ifd35529b44c957737bf422127283c08e['h02c88] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01645] =  Ifd35529b44c957737bf422127283c08e['h02c8a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01646] =  Ifd35529b44c957737bf422127283c08e['h02c8c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01647] =  Ifd35529b44c957737bf422127283c08e['h02c8e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01648] =  Ifd35529b44c957737bf422127283c08e['h02c90] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01649] =  Ifd35529b44c957737bf422127283c08e['h02c92] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0164a] =  Ifd35529b44c957737bf422127283c08e['h02c94] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0164b] =  Ifd35529b44c957737bf422127283c08e['h02c96] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0164c] =  Ifd35529b44c957737bf422127283c08e['h02c98] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0164d] =  Ifd35529b44c957737bf422127283c08e['h02c9a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0164e] =  Ifd35529b44c957737bf422127283c08e['h02c9c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0164f] =  Ifd35529b44c957737bf422127283c08e['h02c9e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01650] =  Ifd35529b44c957737bf422127283c08e['h02ca0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01651] =  Ifd35529b44c957737bf422127283c08e['h02ca2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01652] =  Ifd35529b44c957737bf422127283c08e['h02ca4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01653] =  Ifd35529b44c957737bf422127283c08e['h02ca6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01654] =  Ifd35529b44c957737bf422127283c08e['h02ca8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01655] =  Ifd35529b44c957737bf422127283c08e['h02caa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01656] =  Ifd35529b44c957737bf422127283c08e['h02cac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01657] =  Ifd35529b44c957737bf422127283c08e['h02cae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01658] =  Ifd35529b44c957737bf422127283c08e['h02cb0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01659] =  Ifd35529b44c957737bf422127283c08e['h02cb2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0165a] =  Ifd35529b44c957737bf422127283c08e['h02cb4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0165b] =  Ifd35529b44c957737bf422127283c08e['h02cb6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0165c] =  Ifd35529b44c957737bf422127283c08e['h02cb8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0165d] =  Ifd35529b44c957737bf422127283c08e['h02cba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0165e] =  Ifd35529b44c957737bf422127283c08e['h02cbc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0165f] =  Ifd35529b44c957737bf422127283c08e['h02cbe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01660] =  Ifd35529b44c957737bf422127283c08e['h02cc0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01661] =  Ifd35529b44c957737bf422127283c08e['h02cc2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01662] =  Ifd35529b44c957737bf422127283c08e['h02cc4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01663] =  Ifd35529b44c957737bf422127283c08e['h02cc6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01664] =  Ifd35529b44c957737bf422127283c08e['h02cc8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01665] =  Ifd35529b44c957737bf422127283c08e['h02cca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01666] =  Ifd35529b44c957737bf422127283c08e['h02ccc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01667] =  Ifd35529b44c957737bf422127283c08e['h02cce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01668] =  Ifd35529b44c957737bf422127283c08e['h02cd0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01669] =  Ifd35529b44c957737bf422127283c08e['h02cd2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0166a] =  Ifd35529b44c957737bf422127283c08e['h02cd4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0166b] =  Ifd35529b44c957737bf422127283c08e['h02cd6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0166c] =  Ifd35529b44c957737bf422127283c08e['h02cd8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0166d] =  Ifd35529b44c957737bf422127283c08e['h02cda] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0166e] =  Ifd35529b44c957737bf422127283c08e['h02cdc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0166f] =  Ifd35529b44c957737bf422127283c08e['h02cde] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01670] =  Ifd35529b44c957737bf422127283c08e['h02ce0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01671] =  Ifd35529b44c957737bf422127283c08e['h02ce2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01672] =  Ifd35529b44c957737bf422127283c08e['h02ce4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01673] =  Ifd35529b44c957737bf422127283c08e['h02ce6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01674] =  Ifd35529b44c957737bf422127283c08e['h02ce8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01675] =  Ifd35529b44c957737bf422127283c08e['h02cea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01676] =  Ifd35529b44c957737bf422127283c08e['h02cec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01677] =  Ifd35529b44c957737bf422127283c08e['h02cee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01678] =  Ifd35529b44c957737bf422127283c08e['h02cf0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01679] =  Ifd35529b44c957737bf422127283c08e['h02cf2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0167a] =  Ifd35529b44c957737bf422127283c08e['h02cf4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0167b] =  Ifd35529b44c957737bf422127283c08e['h02cf6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0167c] =  Ifd35529b44c957737bf422127283c08e['h02cf8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0167d] =  Ifd35529b44c957737bf422127283c08e['h02cfa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0167e] =  Ifd35529b44c957737bf422127283c08e['h02cfc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0167f] =  Ifd35529b44c957737bf422127283c08e['h02cfe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01680] =  Ifd35529b44c957737bf422127283c08e['h02d00] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01681] =  Ifd35529b44c957737bf422127283c08e['h02d02] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01682] =  Ifd35529b44c957737bf422127283c08e['h02d04] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01683] =  Ifd35529b44c957737bf422127283c08e['h02d06] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01684] =  Ifd35529b44c957737bf422127283c08e['h02d08] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01685] =  Ifd35529b44c957737bf422127283c08e['h02d0a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01686] =  Ifd35529b44c957737bf422127283c08e['h02d0c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01687] =  Ifd35529b44c957737bf422127283c08e['h02d0e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01688] =  Ifd35529b44c957737bf422127283c08e['h02d10] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01689] =  Ifd35529b44c957737bf422127283c08e['h02d12] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0168a] =  Ifd35529b44c957737bf422127283c08e['h02d14] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0168b] =  Ifd35529b44c957737bf422127283c08e['h02d16] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0168c] =  Ifd35529b44c957737bf422127283c08e['h02d18] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0168d] =  Ifd35529b44c957737bf422127283c08e['h02d1a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0168e] =  Ifd35529b44c957737bf422127283c08e['h02d1c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0168f] =  Ifd35529b44c957737bf422127283c08e['h02d1e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01690] =  Ifd35529b44c957737bf422127283c08e['h02d20] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01691] =  Ifd35529b44c957737bf422127283c08e['h02d22] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01692] =  Ifd35529b44c957737bf422127283c08e['h02d24] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01693] =  Ifd35529b44c957737bf422127283c08e['h02d26] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01694] =  Ifd35529b44c957737bf422127283c08e['h02d28] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01695] =  Ifd35529b44c957737bf422127283c08e['h02d2a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01696] =  Ifd35529b44c957737bf422127283c08e['h02d2c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01697] =  Ifd35529b44c957737bf422127283c08e['h02d2e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01698] =  Ifd35529b44c957737bf422127283c08e['h02d30] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01699] =  Ifd35529b44c957737bf422127283c08e['h02d32] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0169a] =  Ifd35529b44c957737bf422127283c08e['h02d34] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0169b] =  Ifd35529b44c957737bf422127283c08e['h02d36] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0169c] =  Ifd35529b44c957737bf422127283c08e['h02d38] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0169d] =  Ifd35529b44c957737bf422127283c08e['h02d3a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0169e] =  Ifd35529b44c957737bf422127283c08e['h02d3c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0169f] =  Ifd35529b44c957737bf422127283c08e['h02d3e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016a0] =  Ifd35529b44c957737bf422127283c08e['h02d40] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016a1] =  Ifd35529b44c957737bf422127283c08e['h02d42] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016a2] =  Ifd35529b44c957737bf422127283c08e['h02d44] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016a3] =  Ifd35529b44c957737bf422127283c08e['h02d46] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016a4] =  Ifd35529b44c957737bf422127283c08e['h02d48] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016a5] =  Ifd35529b44c957737bf422127283c08e['h02d4a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016a6] =  Ifd35529b44c957737bf422127283c08e['h02d4c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016a7] =  Ifd35529b44c957737bf422127283c08e['h02d4e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016a8] =  Ifd35529b44c957737bf422127283c08e['h02d50] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016a9] =  Ifd35529b44c957737bf422127283c08e['h02d52] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016aa] =  Ifd35529b44c957737bf422127283c08e['h02d54] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016ab] =  Ifd35529b44c957737bf422127283c08e['h02d56] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016ac] =  Ifd35529b44c957737bf422127283c08e['h02d58] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016ad] =  Ifd35529b44c957737bf422127283c08e['h02d5a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016ae] =  Ifd35529b44c957737bf422127283c08e['h02d5c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016af] =  Ifd35529b44c957737bf422127283c08e['h02d5e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016b0] =  Ifd35529b44c957737bf422127283c08e['h02d60] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016b1] =  Ifd35529b44c957737bf422127283c08e['h02d62] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016b2] =  Ifd35529b44c957737bf422127283c08e['h02d64] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016b3] =  Ifd35529b44c957737bf422127283c08e['h02d66] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016b4] =  Ifd35529b44c957737bf422127283c08e['h02d68] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016b5] =  Ifd35529b44c957737bf422127283c08e['h02d6a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016b6] =  Ifd35529b44c957737bf422127283c08e['h02d6c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016b7] =  Ifd35529b44c957737bf422127283c08e['h02d6e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016b8] =  Ifd35529b44c957737bf422127283c08e['h02d70] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016b9] =  Ifd35529b44c957737bf422127283c08e['h02d72] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016ba] =  Ifd35529b44c957737bf422127283c08e['h02d74] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016bb] =  Ifd35529b44c957737bf422127283c08e['h02d76] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016bc] =  Ifd35529b44c957737bf422127283c08e['h02d78] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016bd] =  Ifd35529b44c957737bf422127283c08e['h02d7a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016be] =  Ifd35529b44c957737bf422127283c08e['h02d7c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016bf] =  Ifd35529b44c957737bf422127283c08e['h02d7e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016c0] =  Ifd35529b44c957737bf422127283c08e['h02d80] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016c1] =  Ifd35529b44c957737bf422127283c08e['h02d82] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016c2] =  Ifd35529b44c957737bf422127283c08e['h02d84] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016c3] =  Ifd35529b44c957737bf422127283c08e['h02d86] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016c4] =  Ifd35529b44c957737bf422127283c08e['h02d88] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016c5] =  Ifd35529b44c957737bf422127283c08e['h02d8a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016c6] =  Ifd35529b44c957737bf422127283c08e['h02d8c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016c7] =  Ifd35529b44c957737bf422127283c08e['h02d8e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016c8] =  Ifd35529b44c957737bf422127283c08e['h02d90] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016c9] =  Ifd35529b44c957737bf422127283c08e['h02d92] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016ca] =  Ifd35529b44c957737bf422127283c08e['h02d94] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016cb] =  Ifd35529b44c957737bf422127283c08e['h02d96] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016cc] =  Ifd35529b44c957737bf422127283c08e['h02d98] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016cd] =  Ifd35529b44c957737bf422127283c08e['h02d9a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016ce] =  Ifd35529b44c957737bf422127283c08e['h02d9c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016cf] =  Ifd35529b44c957737bf422127283c08e['h02d9e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016d0] =  Ifd35529b44c957737bf422127283c08e['h02da0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016d1] =  Ifd35529b44c957737bf422127283c08e['h02da2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016d2] =  Ifd35529b44c957737bf422127283c08e['h02da4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016d3] =  Ifd35529b44c957737bf422127283c08e['h02da6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016d4] =  Ifd35529b44c957737bf422127283c08e['h02da8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016d5] =  Ifd35529b44c957737bf422127283c08e['h02daa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016d6] =  Ifd35529b44c957737bf422127283c08e['h02dac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016d7] =  Ifd35529b44c957737bf422127283c08e['h02dae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016d8] =  Ifd35529b44c957737bf422127283c08e['h02db0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016d9] =  Ifd35529b44c957737bf422127283c08e['h02db2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016da] =  Ifd35529b44c957737bf422127283c08e['h02db4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016db] =  Ifd35529b44c957737bf422127283c08e['h02db6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016dc] =  Ifd35529b44c957737bf422127283c08e['h02db8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016dd] =  Ifd35529b44c957737bf422127283c08e['h02dba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016de] =  Ifd35529b44c957737bf422127283c08e['h02dbc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016df] =  Ifd35529b44c957737bf422127283c08e['h02dbe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016e0] =  Ifd35529b44c957737bf422127283c08e['h02dc0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016e1] =  Ifd35529b44c957737bf422127283c08e['h02dc2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016e2] =  Ifd35529b44c957737bf422127283c08e['h02dc4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016e3] =  Ifd35529b44c957737bf422127283c08e['h02dc6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016e4] =  Ifd35529b44c957737bf422127283c08e['h02dc8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016e5] =  Ifd35529b44c957737bf422127283c08e['h02dca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016e6] =  Ifd35529b44c957737bf422127283c08e['h02dcc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016e7] =  Ifd35529b44c957737bf422127283c08e['h02dce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016e8] =  Ifd35529b44c957737bf422127283c08e['h02dd0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016e9] =  Ifd35529b44c957737bf422127283c08e['h02dd2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016ea] =  Ifd35529b44c957737bf422127283c08e['h02dd4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016eb] =  Ifd35529b44c957737bf422127283c08e['h02dd6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016ec] =  Ifd35529b44c957737bf422127283c08e['h02dd8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016ed] =  Ifd35529b44c957737bf422127283c08e['h02dda] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016ee] =  Ifd35529b44c957737bf422127283c08e['h02ddc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016ef] =  Ifd35529b44c957737bf422127283c08e['h02dde] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016f0] =  Ifd35529b44c957737bf422127283c08e['h02de0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016f1] =  Ifd35529b44c957737bf422127283c08e['h02de2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016f2] =  Ifd35529b44c957737bf422127283c08e['h02de4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016f3] =  Ifd35529b44c957737bf422127283c08e['h02de6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016f4] =  Ifd35529b44c957737bf422127283c08e['h02de8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016f5] =  Ifd35529b44c957737bf422127283c08e['h02dea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016f6] =  Ifd35529b44c957737bf422127283c08e['h02dec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016f7] =  Ifd35529b44c957737bf422127283c08e['h02dee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016f8] =  Ifd35529b44c957737bf422127283c08e['h02df0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016f9] =  Ifd35529b44c957737bf422127283c08e['h02df2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016fa] =  Ifd35529b44c957737bf422127283c08e['h02df4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016fb] =  Ifd35529b44c957737bf422127283c08e['h02df6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016fc] =  Ifd35529b44c957737bf422127283c08e['h02df8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016fd] =  Ifd35529b44c957737bf422127283c08e['h02dfa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016fe] =  Ifd35529b44c957737bf422127283c08e['h02dfc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h016ff] =  Ifd35529b44c957737bf422127283c08e['h02dfe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01700] =  Ifd35529b44c957737bf422127283c08e['h02e00] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01701] =  Ifd35529b44c957737bf422127283c08e['h02e02] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01702] =  Ifd35529b44c957737bf422127283c08e['h02e04] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01703] =  Ifd35529b44c957737bf422127283c08e['h02e06] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01704] =  Ifd35529b44c957737bf422127283c08e['h02e08] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01705] =  Ifd35529b44c957737bf422127283c08e['h02e0a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01706] =  Ifd35529b44c957737bf422127283c08e['h02e0c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01707] =  Ifd35529b44c957737bf422127283c08e['h02e0e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01708] =  Ifd35529b44c957737bf422127283c08e['h02e10] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01709] =  Ifd35529b44c957737bf422127283c08e['h02e12] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0170a] =  Ifd35529b44c957737bf422127283c08e['h02e14] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0170b] =  Ifd35529b44c957737bf422127283c08e['h02e16] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0170c] =  Ifd35529b44c957737bf422127283c08e['h02e18] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0170d] =  Ifd35529b44c957737bf422127283c08e['h02e1a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0170e] =  Ifd35529b44c957737bf422127283c08e['h02e1c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0170f] =  Ifd35529b44c957737bf422127283c08e['h02e1e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01710] =  Ifd35529b44c957737bf422127283c08e['h02e20] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01711] =  Ifd35529b44c957737bf422127283c08e['h02e22] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01712] =  Ifd35529b44c957737bf422127283c08e['h02e24] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01713] =  Ifd35529b44c957737bf422127283c08e['h02e26] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01714] =  Ifd35529b44c957737bf422127283c08e['h02e28] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01715] =  Ifd35529b44c957737bf422127283c08e['h02e2a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01716] =  Ifd35529b44c957737bf422127283c08e['h02e2c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01717] =  Ifd35529b44c957737bf422127283c08e['h02e2e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01718] =  Ifd35529b44c957737bf422127283c08e['h02e30] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01719] =  Ifd35529b44c957737bf422127283c08e['h02e32] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0171a] =  Ifd35529b44c957737bf422127283c08e['h02e34] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0171b] =  Ifd35529b44c957737bf422127283c08e['h02e36] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0171c] =  Ifd35529b44c957737bf422127283c08e['h02e38] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0171d] =  Ifd35529b44c957737bf422127283c08e['h02e3a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0171e] =  Ifd35529b44c957737bf422127283c08e['h02e3c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0171f] =  Ifd35529b44c957737bf422127283c08e['h02e3e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01720] =  Ifd35529b44c957737bf422127283c08e['h02e40] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01721] =  Ifd35529b44c957737bf422127283c08e['h02e42] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01722] =  Ifd35529b44c957737bf422127283c08e['h02e44] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01723] =  Ifd35529b44c957737bf422127283c08e['h02e46] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01724] =  Ifd35529b44c957737bf422127283c08e['h02e48] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01725] =  Ifd35529b44c957737bf422127283c08e['h02e4a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01726] =  Ifd35529b44c957737bf422127283c08e['h02e4c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01727] =  Ifd35529b44c957737bf422127283c08e['h02e4e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01728] =  Ifd35529b44c957737bf422127283c08e['h02e50] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01729] =  Ifd35529b44c957737bf422127283c08e['h02e52] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0172a] =  Ifd35529b44c957737bf422127283c08e['h02e54] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0172b] =  Ifd35529b44c957737bf422127283c08e['h02e56] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0172c] =  Ifd35529b44c957737bf422127283c08e['h02e58] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0172d] =  Ifd35529b44c957737bf422127283c08e['h02e5a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0172e] =  Ifd35529b44c957737bf422127283c08e['h02e5c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0172f] =  Ifd35529b44c957737bf422127283c08e['h02e5e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01730] =  Ifd35529b44c957737bf422127283c08e['h02e60] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01731] =  Ifd35529b44c957737bf422127283c08e['h02e62] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01732] =  Ifd35529b44c957737bf422127283c08e['h02e64] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01733] =  Ifd35529b44c957737bf422127283c08e['h02e66] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01734] =  Ifd35529b44c957737bf422127283c08e['h02e68] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01735] =  Ifd35529b44c957737bf422127283c08e['h02e6a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01736] =  Ifd35529b44c957737bf422127283c08e['h02e6c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01737] =  Ifd35529b44c957737bf422127283c08e['h02e6e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01738] =  Ifd35529b44c957737bf422127283c08e['h02e70] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01739] =  Ifd35529b44c957737bf422127283c08e['h02e72] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0173a] =  Ifd35529b44c957737bf422127283c08e['h02e74] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0173b] =  Ifd35529b44c957737bf422127283c08e['h02e76] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0173c] =  Ifd35529b44c957737bf422127283c08e['h02e78] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0173d] =  Ifd35529b44c957737bf422127283c08e['h02e7a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0173e] =  Ifd35529b44c957737bf422127283c08e['h02e7c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0173f] =  Ifd35529b44c957737bf422127283c08e['h02e7e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01740] =  Ifd35529b44c957737bf422127283c08e['h02e80] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01741] =  Ifd35529b44c957737bf422127283c08e['h02e82] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01742] =  Ifd35529b44c957737bf422127283c08e['h02e84] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01743] =  Ifd35529b44c957737bf422127283c08e['h02e86] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01744] =  Ifd35529b44c957737bf422127283c08e['h02e88] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01745] =  Ifd35529b44c957737bf422127283c08e['h02e8a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01746] =  Ifd35529b44c957737bf422127283c08e['h02e8c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01747] =  Ifd35529b44c957737bf422127283c08e['h02e8e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01748] =  Ifd35529b44c957737bf422127283c08e['h02e90] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01749] =  Ifd35529b44c957737bf422127283c08e['h02e92] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0174a] =  Ifd35529b44c957737bf422127283c08e['h02e94] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0174b] =  Ifd35529b44c957737bf422127283c08e['h02e96] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0174c] =  Ifd35529b44c957737bf422127283c08e['h02e98] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0174d] =  Ifd35529b44c957737bf422127283c08e['h02e9a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0174e] =  Ifd35529b44c957737bf422127283c08e['h02e9c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0174f] =  Ifd35529b44c957737bf422127283c08e['h02e9e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01750] =  Ifd35529b44c957737bf422127283c08e['h02ea0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01751] =  Ifd35529b44c957737bf422127283c08e['h02ea2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01752] =  Ifd35529b44c957737bf422127283c08e['h02ea4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01753] =  Ifd35529b44c957737bf422127283c08e['h02ea6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01754] =  Ifd35529b44c957737bf422127283c08e['h02ea8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01755] =  Ifd35529b44c957737bf422127283c08e['h02eaa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01756] =  Ifd35529b44c957737bf422127283c08e['h02eac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01757] =  Ifd35529b44c957737bf422127283c08e['h02eae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01758] =  Ifd35529b44c957737bf422127283c08e['h02eb0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01759] =  Ifd35529b44c957737bf422127283c08e['h02eb2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0175a] =  Ifd35529b44c957737bf422127283c08e['h02eb4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0175b] =  Ifd35529b44c957737bf422127283c08e['h02eb6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0175c] =  Ifd35529b44c957737bf422127283c08e['h02eb8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0175d] =  Ifd35529b44c957737bf422127283c08e['h02eba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0175e] =  Ifd35529b44c957737bf422127283c08e['h02ebc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0175f] =  Ifd35529b44c957737bf422127283c08e['h02ebe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01760] =  Ifd35529b44c957737bf422127283c08e['h02ec0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01761] =  Ifd35529b44c957737bf422127283c08e['h02ec2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01762] =  Ifd35529b44c957737bf422127283c08e['h02ec4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01763] =  Ifd35529b44c957737bf422127283c08e['h02ec6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01764] =  Ifd35529b44c957737bf422127283c08e['h02ec8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01765] =  Ifd35529b44c957737bf422127283c08e['h02eca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01766] =  Ifd35529b44c957737bf422127283c08e['h02ecc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01767] =  Ifd35529b44c957737bf422127283c08e['h02ece] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01768] =  Ifd35529b44c957737bf422127283c08e['h02ed0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01769] =  Ifd35529b44c957737bf422127283c08e['h02ed2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0176a] =  Ifd35529b44c957737bf422127283c08e['h02ed4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0176b] =  Ifd35529b44c957737bf422127283c08e['h02ed6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0176c] =  Ifd35529b44c957737bf422127283c08e['h02ed8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0176d] =  Ifd35529b44c957737bf422127283c08e['h02eda] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0176e] =  Ifd35529b44c957737bf422127283c08e['h02edc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0176f] =  Ifd35529b44c957737bf422127283c08e['h02ede] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01770] =  Ifd35529b44c957737bf422127283c08e['h02ee0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01771] =  Ifd35529b44c957737bf422127283c08e['h02ee2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01772] =  Ifd35529b44c957737bf422127283c08e['h02ee4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01773] =  Ifd35529b44c957737bf422127283c08e['h02ee6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01774] =  Ifd35529b44c957737bf422127283c08e['h02ee8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01775] =  Ifd35529b44c957737bf422127283c08e['h02eea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01776] =  Ifd35529b44c957737bf422127283c08e['h02eec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01777] =  Ifd35529b44c957737bf422127283c08e['h02eee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01778] =  Ifd35529b44c957737bf422127283c08e['h02ef0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01779] =  Ifd35529b44c957737bf422127283c08e['h02ef2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0177a] =  Ifd35529b44c957737bf422127283c08e['h02ef4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0177b] =  Ifd35529b44c957737bf422127283c08e['h02ef6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0177c] =  Ifd35529b44c957737bf422127283c08e['h02ef8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0177d] =  Ifd35529b44c957737bf422127283c08e['h02efa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0177e] =  Ifd35529b44c957737bf422127283c08e['h02efc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0177f] =  Ifd35529b44c957737bf422127283c08e['h02efe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01780] =  Ifd35529b44c957737bf422127283c08e['h02f00] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01781] =  Ifd35529b44c957737bf422127283c08e['h02f02] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01782] =  Ifd35529b44c957737bf422127283c08e['h02f04] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01783] =  Ifd35529b44c957737bf422127283c08e['h02f06] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01784] =  Ifd35529b44c957737bf422127283c08e['h02f08] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01785] =  Ifd35529b44c957737bf422127283c08e['h02f0a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01786] =  Ifd35529b44c957737bf422127283c08e['h02f0c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01787] =  Ifd35529b44c957737bf422127283c08e['h02f0e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01788] =  Ifd35529b44c957737bf422127283c08e['h02f10] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01789] =  Ifd35529b44c957737bf422127283c08e['h02f12] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0178a] =  Ifd35529b44c957737bf422127283c08e['h02f14] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0178b] =  Ifd35529b44c957737bf422127283c08e['h02f16] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0178c] =  Ifd35529b44c957737bf422127283c08e['h02f18] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0178d] =  Ifd35529b44c957737bf422127283c08e['h02f1a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0178e] =  Ifd35529b44c957737bf422127283c08e['h02f1c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0178f] =  Ifd35529b44c957737bf422127283c08e['h02f1e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01790] =  Ifd35529b44c957737bf422127283c08e['h02f20] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01791] =  Ifd35529b44c957737bf422127283c08e['h02f22] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01792] =  Ifd35529b44c957737bf422127283c08e['h02f24] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01793] =  Ifd35529b44c957737bf422127283c08e['h02f26] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01794] =  Ifd35529b44c957737bf422127283c08e['h02f28] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01795] =  Ifd35529b44c957737bf422127283c08e['h02f2a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01796] =  Ifd35529b44c957737bf422127283c08e['h02f2c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01797] =  Ifd35529b44c957737bf422127283c08e['h02f2e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01798] =  Ifd35529b44c957737bf422127283c08e['h02f30] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01799] =  Ifd35529b44c957737bf422127283c08e['h02f32] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0179a] =  Ifd35529b44c957737bf422127283c08e['h02f34] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0179b] =  Ifd35529b44c957737bf422127283c08e['h02f36] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0179c] =  Ifd35529b44c957737bf422127283c08e['h02f38] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0179d] =  Ifd35529b44c957737bf422127283c08e['h02f3a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0179e] =  Ifd35529b44c957737bf422127283c08e['h02f3c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0179f] =  Ifd35529b44c957737bf422127283c08e['h02f3e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017a0] =  Ifd35529b44c957737bf422127283c08e['h02f40] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017a1] =  Ifd35529b44c957737bf422127283c08e['h02f42] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017a2] =  Ifd35529b44c957737bf422127283c08e['h02f44] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017a3] =  Ifd35529b44c957737bf422127283c08e['h02f46] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017a4] =  Ifd35529b44c957737bf422127283c08e['h02f48] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017a5] =  Ifd35529b44c957737bf422127283c08e['h02f4a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017a6] =  Ifd35529b44c957737bf422127283c08e['h02f4c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017a7] =  Ifd35529b44c957737bf422127283c08e['h02f4e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017a8] =  Ifd35529b44c957737bf422127283c08e['h02f50] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017a9] =  Ifd35529b44c957737bf422127283c08e['h02f52] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017aa] =  Ifd35529b44c957737bf422127283c08e['h02f54] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017ab] =  Ifd35529b44c957737bf422127283c08e['h02f56] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017ac] =  Ifd35529b44c957737bf422127283c08e['h02f58] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017ad] =  Ifd35529b44c957737bf422127283c08e['h02f5a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017ae] =  Ifd35529b44c957737bf422127283c08e['h02f5c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017af] =  Ifd35529b44c957737bf422127283c08e['h02f5e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017b0] =  Ifd35529b44c957737bf422127283c08e['h02f60] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017b1] =  Ifd35529b44c957737bf422127283c08e['h02f62] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017b2] =  Ifd35529b44c957737bf422127283c08e['h02f64] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017b3] =  Ifd35529b44c957737bf422127283c08e['h02f66] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017b4] =  Ifd35529b44c957737bf422127283c08e['h02f68] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017b5] =  Ifd35529b44c957737bf422127283c08e['h02f6a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017b6] =  Ifd35529b44c957737bf422127283c08e['h02f6c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017b7] =  Ifd35529b44c957737bf422127283c08e['h02f6e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017b8] =  Ifd35529b44c957737bf422127283c08e['h02f70] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017b9] =  Ifd35529b44c957737bf422127283c08e['h02f72] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017ba] =  Ifd35529b44c957737bf422127283c08e['h02f74] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017bb] =  Ifd35529b44c957737bf422127283c08e['h02f76] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017bc] =  Ifd35529b44c957737bf422127283c08e['h02f78] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017bd] =  Ifd35529b44c957737bf422127283c08e['h02f7a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017be] =  Ifd35529b44c957737bf422127283c08e['h02f7c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017bf] =  Ifd35529b44c957737bf422127283c08e['h02f7e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017c0] =  Ifd35529b44c957737bf422127283c08e['h02f80] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017c1] =  Ifd35529b44c957737bf422127283c08e['h02f82] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017c2] =  Ifd35529b44c957737bf422127283c08e['h02f84] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017c3] =  Ifd35529b44c957737bf422127283c08e['h02f86] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017c4] =  Ifd35529b44c957737bf422127283c08e['h02f88] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017c5] =  Ifd35529b44c957737bf422127283c08e['h02f8a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017c6] =  Ifd35529b44c957737bf422127283c08e['h02f8c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017c7] =  Ifd35529b44c957737bf422127283c08e['h02f8e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017c8] =  Ifd35529b44c957737bf422127283c08e['h02f90] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017c9] =  Ifd35529b44c957737bf422127283c08e['h02f92] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017ca] =  Ifd35529b44c957737bf422127283c08e['h02f94] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017cb] =  Ifd35529b44c957737bf422127283c08e['h02f96] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017cc] =  Ifd35529b44c957737bf422127283c08e['h02f98] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017cd] =  Ifd35529b44c957737bf422127283c08e['h02f9a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017ce] =  Ifd35529b44c957737bf422127283c08e['h02f9c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017cf] =  Ifd35529b44c957737bf422127283c08e['h02f9e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017d0] =  Ifd35529b44c957737bf422127283c08e['h02fa0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017d1] =  Ifd35529b44c957737bf422127283c08e['h02fa2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017d2] =  Ifd35529b44c957737bf422127283c08e['h02fa4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017d3] =  Ifd35529b44c957737bf422127283c08e['h02fa6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017d4] =  Ifd35529b44c957737bf422127283c08e['h02fa8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017d5] =  Ifd35529b44c957737bf422127283c08e['h02faa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017d6] =  Ifd35529b44c957737bf422127283c08e['h02fac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017d7] =  Ifd35529b44c957737bf422127283c08e['h02fae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017d8] =  Ifd35529b44c957737bf422127283c08e['h02fb0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017d9] =  Ifd35529b44c957737bf422127283c08e['h02fb2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017da] =  Ifd35529b44c957737bf422127283c08e['h02fb4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017db] =  Ifd35529b44c957737bf422127283c08e['h02fb6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017dc] =  Ifd35529b44c957737bf422127283c08e['h02fb8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017dd] =  Ifd35529b44c957737bf422127283c08e['h02fba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017de] =  Ifd35529b44c957737bf422127283c08e['h02fbc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017df] =  Ifd35529b44c957737bf422127283c08e['h02fbe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017e0] =  Ifd35529b44c957737bf422127283c08e['h02fc0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017e1] =  Ifd35529b44c957737bf422127283c08e['h02fc2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017e2] =  Ifd35529b44c957737bf422127283c08e['h02fc4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017e3] =  Ifd35529b44c957737bf422127283c08e['h02fc6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017e4] =  Ifd35529b44c957737bf422127283c08e['h02fc8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017e5] =  Ifd35529b44c957737bf422127283c08e['h02fca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017e6] =  Ifd35529b44c957737bf422127283c08e['h02fcc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017e7] =  Ifd35529b44c957737bf422127283c08e['h02fce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017e8] =  Ifd35529b44c957737bf422127283c08e['h02fd0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017e9] =  Ifd35529b44c957737bf422127283c08e['h02fd2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017ea] =  Ifd35529b44c957737bf422127283c08e['h02fd4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017eb] =  Ifd35529b44c957737bf422127283c08e['h02fd6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017ec] =  Ifd35529b44c957737bf422127283c08e['h02fd8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017ed] =  Ifd35529b44c957737bf422127283c08e['h02fda] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017ee] =  Ifd35529b44c957737bf422127283c08e['h02fdc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017ef] =  Ifd35529b44c957737bf422127283c08e['h02fde] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017f0] =  Ifd35529b44c957737bf422127283c08e['h02fe0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017f1] =  Ifd35529b44c957737bf422127283c08e['h02fe2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017f2] =  Ifd35529b44c957737bf422127283c08e['h02fe4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017f3] =  Ifd35529b44c957737bf422127283c08e['h02fe6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017f4] =  Ifd35529b44c957737bf422127283c08e['h02fe8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017f5] =  Ifd35529b44c957737bf422127283c08e['h02fea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017f6] =  Ifd35529b44c957737bf422127283c08e['h02fec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017f7] =  Ifd35529b44c957737bf422127283c08e['h02fee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017f8] =  Ifd35529b44c957737bf422127283c08e['h02ff0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017f9] =  Ifd35529b44c957737bf422127283c08e['h02ff2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017fa] =  Ifd35529b44c957737bf422127283c08e['h02ff4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017fb] =  Ifd35529b44c957737bf422127283c08e['h02ff6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017fc] =  Ifd35529b44c957737bf422127283c08e['h02ff8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017fd] =  Ifd35529b44c957737bf422127283c08e['h02ffa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017fe] =  Ifd35529b44c957737bf422127283c08e['h02ffc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h017ff] =  Ifd35529b44c957737bf422127283c08e['h02ffe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01800] =  Ifd35529b44c957737bf422127283c08e['h03000] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01801] =  Ifd35529b44c957737bf422127283c08e['h03002] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01802] =  Ifd35529b44c957737bf422127283c08e['h03004] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01803] =  Ifd35529b44c957737bf422127283c08e['h03006] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01804] =  Ifd35529b44c957737bf422127283c08e['h03008] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01805] =  Ifd35529b44c957737bf422127283c08e['h0300a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01806] =  Ifd35529b44c957737bf422127283c08e['h0300c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01807] =  Ifd35529b44c957737bf422127283c08e['h0300e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01808] =  Ifd35529b44c957737bf422127283c08e['h03010] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01809] =  Ifd35529b44c957737bf422127283c08e['h03012] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0180a] =  Ifd35529b44c957737bf422127283c08e['h03014] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0180b] =  Ifd35529b44c957737bf422127283c08e['h03016] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0180c] =  Ifd35529b44c957737bf422127283c08e['h03018] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0180d] =  Ifd35529b44c957737bf422127283c08e['h0301a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0180e] =  Ifd35529b44c957737bf422127283c08e['h0301c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0180f] =  Ifd35529b44c957737bf422127283c08e['h0301e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01810] =  Ifd35529b44c957737bf422127283c08e['h03020] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01811] =  Ifd35529b44c957737bf422127283c08e['h03022] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01812] =  Ifd35529b44c957737bf422127283c08e['h03024] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01813] =  Ifd35529b44c957737bf422127283c08e['h03026] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01814] =  Ifd35529b44c957737bf422127283c08e['h03028] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01815] =  Ifd35529b44c957737bf422127283c08e['h0302a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01816] =  Ifd35529b44c957737bf422127283c08e['h0302c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01817] =  Ifd35529b44c957737bf422127283c08e['h0302e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01818] =  Ifd35529b44c957737bf422127283c08e['h03030] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01819] =  Ifd35529b44c957737bf422127283c08e['h03032] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0181a] =  Ifd35529b44c957737bf422127283c08e['h03034] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0181b] =  Ifd35529b44c957737bf422127283c08e['h03036] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0181c] =  Ifd35529b44c957737bf422127283c08e['h03038] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0181d] =  Ifd35529b44c957737bf422127283c08e['h0303a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0181e] =  Ifd35529b44c957737bf422127283c08e['h0303c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0181f] =  Ifd35529b44c957737bf422127283c08e['h0303e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01820] =  Ifd35529b44c957737bf422127283c08e['h03040] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01821] =  Ifd35529b44c957737bf422127283c08e['h03042] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01822] =  Ifd35529b44c957737bf422127283c08e['h03044] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01823] =  Ifd35529b44c957737bf422127283c08e['h03046] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01824] =  Ifd35529b44c957737bf422127283c08e['h03048] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01825] =  Ifd35529b44c957737bf422127283c08e['h0304a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01826] =  Ifd35529b44c957737bf422127283c08e['h0304c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01827] =  Ifd35529b44c957737bf422127283c08e['h0304e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01828] =  Ifd35529b44c957737bf422127283c08e['h03050] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01829] =  Ifd35529b44c957737bf422127283c08e['h03052] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0182a] =  Ifd35529b44c957737bf422127283c08e['h03054] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0182b] =  Ifd35529b44c957737bf422127283c08e['h03056] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0182c] =  Ifd35529b44c957737bf422127283c08e['h03058] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0182d] =  Ifd35529b44c957737bf422127283c08e['h0305a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0182e] =  Ifd35529b44c957737bf422127283c08e['h0305c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0182f] =  Ifd35529b44c957737bf422127283c08e['h0305e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01830] =  Ifd35529b44c957737bf422127283c08e['h03060] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01831] =  Ifd35529b44c957737bf422127283c08e['h03062] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01832] =  Ifd35529b44c957737bf422127283c08e['h03064] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01833] =  Ifd35529b44c957737bf422127283c08e['h03066] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01834] =  Ifd35529b44c957737bf422127283c08e['h03068] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01835] =  Ifd35529b44c957737bf422127283c08e['h0306a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01836] =  Ifd35529b44c957737bf422127283c08e['h0306c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01837] =  Ifd35529b44c957737bf422127283c08e['h0306e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01838] =  Ifd35529b44c957737bf422127283c08e['h03070] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01839] =  Ifd35529b44c957737bf422127283c08e['h03072] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0183a] =  Ifd35529b44c957737bf422127283c08e['h03074] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0183b] =  Ifd35529b44c957737bf422127283c08e['h03076] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0183c] =  Ifd35529b44c957737bf422127283c08e['h03078] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0183d] =  Ifd35529b44c957737bf422127283c08e['h0307a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0183e] =  Ifd35529b44c957737bf422127283c08e['h0307c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0183f] =  Ifd35529b44c957737bf422127283c08e['h0307e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01840] =  Ifd35529b44c957737bf422127283c08e['h03080] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01841] =  Ifd35529b44c957737bf422127283c08e['h03082] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01842] =  Ifd35529b44c957737bf422127283c08e['h03084] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01843] =  Ifd35529b44c957737bf422127283c08e['h03086] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01844] =  Ifd35529b44c957737bf422127283c08e['h03088] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01845] =  Ifd35529b44c957737bf422127283c08e['h0308a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01846] =  Ifd35529b44c957737bf422127283c08e['h0308c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01847] =  Ifd35529b44c957737bf422127283c08e['h0308e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01848] =  Ifd35529b44c957737bf422127283c08e['h03090] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01849] =  Ifd35529b44c957737bf422127283c08e['h03092] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0184a] =  Ifd35529b44c957737bf422127283c08e['h03094] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0184b] =  Ifd35529b44c957737bf422127283c08e['h03096] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0184c] =  Ifd35529b44c957737bf422127283c08e['h03098] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0184d] =  Ifd35529b44c957737bf422127283c08e['h0309a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0184e] =  Ifd35529b44c957737bf422127283c08e['h0309c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0184f] =  Ifd35529b44c957737bf422127283c08e['h0309e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01850] =  Ifd35529b44c957737bf422127283c08e['h030a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01851] =  Ifd35529b44c957737bf422127283c08e['h030a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01852] =  Ifd35529b44c957737bf422127283c08e['h030a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01853] =  Ifd35529b44c957737bf422127283c08e['h030a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01854] =  Ifd35529b44c957737bf422127283c08e['h030a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01855] =  Ifd35529b44c957737bf422127283c08e['h030aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01856] =  Ifd35529b44c957737bf422127283c08e['h030ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01857] =  Ifd35529b44c957737bf422127283c08e['h030ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01858] =  Ifd35529b44c957737bf422127283c08e['h030b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01859] =  Ifd35529b44c957737bf422127283c08e['h030b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0185a] =  Ifd35529b44c957737bf422127283c08e['h030b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0185b] =  Ifd35529b44c957737bf422127283c08e['h030b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0185c] =  Ifd35529b44c957737bf422127283c08e['h030b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0185d] =  Ifd35529b44c957737bf422127283c08e['h030ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0185e] =  Ifd35529b44c957737bf422127283c08e['h030bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0185f] =  Ifd35529b44c957737bf422127283c08e['h030be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01860] =  Ifd35529b44c957737bf422127283c08e['h030c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01861] =  Ifd35529b44c957737bf422127283c08e['h030c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01862] =  Ifd35529b44c957737bf422127283c08e['h030c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01863] =  Ifd35529b44c957737bf422127283c08e['h030c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01864] =  Ifd35529b44c957737bf422127283c08e['h030c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01865] =  Ifd35529b44c957737bf422127283c08e['h030ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01866] =  Ifd35529b44c957737bf422127283c08e['h030cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01867] =  Ifd35529b44c957737bf422127283c08e['h030ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01868] =  Ifd35529b44c957737bf422127283c08e['h030d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01869] =  Ifd35529b44c957737bf422127283c08e['h030d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0186a] =  Ifd35529b44c957737bf422127283c08e['h030d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0186b] =  Ifd35529b44c957737bf422127283c08e['h030d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0186c] =  Ifd35529b44c957737bf422127283c08e['h030d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0186d] =  Ifd35529b44c957737bf422127283c08e['h030da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0186e] =  Ifd35529b44c957737bf422127283c08e['h030dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0186f] =  Ifd35529b44c957737bf422127283c08e['h030de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01870] =  Ifd35529b44c957737bf422127283c08e['h030e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01871] =  Ifd35529b44c957737bf422127283c08e['h030e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01872] =  Ifd35529b44c957737bf422127283c08e['h030e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01873] =  Ifd35529b44c957737bf422127283c08e['h030e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01874] =  Ifd35529b44c957737bf422127283c08e['h030e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01875] =  Ifd35529b44c957737bf422127283c08e['h030ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01876] =  Ifd35529b44c957737bf422127283c08e['h030ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01877] =  Ifd35529b44c957737bf422127283c08e['h030ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01878] =  Ifd35529b44c957737bf422127283c08e['h030f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01879] =  Ifd35529b44c957737bf422127283c08e['h030f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0187a] =  Ifd35529b44c957737bf422127283c08e['h030f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0187b] =  Ifd35529b44c957737bf422127283c08e['h030f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0187c] =  Ifd35529b44c957737bf422127283c08e['h030f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0187d] =  Ifd35529b44c957737bf422127283c08e['h030fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0187e] =  Ifd35529b44c957737bf422127283c08e['h030fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0187f] =  Ifd35529b44c957737bf422127283c08e['h030fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01880] =  Ifd35529b44c957737bf422127283c08e['h03100] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01881] =  Ifd35529b44c957737bf422127283c08e['h03102] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01882] =  Ifd35529b44c957737bf422127283c08e['h03104] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01883] =  Ifd35529b44c957737bf422127283c08e['h03106] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01884] =  Ifd35529b44c957737bf422127283c08e['h03108] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01885] =  Ifd35529b44c957737bf422127283c08e['h0310a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01886] =  Ifd35529b44c957737bf422127283c08e['h0310c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01887] =  Ifd35529b44c957737bf422127283c08e['h0310e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01888] =  Ifd35529b44c957737bf422127283c08e['h03110] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01889] =  Ifd35529b44c957737bf422127283c08e['h03112] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0188a] =  Ifd35529b44c957737bf422127283c08e['h03114] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0188b] =  Ifd35529b44c957737bf422127283c08e['h03116] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0188c] =  Ifd35529b44c957737bf422127283c08e['h03118] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0188d] =  Ifd35529b44c957737bf422127283c08e['h0311a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0188e] =  Ifd35529b44c957737bf422127283c08e['h0311c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0188f] =  Ifd35529b44c957737bf422127283c08e['h0311e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01890] =  Ifd35529b44c957737bf422127283c08e['h03120] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01891] =  Ifd35529b44c957737bf422127283c08e['h03122] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01892] =  Ifd35529b44c957737bf422127283c08e['h03124] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01893] =  Ifd35529b44c957737bf422127283c08e['h03126] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01894] =  Ifd35529b44c957737bf422127283c08e['h03128] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01895] =  Ifd35529b44c957737bf422127283c08e['h0312a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01896] =  Ifd35529b44c957737bf422127283c08e['h0312c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01897] =  Ifd35529b44c957737bf422127283c08e['h0312e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01898] =  Ifd35529b44c957737bf422127283c08e['h03130] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01899] =  Ifd35529b44c957737bf422127283c08e['h03132] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0189a] =  Ifd35529b44c957737bf422127283c08e['h03134] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0189b] =  Ifd35529b44c957737bf422127283c08e['h03136] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0189c] =  Ifd35529b44c957737bf422127283c08e['h03138] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0189d] =  Ifd35529b44c957737bf422127283c08e['h0313a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0189e] =  Ifd35529b44c957737bf422127283c08e['h0313c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0189f] =  Ifd35529b44c957737bf422127283c08e['h0313e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018a0] =  Ifd35529b44c957737bf422127283c08e['h03140] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018a1] =  Ifd35529b44c957737bf422127283c08e['h03142] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018a2] =  Ifd35529b44c957737bf422127283c08e['h03144] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018a3] =  Ifd35529b44c957737bf422127283c08e['h03146] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018a4] =  Ifd35529b44c957737bf422127283c08e['h03148] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018a5] =  Ifd35529b44c957737bf422127283c08e['h0314a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018a6] =  Ifd35529b44c957737bf422127283c08e['h0314c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018a7] =  Ifd35529b44c957737bf422127283c08e['h0314e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018a8] =  Ifd35529b44c957737bf422127283c08e['h03150] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018a9] =  Ifd35529b44c957737bf422127283c08e['h03152] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018aa] =  Ifd35529b44c957737bf422127283c08e['h03154] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018ab] =  Ifd35529b44c957737bf422127283c08e['h03156] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018ac] =  Ifd35529b44c957737bf422127283c08e['h03158] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018ad] =  Ifd35529b44c957737bf422127283c08e['h0315a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018ae] =  Ifd35529b44c957737bf422127283c08e['h0315c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018af] =  Ifd35529b44c957737bf422127283c08e['h0315e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018b0] =  Ifd35529b44c957737bf422127283c08e['h03160] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018b1] =  Ifd35529b44c957737bf422127283c08e['h03162] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018b2] =  Ifd35529b44c957737bf422127283c08e['h03164] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018b3] =  Ifd35529b44c957737bf422127283c08e['h03166] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018b4] =  Ifd35529b44c957737bf422127283c08e['h03168] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018b5] =  Ifd35529b44c957737bf422127283c08e['h0316a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018b6] =  Ifd35529b44c957737bf422127283c08e['h0316c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018b7] =  Ifd35529b44c957737bf422127283c08e['h0316e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018b8] =  Ifd35529b44c957737bf422127283c08e['h03170] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018b9] =  Ifd35529b44c957737bf422127283c08e['h03172] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018ba] =  Ifd35529b44c957737bf422127283c08e['h03174] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018bb] =  Ifd35529b44c957737bf422127283c08e['h03176] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018bc] =  Ifd35529b44c957737bf422127283c08e['h03178] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018bd] =  Ifd35529b44c957737bf422127283c08e['h0317a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018be] =  Ifd35529b44c957737bf422127283c08e['h0317c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018bf] =  Ifd35529b44c957737bf422127283c08e['h0317e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018c0] =  Ifd35529b44c957737bf422127283c08e['h03180] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018c1] =  Ifd35529b44c957737bf422127283c08e['h03182] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018c2] =  Ifd35529b44c957737bf422127283c08e['h03184] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018c3] =  Ifd35529b44c957737bf422127283c08e['h03186] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018c4] =  Ifd35529b44c957737bf422127283c08e['h03188] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018c5] =  Ifd35529b44c957737bf422127283c08e['h0318a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018c6] =  Ifd35529b44c957737bf422127283c08e['h0318c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018c7] =  Ifd35529b44c957737bf422127283c08e['h0318e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018c8] =  Ifd35529b44c957737bf422127283c08e['h03190] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018c9] =  Ifd35529b44c957737bf422127283c08e['h03192] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018ca] =  Ifd35529b44c957737bf422127283c08e['h03194] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018cb] =  Ifd35529b44c957737bf422127283c08e['h03196] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018cc] =  Ifd35529b44c957737bf422127283c08e['h03198] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018cd] =  Ifd35529b44c957737bf422127283c08e['h0319a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018ce] =  Ifd35529b44c957737bf422127283c08e['h0319c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018cf] =  Ifd35529b44c957737bf422127283c08e['h0319e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018d0] =  Ifd35529b44c957737bf422127283c08e['h031a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018d1] =  Ifd35529b44c957737bf422127283c08e['h031a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018d2] =  Ifd35529b44c957737bf422127283c08e['h031a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018d3] =  Ifd35529b44c957737bf422127283c08e['h031a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018d4] =  Ifd35529b44c957737bf422127283c08e['h031a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018d5] =  Ifd35529b44c957737bf422127283c08e['h031aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018d6] =  Ifd35529b44c957737bf422127283c08e['h031ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018d7] =  Ifd35529b44c957737bf422127283c08e['h031ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018d8] =  Ifd35529b44c957737bf422127283c08e['h031b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018d9] =  Ifd35529b44c957737bf422127283c08e['h031b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018da] =  Ifd35529b44c957737bf422127283c08e['h031b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018db] =  Ifd35529b44c957737bf422127283c08e['h031b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018dc] =  Ifd35529b44c957737bf422127283c08e['h031b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018dd] =  Ifd35529b44c957737bf422127283c08e['h031ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018de] =  Ifd35529b44c957737bf422127283c08e['h031bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018df] =  Ifd35529b44c957737bf422127283c08e['h031be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018e0] =  Ifd35529b44c957737bf422127283c08e['h031c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018e1] =  Ifd35529b44c957737bf422127283c08e['h031c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018e2] =  Ifd35529b44c957737bf422127283c08e['h031c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018e3] =  Ifd35529b44c957737bf422127283c08e['h031c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018e4] =  Ifd35529b44c957737bf422127283c08e['h031c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018e5] =  Ifd35529b44c957737bf422127283c08e['h031ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018e6] =  Ifd35529b44c957737bf422127283c08e['h031cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018e7] =  Ifd35529b44c957737bf422127283c08e['h031ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018e8] =  Ifd35529b44c957737bf422127283c08e['h031d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018e9] =  Ifd35529b44c957737bf422127283c08e['h031d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018ea] =  Ifd35529b44c957737bf422127283c08e['h031d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018eb] =  Ifd35529b44c957737bf422127283c08e['h031d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018ec] =  Ifd35529b44c957737bf422127283c08e['h031d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018ed] =  Ifd35529b44c957737bf422127283c08e['h031da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018ee] =  Ifd35529b44c957737bf422127283c08e['h031dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018ef] =  Ifd35529b44c957737bf422127283c08e['h031de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018f0] =  Ifd35529b44c957737bf422127283c08e['h031e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018f1] =  Ifd35529b44c957737bf422127283c08e['h031e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018f2] =  Ifd35529b44c957737bf422127283c08e['h031e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018f3] =  Ifd35529b44c957737bf422127283c08e['h031e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018f4] =  Ifd35529b44c957737bf422127283c08e['h031e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018f5] =  Ifd35529b44c957737bf422127283c08e['h031ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018f6] =  Ifd35529b44c957737bf422127283c08e['h031ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018f7] =  Ifd35529b44c957737bf422127283c08e['h031ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018f8] =  Ifd35529b44c957737bf422127283c08e['h031f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018f9] =  Ifd35529b44c957737bf422127283c08e['h031f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018fa] =  Ifd35529b44c957737bf422127283c08e['h031f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018fb] =  Ifd35529b44c957737bf422127283c08e['h031f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018fc] =  Ifd35529b44c957737bf422127283c08e['h031f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018fd] =  Ifd35529b44c957737bf422127283c08e['h031fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018fe] =  Ifd35529b44c957737bf422127283c08e['h031fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h018ff] =  Ifd35529b44c957737bf422127283c08e['h031fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01900] =  Ifd35529b44c957737bf422127283c08e['h03200] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01901] =  Ifd35529b44c957737bf422127283c08e['h03202] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01902] =  Ifd35529b44c957737bf422127283c08e['h03204] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01903] =  Ifd35529b44c957737bf422127283c08e['h03206] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01904] =  Ifd35529b44c957737bf422127283c08e['h03208] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01905] =  Ifd35529b44c957737bf422127283c08e['h0320a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01906] =  Ifd35529b44c957737bf422127283c08e['h0320c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01907] =  Ifd35529b44c957737bf422127283c08e['h0320e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01908] =  Ifd35529b44c957737bf422127283c08e['h03210] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01909] =  Ifd35529b44c957737bf422127283c08e['h03212] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0190a] =  Ifd35529b44c957737bf422127283c08e['h03214] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0190b] =  Ifd35529b44c957737bf422127283c08e['h03216] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0190c] =  Ifd35529b44c957737bf422127283c08e['h03218] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0190d] =  Ifd35529b44c957737bf422127283c08e['h0321a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0190e] =  Ifd35529b44c957737bf422127283c08e['h0321c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0190f] =  Ifd35529b44c957737bf422127283c08e['h0321e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01910] =  Ifd35529b44c957737bf422127283c08e['h03220] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01911] =  Ifd35529b44c957737bf422127283c08e['h03222] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01912] =  Ifd35529b44c957737bf422127283c08e['h03224] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01913] =  Ifd35529b44c957737bf422127283c08e['h03226] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01914] =  Ifd35529b44c957737bf422127283c08e['h03228] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01915] =  Ifd35529b44c957737bf422127283c08e['h0322a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01916] =  Ifd35529b44c957737bf422127283c08e['h0322c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01917] =  Ifd35529b44c957737bf422127283c08e['h0322e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01918] =  Ifd35529b44c957737bf422127283c08e['h03230] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01919] =  Ifd35529b44c957737bf422127283c08e['h03232] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0191a] =  Ifd35529b44c957737bf422127283c08e['h03234] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0191b] =  Ifd35529b44c957737bf422127283c08e['h03236] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0191c] =  Ifd35529b44c957737bf422127283c08e['h03238] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0191d] =  Ifd35529b44c957737bf422127283c08e['h0323a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0191e] =  Ifd35529b44c957737bf422127283c08e['h0323c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0191f] =  Ifd35529b44c957737bf422127283c08e['h0323e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01920] =  Ifd35529b44c957737bf422127283c08e['h03240] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01921] =  Ifd35529b44c957737bf422127283c08e['h03242] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01922] =  Ifd35529b44c957737bf422127283c08e['h03244] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01923] =  Ifd35529b44c957737bf422127283c08e['h03246] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01924] =  Ifd35529b44c957737bf422127283c08e['h03248] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01925] =  Ifd35529b44c957737bf422127283c08e['h0324a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01926] =  Ifd35529b44c957737bf422127283c08e['h0324c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01927] =  Ifd35529b44c957737bf422127283c08e['h0324e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01928] =  Ifd35529b44c957737bf422127283c08e['h03250] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01929] =  Ifd35529b44c957737bf422127283c08e['h03252] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0192a] =  Ifd35529b44c957737bf422127283c08e['h03254] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0192b] =  Ifd35529b44c957737bf422127283c08e['h03256] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0192c] =  Ifd35529b44c957737bf422127283c08e['h03258] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0192d] =  Ifd35529b44c957737bf422127283c08e['h0325a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0192e] =  Ifd35529b44c957737bf422127283c08e['h0325c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0192f] =  Ifd35529b44c957737bf422127283c08e['h0325e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01930] =  Ifd35529b44c957737bf422127283c08e['h03260] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01931] =  Ifd35529b44c957737bf422127283c08e['h03262] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01932] =  Ifd35529b44c957737bf422127283c08e['h03264] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01933] =  Ifd35529b44c957737bf422127283c08e['h03266] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01934] =  Ifd35529b44c957737bf422127283c08e['h03268] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01935] =  Ifd35529b44c957737bf422127283c08e['h0326a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01936] =  Ifd35529b44c957737bf422127283c08e['h0326c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01937] =  Ifd35529b44c957737bf422127283c08e['h0326e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01938] =  Ifd35529b44c957737bf422127283c08e['h03270] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01939] =  Ifd35529b44c957737bf422127283c08e['h03272] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0193a] =  Ifd35529b44c957737bf422127283c08e['h03274] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0193b] =  Ifd35529b44c957737bf422127283c08e['h03276] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0193c] =  Ifd35529b44c957737bf422127283c08e['h03278] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0193d] =  Ifd35529b44c957737bf422127283c08e['h0327a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0193e] =  Ifd35529b44c957737bf422127283c08e['h0327c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0193f] =  Ifd35529b44c957737bf422127283c08e['h0327e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01940] =  Ifd35529b44c957737bf422127283c08e['h03280] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01941] =  Ifd35529b44c957737bf422127283c08e['h03282] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01942] =  Ifd35529b44c957737bf422127283c08e['h03284] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01943] =  Ifd35529b44c957737bf422127283c08e['h03286] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01944] =  Ifd35529b44c957737bf422127283c08e['h03288] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01945] =  Ifd35529b44c957737bf422127283c08e['h0328a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01946] =  Ifd35529b44c957737bf422127283c08e['h0328c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01947] =  Ifd35529b44c957737bf422127283c08e['h0328e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01948] =  Ifd35529b44c957737bf422127283c08e['h03290] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01949] =  Ifd35529b44c957737bf422127283c08e['h03292] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0194a] =  Ifd35529b44c957737bf422127283c08e['h03294] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0194b] =  Ifd35529b44c957737bf422127283c08e['h03296] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0194c] =  Ifd35529b44c957737bf422127283c08e['h03298] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0194d] =  Ifd35529b44c957737bf422127283c08e['h0329a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0194e] =  Ifd35529b44c957737bf422127283c08e['h0329c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0194f] =  Ifd35529b44c957737bf422127283c08e['h0329e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01950] =  Ifd35529b44c957737bf422127283c08e['h032a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01951] =  Ifd35529b44c957737bf422127283c08e['h032a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01952] =  Ifd35529b44c957737bf422127283c08e['h032a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01953] =  Ifd35529b44c957737bf422127283c08e['h032a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01954] =  Ifd35529b44c957737bf422127283c08e['h032a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01955] =  Ifd35529b44c957737bf422127283c08e['h032aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01956] =  Ifd35529b44c957737bf422127283c08e['h032ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01957] =  Ifd35529b44c957737bf422127283c08e['h032ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01958] =  Ifd35529b44c957737bf422127283c08e['h032b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01959] =  Ifd35529b44c957737bf422127283c08e['h032b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0195a] =  Ifd35529b44c957737bf422127283c08e['h032b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0195b] =  Ifd35529b44c957737bf422127283c08e['h032b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0195c] =  Ifd35529b44c957737bf422127283c08e['h032b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0195d] =  Ifd35529b44c957737bf422127283c08e['h032ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0195e] =  Ifd35529b44c957737bf422127283c08e['h032bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0195f] =  Ifd35529b44c957737bf422127283c08e['h032be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01960] =  Ifd35529b44c957737bf422127283c08e['h032c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01961] =  Ifd35529b44c957737bf422127283c08e['h032c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01962] =  Ifd35529b44c957737bf422127283c08e['h032c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01963] =  Ifd35529b44c957737bf422127283c08e['h032c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01964] =  Ifd35529b44c957737bf422127283c08e['h032c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01965] =  Ifd35529b44c957737bf422127283c08e['h032ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01966] =  Ifd35529b44c957737bf422127283c08e['h032cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01967] =  Ifd35529b44c957737bf422127283c08e['h032ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01968] =  Ifd35529b44c957737bf422127283c08e['h032d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01969] =  Ifd35529b44c957737bf422127283c08e['h032d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0196a] =  Ifd35529b44c957737bf422127283c08e['h032d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0196b] =  Ifd35529b44c957737bf422127283c08e['h032d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0196c] =  Ifd35529b44c957737bf422127283c08e['h032d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0196d] =  Ifd35529b44c957737bf422127283c08e['h032da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0196e] =  Ifd35529b44c957737bf422127283c08e['h032dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0196f] =  Ifd35529b44c957737bf422127283c08e['h032de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01970] =  Ifd35529b44c957737bf422127283c08e['h032e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01971] =  Ifd35529b44c957737bf422127283c08e['h032e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01972] =  Ifd35529b44c957737bf422127283c08e['h032e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01973] =  Ifd35529b44c957737bf422127283c08e['h032e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01974] =  Ifd35529b44c957737bf422127283c08e['h032e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01975] =  Ifd35529b44c957737bf422127283c08e['h032ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01976] =  Ifd35529b44c957737bf422127283c08e['h032ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01977] =  Ifd35529b44c957737bf422127283c08e['h032ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01978] =  Ifd35529b44c957737bf422127283c08e['h032f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01979] =  Ifd35529b44c957737bf422127283c08e['h032f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0197a] =  Ifd35529b44c957737bf422127283c08e['h032f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0197b] =  Ifd35529b44c957737bf422127283c08e['h032f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0197c] =  Ifd35529b44c957737bf422127283c08e['h032f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0197d] =  Ifd35529b44c957737bf422127283c08e['h032fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0197e] =  Ifd35529b44c957737bf422127283c08e['h032fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0197f] =  Ifd35529b44c957737bf422127283c08e['h032fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01980] =  Ifd35529b44c957737bf422127283c08e['h03300] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01981] =  Ifd35529b44c957737bf422127283c08e['h03302] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01982] =  Ifd35529b44c957737bf422127283c08e['h03304] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01983] =  Ifd35529b44c957737bf422127283c08e['h03306] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01984] =  Ifd35529b44c957737bf422127283c08e['h03308] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01985] =  Ifd35529b44c957737bf422127283c08e['h0330a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01986] =  Ifd35529b44c957737bf422127283c08e['h0330c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01987] =  Ifd35529b44c957737bf422127283c08e['h0330e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01988] =  Ifd35529b44c957737bf422127283c08e['h03310] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01989] =  Ifd35529b44c957737bf422127283c08e['h03312] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0198a] =  Ifd35529b44c957737bf422127283c08e['h03314] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0198b] =  Ifd35529b44c957737bf422127283c08e['h03316] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0198c] =  Ifd35529b44c957737bf422127283c08e['h03318] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0198d] =  Ifd35529b44c957737bf422127283c08e['h0331a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0198e] =  Ifd35529b44c957737bf422127283c08e['h0331c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0198f] =  Ifd35529b44c957737bf422127283c08e['h0331e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01990] =  Ifd35529b44c957737bf422127283c08e['h03320] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01991] =  Ifd35529b44c957737bf422127283c08e['h03322] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01992] =  Ifd35529b44c957737bf422127283c08e['h03324] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01993] =  Ifd35529b44c957737bf422127283c08e['h03326] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01994] =  Ifd35529b44c957737bf422127283c08e['h03328] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01995] =  Ifd35529b44c957737bf422127283c08e['h0332a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01996] =  Ifd35529b44c957737bf422127283c08e['h0332c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01997] =  Ifd35529b44c957737bf422127283c08e['h0332e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01998] =  Ifd35529b44c957737bf422127283c08e['h03330] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01999] =  Ifd35529b44c957737bf422127283c08e['h03332] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0199a] =  Ifd35529b44c957737bf422127283c08e['h03334] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0199b] =  Ifd35529b44c957737bf422127283c08e['h03336] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0199c] =  Ifd35529b44c957737bf422127283c08e['h03338] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0199d] =  Ifd35529b44c957737bf422127283c08e['h0333a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0199e] =  Ifd35529b44c957737bf422127283c08e['h0333c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h0199f] =  Ifd35529b44c957737bf422127283c08e['h0333e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019a0] =  Ifd35529b44c957737bf422127283c08e['h03340] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019a1] =  Ifd35529b44c957737bf422127283c08e['h03342] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019a2] =  Ifd35529b44c957737bf422127283c08e['h03344] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019a3] =  Ifd35529b44c957737bf422127283c08e['h03346] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019a4] =  Ifd35529b44c957737bf422127283c08e['h03348] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019a5] =  Ifd35529b44c957737bf422127283c08e['h0334a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019a6] =  Ifd35529b44c957737bf422127283c08e['h0334c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019a7] =  Ifd35529b44c957737bf422127283c08e['h0334e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019a8] =  Ifd35529b44c957737bf422127283c08e['h03350] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019a9] =  Ifd35529b44c957737bf422127283c08e['h03352] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019aa] =  Ifd35529b44c957737bf422127283c08e['h03354] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019ab] =  Ifd35529b44c957737bf422127283c08e['h03356] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019ac] =  Ifd35529b44c957737bf422127283c08e['h03358] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019ad] =  Ifd35529b44c957737bf422127283c08e['h0335a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019ae] =  Ifd35529b44c957737bf422127283c08e['h0335c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019af] =  Ifd35529b44c957737bf422127283c08e['h0335e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019b0] =  Ifd35529b44c957737bf422127283c08e['h03360] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019b1] =  Ifd35529b44c957737bf422127283c08e['h03362] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019b2] =  Ifd35529b44c957737bf422127283c08e['h03364] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019b3] =  Ifd35529b44c957737bf422127283c08e['h03366] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019b4] =  Ifd35529b44c957737bf422127283c08e['h03368] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019b5] =  Ifd35529b44c957737bf422127283c08e['h0336a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019b6] =  Ifd35529b44c957737bf422127283c08e['h0336c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019b7] =  Ifd35529b44c957737bf422127283c08e['h0336e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019b8] =  Ifd35529b44c957737bf422127283c08e['h03370] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019b9] =  Ifd35529b44c957737bf422127283c08e['h03372] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019ba] =  Ifd35529b44c957737bf422127283c08e['h03374] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019bb] =  Ifd35529b44c957737bf422127283c08e['h03376] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019bc] =  Ifd35529b44c957737bf422127283c08e['h03378] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019bd] =  Ifd35529b44c957737bf422127283c08e['h0337a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019be] =  Ifd35529b44c957737bf422127283c08e['h0337c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019bf] =  Ifd35529b44c957737bf422127283c08e['h0337e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019c0] =  Ifd35529b44c957737bf422127283c08e['h03380] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019c1] =  Ifd35529b44c957737bf422127283c08e['h03382] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019c2] =  Ifd35529b44c957737bf422127283c08e['h03384] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019c3] =  Ifd35529b44c957737bf422127283c08e['h03386] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019c4] =  Ifd35529b44c957737bf422127283c08e['h03388] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019c5] =  Ifd35529b44c957737bf422127283c08e['h0338a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019c6] =  Ifd35529b44c957737bf422127283c08e['h0338c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019c7] =  Ifd35529b44c957737bf422127283c08e['h0338e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019c8] =  Ifd35529b44c957737bf422127283c08e['h03390] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019c9] =  Ifd35529b44c957737bf422127283c08e['h03392] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019ca] =  Ifd35529b44c957737bf422127283c08e['h03394] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019cb] =  Ifd35529b44c957737bf422127283c08e['h03396] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019cc] =  Ifd35529b44c957737bf422127283c08e['h03398] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019cd] =  Ifd35529b44c957737bf422127283c08e['h0339a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019ce] =  Ifd35529b44c957737bf422127283c08e['h0339c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019cf] =  Ifd35529b44c957737bf422127283c08e['h0339e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019d0] =  Ifd35529b44c957737bf422127283c08e['h033a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019d1] =  Ifd35529b44c957737bf422127283c08e['h033a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019d2] =  Ifd35529b44c957737bf422127283c08e['h033a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019d3] =  Ifd35529b44c957737bf422127283c08e['h033a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019d4] =  Ifd35529b44c957737bf422127283c08e['h033a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019d5] =  Ifd35529b44c957737bf422127283c08e['h033aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019d6] =  Ifd35529b44c957737bf422127283c08e['h033ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019d7] =  Ifd35529b44c957737bf422127283c08e['h033ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019d8] =  Ifd35529b44c957737bf422127283c08e['h033b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019d9] =  Ifd35529b44c957737bf422127283c08e['h033b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019da] =  Ifd35529b44c957737bf422127283c08e['h033b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019db] =  Ifd35529b44c957737bf422127283c08e['h033b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019dc] =  Ifd35529b44c957737bf422127283c08e['h033b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019dd] =  Ifd35529b44c957737bf422127283c08e['h033ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019de] =  Ifd35529b44c957737bf422127283c08e['h033bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019df] =  Ifd35529b44c957737bf422127283c08e['h033be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019e0] =  Ifd35529b44c957737bf422127283c08e['h033c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019e1] =  Ifd35529b44c957737bf422127283c08e['h033c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019e2] =  Ifd35529b44c957737bf422127283c08e['h033c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019e3] =  Ifd35529b44c957737bf422127283c08e['h033c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019e4] =  Ifd35529b44c957737bf422127283c08e['h033c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019e5] =  Ifd35529b44c957737bf422127283c08e['h033ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019e6] =  Ifd35529b44c957737bf422127283c08e['h033cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019e7] =  Ifd35529b44c957737bf422127283c08e['h033ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019e8] =  Ifd35529b44c957737bf422127283c08e['h033d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019e9] =  Ifd35529b44c957737bf422127283c08e['h033d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019ea] =  Ifd35529b44c957737bf422127283c08e['h033d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019eb] =  Ifd35529b44c957737bf422127283c08e['h033d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019ec] =  Ifd35529b44c957737bf422127283c08e['h033d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019ed] =  Ifd35529b44c957737bf422127283c08e['h033da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019ee] =  Ifd35529b44c957737bf422127283c08e['h033dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019ef] =  Ifd35529b44c957737bf422127283c08e['h033de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019f0] =  Ifd35529b44c957737bf422127283c08e['h033e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019f1] =  Ifd35529b44c957737bf422127283c08e['h033e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019f2] =  Ifd35529b44c957737bf422127283c08e['h033e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019f3] =  Ifd35529b44c957737bf422127283c08e['h033e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019f4] =  Ifd35529b44c957737bf422127283c08e['h033e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019f5] =  Ifd35529b44c957737bf422127283c08e['h033ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019f6] =  Ifd35529b44c957737bf422127283c08e['h033ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019f7] =  Ifd35529b44c957737bf422127283c08e['h033ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019f8] =  Ifd35529b44c957737bf422127283c08e['h033f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019f9] =  Ifd35529b44c957737bf422127283c08e['h033f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019fa] =  Ifd35529b44c957737bf422127283c08e['h033f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019fb] =  Ifd35529b44c957737bf422127283c08e['h033f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019fc] =  Ifd35529b44c957737bf422127283c08e['h033f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019fd] =  Ifd35529b44c957737bf422127283c08e['h033fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019fe] =  Ifd35529b44c957737bf422127283c08e['h033fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h019ff] =  Ifd35529b44c957737bf422127283c08e['h033fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a00] =  Ifd35529b44c957737bf422127283c08e['h03400] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a01] =  Ifd35529b44c957737bf422127283c08e['h03402] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a02] =  Ifd35529b44c957737bf422127283c08e['h03404] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a03] =  Ifd35529b44c957737bf422127283c08e['h03406] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a04] =  Ifd35529b44c957737bf422127283c08e['h03408] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a05] =  Ifd35529b44c957737bf422127283c08e['h0340a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a06] =  Ifd35529b44c957737bf422127283c08e['h0340c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a07] =  Ifd35529b44c957737bf422127283c08e['h0340e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a08] =  Ifd35529b44c957737bf422127283c08e['h03410] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a09] =  Ifd35529b44c957737bf422127283c08e['h03412] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a0a] =  Ifd35529b44c957737bf422127283c08e['h03414] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a0b] =  Ifd35529b44c957737bf422127283c08e['h03416] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a0c] =  Ifd35529b44c957737bf422127283c08e['h03418] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a0d] =  Ifd35529b44c957737bf422127283c08e['h0341a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a0e] =  Ifd35529b44c957737bf422127283c08e['h0341c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a0f] =  Ifd35529b44c957737bf422127283c08e['h0341e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a10] =  Ifd35529b44c957737bf422127283c08e['h03420] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a11] =  Ifd35529b44c957737bf422127283c08e['h03422] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a12] =  Ifd35529b44c957737bf422127283c08e['h03424] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a13] =  Ifd35529b44c957737bf422127283c08e['h03426] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a14] =  Ifd35529b44c957737bf422127283c08e['h03428] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a15] =  Ifd35529b44c957737bf422127283c08e['h0342a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a16] =  Ifd35529b44c957737bf422127283c08e['h0342c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a17] =  Ifd35529b44c957737bf422127283c08e['h0342e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a18] =  Ifd35529b44c957737bf422127283c08e['h03430] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a19] =  Ifd35529b44c957737bf422127283c08e['h03432] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a1a] =  Ifd35529b44c957737bf422127283c08e['h03434] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a1b] =  Ifd35529b44c957737bf422127283c08e['h03436] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a1c] =  Ifd35529b44c957737bf422127283c08e['h03438] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a1d] =  Ifd35529b44c957737bf422127283c08e['h0343a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a1e] =  Ifd35529b44c957737bf422127283c08e['h0343c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a1f] =  Ifd35529b44c957737bf422127283c08e['h0343e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a20] =  Ifd35529b44c957737bf422127283c08e['h03440] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a21] =  Ifd35529b44c957737bf422127283c08e['h03442] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a22] =  Ifd35529b44c957737bf422127283c08e['h03444] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a23] =  Ifd35529b44c957737bf422127283c08e['h03446] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a24] =  Ifd35529b44c957737bf422127283c08e['h03448] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a25] =  Ifd35529b44c957737bf422127283c08e['h0344a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a26] =  Ifd35529b44c957737bf422127283c08e['h0344c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a27] =  Ifd35529b44c957737bf422127283c08e['h0344e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a28] =  Ifd35529b44c957737bf422127283c08e['h03450] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a29] =  Ifd35529b44c957737bf422127283c08e['h03452] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a2a] =  Ifd35529b44c957737bf422127283c08e['h03454] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a2b] =  Ifd35529b44c957737bf422127283c08e['h03456] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a2c] =  Ifd35529b44c957737bf422127283c08e['h03458] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a2d] =  Ifd35529b44c957737bf422127283c08e['h0345a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a2e] =  Ifd35529b44c957737bf422127283c08e['h0345c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a2f] =  Ifd35529b44c957737bf422127283c08e['h0345e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a30] =  Ifd35529b44c957737bf422127283c08e['h03460] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a31] =  Ifd35529b44c957737bf422127283c08e['h03462] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a32] =  Ifd35529b44c957737bf422127283c08e['h03464] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a33] =  Ifd35529b44c957737bf422127283c08e['h03466] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a34] =  Ifd35529b44c957737bf422127283c08e['h03468] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a35] =  Ifd35529b44c957737bf422127283c08e['h0346a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a36] =  Ifd35529b44c957737bf422127283c08e['h0346c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a37] =  Ifd35529b44c957737bf422127283c08e['h0346e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a38] =  Ifd35529b44c957737bf422127283c08e['h03470] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a39] =  Ifd35529b44c957737bf422127283c08e['h03472] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a3a] =  Ifd35529b44c957737bf422127283c08e['h03474] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a3b] =  Ifd35529b44c957737bf422127283c08e['h03476] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a3c] =  Ifd35529b44c957737bf422127283c08e['h03478] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a3d] =  Ifd35529b44c957737bf422127283c08e['h0347a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a3e] =  Ifd35529b44c957737bf422127283c08e['h0347c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a3f] =  Ifd35529b44c957737bf422127283c08e['h0347e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a40] =  Ifd35529b44c957737bf422127283c08e['h03480] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a41] =  Ifd35529b44c957737bf422127283c08e['h03482] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a42] =  Ifd35529b44c957737bf422127283c08e['h03484] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a43] =  Ifd35529b44c957737bf422127283c08e['h03486] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a44] =  Ifd35529b44c957737bf422127283c08e['h03488] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a45] =  Ifd35529b44c957737bf422127283c08e['h0348a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a46] =  Ifd35529b44c957737bf422127283c08e['h0348c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a47] =  Ifd35529b44c957737bf422127283c08e['h0348e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a48] =  Ifd35529b44c957737bf422127283c08e['h03490] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a49] =  Ifd35529b44c957737bf422127283c08e['h03492] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a4a] =  Ifd35529b44c957737bf422127283c08e['h03494] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a4b] =  Ifd35529b44c957737bf422127283c08e['h03496] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a4c] =  Ifd35529b44c957737bf422127283c08e['h03498] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a4d] =  Ifd35529b44c957737bf422127283c08e['h0349a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a4e] =  Ifd35529b44c957737bf422127283c08e['h0349c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a4f] =  Ifd35529b44c957737bf422127283c08e['h0349e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a50] =  Ifd35529b44c957737bf422127283c08e['h034a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a51] =  Ifd35529b44c957737bf422127283c08e['h034a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a52] =  Ifd35529b44c957737bf422127283c08e['h034a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a53] =  Ifd35529b44c957737bf422127283c08e['h034a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a54] =  Ifd35529b44c957737bf422127283c08e['h034a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a55] =  Ifd35529b44c957737bf422127283c08e['h034aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a56] =  Ifd35529b44c957737bf422127283c08e['h034ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a57] =  Ifd35529b44c957737bf422127283c08e['h034ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a58] =  Ifd35529b44c957737bf422127283c08e['h034b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a59] =  Ifd35529b44c957737bf422127283c08e['h034b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a5a] =  Ifd35529b44c957737bf422127283c08e['h034b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a5b] =  Ifd35529b44c957737bf422127283c08e['h034b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a5c] =  Ifd35529b44c957737bf422127283c08e['h034b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a5d] =  Ifd35529b44c957737bf422127283c08e['h034ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a5e] =  Ifd35529b44c957737bf422127283c08e['h034bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a5f] =  Ifd35529b44c957737bf422127283c08e['h034be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a60] =  Ifd35529b44c957737bf422127283c08e['h034c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a61] =  Ifd35529b44c957737bf422127283c08e['h034c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a62] =  Ifd35529b44c957737bf422127283c08e['h034c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a63] =  Ifd35529b44c957737bf422127283c08e['h034c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a64] =  Ifd35529b44c957737bf422127283c08e['h034c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a65] =  Ifd35529b44c957737bf422127283c08e['h034ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a66] =  Ifd35529b44c957737bf422127283c08e['h034cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a67] =  Ifd35529b44c957737bf422127283c08e['h034ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a68] =  Ifd35529b44c957737bf422127283c08e['h034d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a69] =  Ifd35529b44c957737bf422127283c08e['h034d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a6a] =  Ifd35529b44c957737bf422127283c08e['h034d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a6b] =  Ifd35529b44c957737bf422127283c08e['h034d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a6c] =  Ifd35529b44c957737bf422127283c08e['h034d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a6d] =  Ifd35529b44c957737bf422127283c08e['h034da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a6e] =  Ifd35529b44c957737bf422127283c08e['h034dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a6f] =  Ifd35529b44c957737bf422127283c08e['h034de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a70] =  Ifd35529b44c957737bf422127283c08e['h034e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a71] =  Ifd35529b44c957737bf422127283c08e['h034e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a72] =  Ifd35529b44c957737bf422127283c08e['h034e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a73] =  Ifd35529b44c957737bf422127283c08e['h034e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a74] =  Ifd35529b44c957737bf422127283c08e['h034e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a75] =  Ifd35529b44c957737bf422127283c08e['h034ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a76] =  Ifd35529b44c957737bf422127283c08e['h034ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a77] =  Ifd35529b44c957737bf422127283c08e['h034ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a78] =  Ifd35529b44c957737bf422127283c08e['h034f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a79] =  Ifd35529b44c957737bf422127283c08e['h034f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a7a] =  Ifd35529b44c957737bf422127283c08e['h034f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a7b] =  Ifd35529b44c957737bf422127283c08e['h034f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a7c] =  Ifd35529b44c957737bf422127283c08e['h034f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a7d] =  Ifd35529b44c957737bf422127283c08e['h034fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a7e] =  Ifd35529b44c957737bf422127283c08e['h034fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a7f] =  Ifd35529b44c957737bf422127283c08e['h034fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a80] =  Ifd35529b44c957737bf422127283c08e['h03500] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a81] =  Ifd35529b44c957737bf422127283c08e['h03502] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a82] =  Ifd35529b44c957737bf422127283c08e['h03504] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a83] =  Ifd35529b44c957737bf422127283c08e['h03506] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a84] =  Ifd35529b44c957737bf422127283c08e['h03508] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a85] =  Ifd35529b44c957737bf422127283c08e['h0350a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a86] =  Ifd35529b44c957737bf422127283c08e['h0350c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a87] =  Ifd35529b44c957737bf422127283c08e['h0350e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a88] =  Ifd35529b44c957737bf422127283c08e['h03510] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a89] =  Ifd35529b44c957737bf422127283c08e['h03512] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a8a] =  Ifd35529b44c957737bf422127283c08e['h03514] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a8b] =  Ifd35529b44c957737bf422127283c08e['h03516] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a8c] =  Ifd35529b44c957737bf422127283c08e['h03518] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a8d] =  Ifd35529b44c957737bf422127283c08e['h0351a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a8e] =  Ifd35529b44c957737bf422127283c08e['h0351c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a8f] =  Ifd35529b44c957737bf422127283c08e['h0351e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a90] =  Ifd35529b44c957737bf422127283c08e['h03520] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a91] =  Ifd35529b44c957737bf422127283c08e['h03522] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a92] =  Ifd35529b44c957737bf422127283c08e['h03524] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a93] =  Ifd35529b44c957737bf422127283c08e['h03526] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a94] =  Ifd35529b44c957737bf422127283c08e['h03528] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a95] =  Ifd35529b44c957737bf422127283c08e['h0352a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a96] =  Ifd35529b44c957737bf422127283c08e['h0352c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a97] =  Ifd35529b44c957737bf422127283c08e['h0352e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a98] =  Ifd35529b44c957737bf422127283c08e['h03530] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a99] =  Ifd35529b44c957737bf422127283c08e['h03532] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a9a] =  Ifd35529b44c957737bf422127283c08e['h03534] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a9b] =  Ifd35529b44c957737bf422127283c08e['h03536] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a9c] =  Ifd35529b44c957737bf422127283c08e['h03538] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a9d] =  Ifd35529b44c957737bf422127283c08e['h0353a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a9e] =  Ifd35529b44c957737bf422127283c08e['h0353c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01a9f] =  Ifd35529b44c957737bf422127283c08e['h0353e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01aa0] =  Ifd35529b44c957737bf422127283c08e['h03540] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01aa1] =  Ifd35529b44c957737bf422127283c08e['h03542] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01aa2] =  Ifd35529b44c957737bf422127283c08e['h03544] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01aa3] =  Ifd35529b44c957737bf422127283c08e['h03546] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01aa4] =  Ifd35529b44c957737bf422127283c08e['h03548] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01aa5] =  Ifd35529b44c957737bf422127283c08e['h0354a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01aa6] =  Ifd35529b44c957737bf422127283c08e['h0354c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01aa7] =  Ifd35529b44c957737bf422127283c08e['h0354e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01aa8] =  Ifd35529b44c957737bf422127283c08e['h03550] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01aa9] =  Ifd35529b44c957737bf422127283c08e['h03552] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01aaa] =  Ifd35529b44c957737bf422127283c08e['h03554] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01aab] =  Ifd35529b44c957737bf422127283c08e['h03556] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01aac] =  Ifd35529b44c957737bf422127283c08e['h03558] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01aad] =  Ifd35529b44c957737bf422127283c08e['h0355a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01aae] =  Ifd35529b44c957737bf422127283c08e['h0355c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01aaf] =  Ifd35529b44c957737bf422127283c08e['h0355e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ab0] =  Ifd35529b44c957737bf422127283c08e['h03560] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ab1] =  Ifd35529b44c957737bf422127283c08e['h03562] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ab2] =  Ifd35529b44c957737bf422127283c08e['h03564] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ab3] =  Ifd35529b44c957737bf422127283c08e['h03566] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ab4] =  Ifd35529b44c957737bf422127283c08e['h03568] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ab5] =  Ifd35529b44c957737bf422127283c08e['h0356a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ab6] =  Ifd35529b44c957737bf422127283c08e['h0356c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ab7] =  Ifd35529b44c957737bf422127283c08e['h0356e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ab8] =  Ifd35529b44c957737bf422127283c08e['h03570] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ab9] =  Ifd35529b44c957737bf422127283c08e['h03572] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01aba] =  Ifd35529b44c957737bf422127283c08e['h03574] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01abb] =  Ifd35529b44c957737bf422127283c08e['h03576] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01abc] =  Ifd35529b44c957737bf422127283c08e['h03578] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01abd] =  Ifd35529b44c957737bf422127283c08e['h0357a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01abe] =  Ifd35529b44c957737bf422127283c08e['h0357c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01abf] =  Ifd35529b44c957737bf422127283c08e['h0357e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ac0] =  Ifd35529b44c957737bf422127283c08e['h03580] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ac1] =  Ifd35529b44c957737bf422127283c08e['h03582] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ac2] =  Ifd35529b44c957737bf422127283c08e['h03584] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ac3] =  Ifd35529b44c957737bf422127283c08e['h03586] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ac4] =  Ifd35529b44c957737bf422127283c08e['h03588] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ac5] =  Ifd35529b44c957737bf422127283c08e['h0358a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ac6] =  Ifd35529b44c957737bf422127283c08e['h0358c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ac7] =  Ifd35529b44c957737bf422127283c08e['h0358e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ac8] =  Ifd35529b44c957737bf422127283c08e['h03590] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ac9] =  Ifd35529b44c957737bf422127283c08e['h03592] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01aca] =  Ifd35529b44c957737bf422127283c08e['h03594] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01acb] =  Ifd35529b44c957737bf422127283c08e['h03596] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01acc] =  Ifd35529b44c957737bf422127283c08e['h03598] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01acd] =  Ifd35529b44c957737bf422127283c08e['h0359a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ace] =  Ifd35529b44c957737bf422127283c08e['h0359c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01acf] =  Ifd35529b44c957737bf422127283c08e['h0359e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ad0] =  Ifd35529b44c957737bf422127283c08e['h035a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ad1] =  Ifd35529b44c957737bf422127283c08e['h035a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ad2] =  Ifd35529b44c957737bf422127283c08e['h035a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ad3] =  Ifd35529b44c957737bf422127283c08e['h035a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ad4] =  Ifd35529b44c957737bf422127283c08e['h035a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ad5] =  Ifd35529b44c957737bf422127283c08e['h035aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ad6] =  Ifd35529b44c957737bf422127283c08e['h035ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ad7] =  Ifd35529b44c957737bf422127283c08e['h035ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ad8] =  Ifd35529b44c957737bf422127283c08e['h035b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ad9] =  Ifd35529b44c957737bf422127283c08e['h035b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ada] =  Ifd35529b44c957737bf422127283c08e['h035b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01adb] =  Ifd35529b44c957737bf422127283c08e['h035b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01adc] =  Ifd35529b44c957737bf422127283c08e['h035b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01add] =  Ifd35529b44c957737bf422127283c08e['h035ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ade] =  Ifd35529b44c957737bf422127283c08e['h035bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01adf] =  Ifd35529b44c957737bf422127283c08e['h035be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ae0] =  Ifd35529b44c957737bf422127283c08e['h035c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ae1] =  Ifd35529b44c957737bf422127283c08e['h035c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ae2] =  Ifd35529b44c957737bf422127283c08e['h035c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ae3] =  Ifd35529b44c957737bf422127283c08e['h035c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ae4] =  Ifd35529b44c957737bf422127283c08e['h035c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ae5] =  Ifd35529b44c957737bf422127283c08e['h035ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ae6] =  Ifd35529b44c957737bf422127283c08e['h035cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ae7] =  Ifd35529b44c957737bf422127283c08e['h035ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ae8] =  Ifd35529b44c957737bf422127283c08e['h035d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ae9] =  Ifd35529b44c957737bf422127283c08e['h035d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01aea] =  Ifd35529b44c957737bf422127283c08e['h035d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01aeb] =  Ifd35529b44c957737bf422127283c08e['h035d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01aec] =  Ifd35529b44c957737bf422127283c08e['h035d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01aed] =  Ifd35529b44c957737bf422127283c08e['h035da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01aee] =  Ifd35529b44c957737bf422127283c08e['h035dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01aef] =  Ifd35529b44c957737bf422127283c08e['h035de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01af0] =  Ifd35529b44c957737bf422127283c08e['h035e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01af1] =  Ifd35529b44c957737bf422127283c08e['h035e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01af2] =  Ifd35529b44c957737bf422127283c08e['h035e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01af3] =  Ifd35529b44c957737bf422127283c08e['h035e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01af4] =  Ifd35529b44c957737bf422127283c08e['h035e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01af5] =  Ifd35529b44c957737bf422127283c08e['h035ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01af6] =  Ifd35529b44c957737bf422127283c08e['h035ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01af7] =  Ifd35529b44c957737bf422127283c08e['h035ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01af8] =  Ifd35529b44c957737bf422127283c08e['h035f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01af9] =  Ifd35529b44c957737bf422127283c08e['h035f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01afa] =  Ifd35529b44c957737bf422127283c08e['h035f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01afb] =  Ifd35529b44c957737bf422127283c08e['h035f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01afc] =  Ifd35529b44c957737bf422127283c08e['h035f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01afd] =  Ifd35529b44c957737bf422127283c08e['h035fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01afe] =  Ifd35529b44c957737bf422127283c08e['h035fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01aff] =  Ifd35529b44c957737bf422127283c08e['h035fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b00] =  Ifd35529b44c957737bf422127283c08e['h03600] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b01] =  Ifd35529b44c957737bf422127283c08e['h03602] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b02] =  Ifd35529b44c957737bf422127283c08e['h03604] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b03] =  Ifd35529b44c957737bf422127283c08e['h03606] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b04] =  Ifd35529b44c957737bf422127283c08e['h03608] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b05] =  Ifd35529b44c957737bf422127283c08e['h0360a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b06] =  Ifd35529b44c957737bf422127283c08e['h0360c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b07] =  Ifd35529b44c957737bf422127283c08e['h0360e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b08] =  Ifd35529b44c957737bf422127283c08e['h03610] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b09] =  Ifd35529b44c957737bf422127283c08e['h03612] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b0a] =  Ifd35529b44c957737bf422127283c08e['h03614] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b0b] =  Ifd35529b44c957737bf422127283c08e['h03616] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b0c] =  Ifd35529b44c957737bf422127283c08e['h03618] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b0d] =  Ifd35529b44c957737bf422127283c08e['h0361a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b0e] =  Ifd35529b44c957737bf422127283c08e['h0361c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b0f] =  Ifd35529b44c957737bf422127283c08e['h0361e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b10] =  Ifd35529b44c957737bf422127283c08e['h03620] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b11] =  Ifd35529b44c957737bf422127283c08e['h03622] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b12] =  Ifd35529b44c957737bf422127283c08e['h03624] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b13] =  Ifd35529b44c957737bf422127283c08e['h03626] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b14] =  Ifd35529b44c957737bf422127283c08e['h03628] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b15] =  Ifd35529b44c957737bf422127283c08e['h0362a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b16] =  Ifd35529b44c957737bf422127283c08e['h0362c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b17] =  Ifd35529b44c957737bf422127283c08e['h0362e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b18] =  Ifd35529b44c957737bf422127283c08e['h03630] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b19] =  Ifd35529b44c957737bf422127283c08e['h03632] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b1a] =  Ifd35529b44c957737bf422127283c08e['h03634] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b1b] =  Ifd35529b44c957737bf422127283c08e['h03636] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b1c] =  Ifd35529b44c957737bf422127283c08e['h03638] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b1d] =  Ifd35529b44c957737bf422127283c08e['h0363a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b1e] =  Ifd35529b44c957737bf422127283c08e['h0363c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b1f] =  Ifd35529b44c957737bf422127283c08e['h0363e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b20] =  Ifd35529b44c957737bf422127283c08e['h03640] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b21] =  Ifd35529b44c957737bf422127283c08e['h03642] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b22] =  Ifd35529b44c957737bf422127283c08e['h03644] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b23] =  Ifd35529b44c957737bf422127283c08e['h03646] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b24] =  Ifd35529b44c957737bf422127283c08e['h03648] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b25] =  Ifd35529b44c957737bf422127283c08e['h0364a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b26] =  Ifd35529b44c957737bf422127283c08e['h0364c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b27] =  Ifd35529b44c957737bf422127283c08e['h0364e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b28] =  Ifd35529b44c957737bf422127283c08e['h03650] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b29] =  Ifd35529b44c957737bf422127283c08e['h03652] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b2a] =  Ifd35529b44c957737bf422127283c08e['h03654] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b2b] =  Ifd35529b44c957737bf422127283c08e['h03656] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b2c] =  Ifd35529b44c957737bf422127283c08e['h03658] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b2d] =  Ifd35529b44c957737bf422127283c08e['h0365a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b2e] =  Ifd35529b44c957737bf422127283c08e['h0365c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b2f] =  Ifd35529b44c957737bf422127283c08e['h0365e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b30] =  Ifd35529b44c957737bf422127283c08e['h03660] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b31] =  Ifd35529b44c957737bf422127283c08e['h03662] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b32] =  Ifd35529b44c957737bf422127283c08e['h03664] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b33] =  Ifd35529b44c957737bf422127283c08e['h03666] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b34] =  Ifd35529b44c957737bf422127283c08e['h03668] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b35] =  Ifd35529b44c957737bf422127283c08e['h0366a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b36] =  Ifd35529b44c957737bf422127283c08e['h0366c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b37] =  Ifd35529b44c957737bf422127283c08e['h0366e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b38] =  Ifd35529b44c957737bf422127283c08e['h03670] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b39] =  Ifd35529b44c957737bf422127283c08e['h03672] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b3a] =  Ifd35529b44c957737bf422127283c08e['h03674] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b3b] =  Ifd35529b44c957737bf422127283c08e['h03676] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b3c] =  Ifd35529b44c957737bf422127283c08e['h03678] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b3d] =  Ifd35529b44c957737bf422127283c08e['h0367a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b3e] =  Ifd35529b44c957737bf422127283c08e['h0367c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b3f] =  Ifd35529b44c957737bf422127283c08e['h0367e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b40] =  Ifd35529b44c957737bf422127283c08e['h03680] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b41] =  Ifd35529b44c957737bf422127283c08e['h03682] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b42] =  Ifd35529b44c957737bf422127283c08e['h03684] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b43] =  Ifd35529b44c957737bf422127283c08e['h03686] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b44] =  Ifd35529b44c957737bf422127283c08e['h03688] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b45] =  Ifd35529b44c957737bf422127283c08e['h0368a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b46] =  Ifd35529b44c957737bf422127283c08e['h0368c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b47] =  Ifd35529b44c957737bf422127283c08e['h0368e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b48] =  Ifd35529b44c957737bf422127283c08e['h03690] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b49] =  Ifd35529b44c957737bf422127283c08e['h03692] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b4a] =  Ifd35529b44c957737bf422127283c08e['h03694] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b4b] =  Ifd35529b44c957737bf422127283c08e['h03696] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b4c] =  Ifd35529b44c957737bf422127283c08e['h03698] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b4d] =  Ifd35529b44c957737bf422127283c08e['h0369a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b4e] =  Ifd35529b44c957737bf422127283c08e['h0369c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b4f] =  Ifd35529b44c957737bf422127283c08e['h0369e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b50] =  Ifd35529b44c957737bf422127283c08e['h036a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b51] =  Ifd35529b44c957737bf422127283c08e['h036a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b52] =  Ifd35529b44c957737bf422127283c08e['h036a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b53] =  Ifd35529b44c957737bf422127283c08e['h036a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b54] =  Ifd35529b44c957737bf422127283c08e['h036a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b55] =  Ifd35529b44c957737bf422127283c08e['h036aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b56] =  Ifd35529b44c957737bf422127283c08e['h036ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b57] =  Ifd35529b44c957737bf422127283c08e['h036ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b58] =  Ifd35529b44c957737bf422127283c08e['h036b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b59] =  Ifd35529b44c957737bf422127283c08e['h036b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b5a] =  Ifd35529b44c957737bf422127283c08e['h036b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b5b] =  Ifd35529b44c957737bf422127283c08e['h036b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b5c] =  Ifd35529b44c957737bf422127283c08e['h036b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b5d] =  Ifd35529b44c957737bf422127283c08e['h036ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b5e] =  Ifd35529b44c957737bf422127283c08e['h036bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b5f] =  Ifd35529b44c957737bf422127283c08e['h036be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b60] =  Ifd35529b44c957737bf422127283c08e['h036c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b61] =  Ifd35529b44c957737bf422127283c08e['h036c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b62] =  Ifd35529b44c957737bf422127283c08e['h036c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b63] =  Ifd35529b44c957737bf422127283c08e['h036c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b64] =  Ifd35529b44c957737bf422127283c08e['h036c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b65] =  Ifd35529b44c957737bf422127283c08e['h036ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b66] =  Ifd35529b44c957737bf422127283c08e['h036cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b67] =  Ifd35529b44c957737bf422127283c08e['h036ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b68] =  Ifd35529b44c957737bf422127283c08e['h036d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b69] =  Ifd35529b44c957737bf422127283c08e['h036d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b6a] =  Ifd35529b44c957737bf422127283c08e['h036d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b6b] =  Ifd35529b44c957737bf422127283c08e['h036d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b6c] =  Ifd35529b44c957737bf422127283c08e['h036d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b6d] =  Ifd35529b44c957737bf422127283c08e['h036da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b6e] =  Ifd35529b44c957737bf422127283c08e['h036dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b6f] =  Ifd35529b44c957737bf422127283c08e['h036de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b70] =  Ifd35529b44c957737bf422127283c08e['h036e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b71] =  Ifd35529b44c957737bf422127283c08e['h036e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b72] =  Ifd35529b44c957737bf422127283c08e['h036e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b73] =  Ifd35529b44c957737bf422127283c08e['h036e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b74] =  Ifd35529b44c957737bf422127283c08e['h036e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b75] =  Ifd35529b44c957737bf422127283c08e['h036ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b76] =  Ifd35529b44c957737bf422127283c08e['h036ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b77] =  Ifd35529b44c957737bf422127283c08e['h036ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b78] =  Ifd35529b44c957737bf422127283c08e['h036f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b79] =  Ifd35529b44c957737bf422127283c08e['h036f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b7a] =  Ifd35529b44c957737bf422127283c08e['h036f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b7b] =  Ifd35529b44c957737bf422127283c08e['h036f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b7c] =  Ifd35529b44c957737bf422127283c08e['h036f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b7d] =  Ifd35529b44c957737bf422127283c08e['h036fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b7e] =  Ifd35529b44c957737bf422127283c08e['h036fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b7f] =  Ifd35529b44c957737bf422127283c08e['h036fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b80] =  Ifd35529b44c957737bf422127283c08e['h03700] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b81] =  Ifd35529b44c957737bf422127283c08e['h03702] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b82] =  Ifd35529b44c957737bf422127283c08e['h03704] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b83] =  Ifd35529b44c957737bf422127283c08e['h03706] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b84] =  Ifd35529b44c957737bf422127283c08e['h03708] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b85] =  Ifd35529b44c957737bf422127283c08e['h0370a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b86] =  Ifd35529b44c957737bf422127283c08e['h0370c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b87] =  Ifd35529b44c957737bf422127283c08e['h0370e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b88] =  Ifd35529b44c957737bf422127283c08e['h03710] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b89] =  Ifd35529b44c957737bf422127283c08e['h03712] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b8a] =  Ifd35529b44c957737bf422127283c08e['h03714] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b8b] =  Ifd35529b44c957737bf422127283c08e['h03716] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b8c] =  Ifd35529b44c957737bf422127283c08e['h03718] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b8d] =  Ifd35529b44c957737bf422127283c08e['h0371a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b8e] =  Ifd35529b44c957737bf422127283c08e['h0371c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b8f] =  Ifd35529b44c957737bf422127283c08e['h0371e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b90] =  Ifd35529b44c957737bf422127283c08e['h03720] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b91] =  Ifd35529b44c957737bf422127283c08e['h03722] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b92] =  Ifd35529b44c957737bf422127283c08e['h03724] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b93] =  Ifd35529b44c957737bf422127283c08e['h03726] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b94] =  Ifd35529b44c957737bf422127283c08e['h03728] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b95] =  Ifd35529b44c957737bf422127283c08e['h0372a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b96] =  Ifd35529b44c957737bf422127283c08e['h0372c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b97] =  Ifd35529b44c957737bf422127283c08e['h0372e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b98] =  Ifd35529b44c957737bf422127283c08e['h03730] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b99] =  Ifd35529b44c957737bf422127283c08e['h03732] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b9a] =  Ifd35529b44c957737bf422127283c08e['h03734] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b9b] =  Ifd35529b44c957737bf422127283c08e['h03736] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b9c] =  Ifd35529b44c957737bf422127283c08e['h03738] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b9d] =  Ifd35529b44c957737bf422127283c08e['h0373a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b9e] =  Ifd35529b44c957737bf422127283c08e['h0373c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01b9f] =  Ifd35529b44c957737bf422127283c08e['h0373e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ba0] =  Ifd35529b44c957737bf422127283c08e['h03740] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ba1] =  Ifd35529b44c957737bf422127283c08e['h03742] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ba2] =  Ifd35529b44c957737bf422127283c08e['h03744] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ba3] =  Ifd35529b44c957737bf422127283c08e['h03746] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ba4] =  Ifd35529b44c957737bf422127283c08e['h03748] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ba5] =  Ifd35529b44c957737bf422127283c08e['h0374a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ba6] =  Ifd35529b44c957737bf422127283c08e['h0374c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ba7] =  Ifd35529b44c957737bf422127283c08e['h0374e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ba8] =  Ifd35529b44c957737bf422127283c08e['h03750] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ba9] =  Ifd35529b44c957737bf422127283c08e['h03752] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01baa] =  Ifd35529b44c957737bf422127283c08e['h03754] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bab] =  Ifd35529b44c957737bf422127283c08e['h03756] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bac] =  Ifd35529b44c957737bf422127283c08e['h03758] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bad] =  Ifd35529b44c957737bf422127283c08e['h0375a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bae] =  Ifd35529b44c957737bf422127283c08e['h0375c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01baf] =  Ifd35529b44c957737bf422127283c08e['h0375e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bb0] =  Ifd35529b44c957737bf422127283c08e['h03760] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bb1] =  Ifd35529b44c957737bf422127283c08e['h03762] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bb2] =  Ifd35529b44c957737bf422127283c08e['h03764] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bb3] =  Ifd35529b44c957737bf422127283c08e['h03766] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bb4] =  Ifd35529b44c957737bf422127283c08e['h03768] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bb5] =  Ifd35529b44c957737bf422127283c08e['h0376a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bb6] =  Ifd35529b44c957737bf422127283c08e['h0376c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bb7] =  Ifd35529b44c957737bf422127283c08e['h0376e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bb8] =  Ifd35529b44c957737bf422127283c08e['h03770] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bb9] =  Ifd35529b44c957737bf422127283c08e['h03772] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bba] =  Ifd35529b44c957737bf422127283c08e['h03774] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bbb] =  Ifd35529b44c957737bf422127283c08e['h03776] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bbc] =  Ifd35529b44c957737bf422127283c08e['h03778] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bbd] =  Ifd35529b44c957737bf422127283c08e['h0377a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bbe] =  Ifd35529b44c957737bf422127283c08e['h0377c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bbf] =  Ifd35529b44c957737bf422127283c08e['h0377e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bc0] =  Ifd35529b44c957737bf422127283c08e['h03780] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bc1] =  Ifd35529b44c957737bf422127283c08e['h03782] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bc2] =  Ifd35529b44c957737bf422127283c08e['h03784] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bc3] =  Ifd35529b44c957737bf422127283c08e['h03786] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bc4] =  Ifd35529b44c957737bf422127283c08e['h03788] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bc5] =  Ifd35529b44c957737bf422127283c08e['h0378a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bc6] =  Ifd35529b44c957737bf422127283c08e['h0378c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bc7] =  Ifd35529b44c957737bf422127283c08e['h0378e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bc8] =  Ifd35529b44c957737bf422127283c08e['h03790] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bc9] =  Ifd35529b44c957737bf422127283c08e['h03792] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bca] =  Ifd35529b44c957737bf422127283c08e['h03794] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bcb] =  Ifd35529b44c957737bf422127283c08e['h03796] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bcc] =  Ifd35529b44c957737bf422127283c08e['h03798] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bcd] =  Ifd35529b44c957737bf422127283c08e['h0379a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bce] =  Ifd35529b44c957737bf422127283c08e['h0379c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bcf] =  Ifd35529b44c957737bf422127283c08e['h0379e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bd0] =  Ifd35529b44c957737bf422127283c08e['h037a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bd1] =  Ifd35529b44c957737bf422127283c08e['h037a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bd2] =  Ifd35529b44c957737bf422127283c08e['h037a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bd3] =  Ifd35529b44c957737bf422127283c08e['h037a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bd4] =  Ifd35529b44c957737bf422127283c08e['h037a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bd5] =  Ifd35529b44c957737bf422127283c08e['h037aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bd6] =  Ifd35529b44c957737bf422127283c08e['h037ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bd7] =  Ifd35529b44c957737bf422127283c08e['h037ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bd8] =  Ifd35529b44c957737bf422127283c08e['h037b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bd9] =  Ifd35529b44c957737bf422127283c08e['h037b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bda] =  Ifd35529b44c957737bf422127283c08e['h037b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bdb] =  Ifd35529b44c957737bf422127283c08e['h037b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bdc] =  Ifd35529b44c957737bf422127283c08e['h037b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bdd] =  Ifd35529b44c957737bf422127283c08e['h037ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bde] =  Ifd35529b44c957737bf422127283c08e['h037bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bdf] =  Ifd35529b44c957737bf422127283c08e['h037be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01be0] =  Ifd35529b44c957737bf422127283c08e['h037c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01be1] =  Ifd35529b44c957737bf422127283c08e['h037c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01be2] =  Ifd35529b44c957737bf422127283c08e['h037c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01be3] =  Ifd35529b44c957737bf422127283c08e['h037c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01be4] =  Ifd35529b44c957737bf422127283c08e['h037c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01be5] =  Ifd35529b44c957737bf422127283c08e['h037ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01be6] =  Ifd35529b44c957737bf422127283c08e['h037cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01be7] =  Ifd35529b44c957737bf422127283c08e['h037ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01be8] =  Ifd35529b44c957737bf422127283c08e['h037d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01be9] =  Ifd35529b44c957737bf422127283c08e['h037d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bea] =  Ifd35529b44c957737bf422127283c08e['h037d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01beb] =  Ifd35529b44c957737bf422127283c08e['h037d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bec] =  Ifd35529b44c957737bf422127283c08e['h037d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bed] =  Ifd35529b44c957737bf422127283c08e['h037da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bee] =  Ifd35529b44c957737bf422127283c08e['h037dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bef] =  Ifd35529b44c957737bf422127283c08e['h037de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bf0] =  Ifd35529b44c957737bf422127283c08e['h037e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bf1] =  Ifd35529b44c957737bf422127283c08e['h037e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bf2] =  Ifd35529b44c957737bf422127283c08e['h037e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bf3] =  Ifd35529b44c957737bf422127283c08e['h037e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bf4] =  Ifd35529b44c957737bf422127283c08e['h037e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bf5] =  Ifd35529b44c957737bf422127283c08e['h037ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bf6] =  Ifd35529b44c957737bf422127283c08e['h037ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bf7] =  Ifd35529b44c957737bf422127283c08e['h037ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bf8] =  Ifd35529b44c957737bf422127283c08e['h037f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bf9] =  Ifd35529b44c957737bf422127283c08e['h037f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bfa] =  Ifd35529b44c957737bf422127283c08e['h037f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bfb] =  Ifd35529b44c957737bf422127283c08e['h037f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bfc] =  Ifd35529b44c957737bf422127283c08e['h037f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bfd] =  Ifd35529b44c957737bf422127283c08e['h037fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bfe] =  Ifd35529b44c957737bf422127283c08e['h037fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01bff] =  Ifd35529b44c957737bf422127283c08e['h037fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c00] =  Ifd35529b44c957737bf422127283c08e['h03800] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c01] =  Ifd35529b44c957737bf422127283c08e['h03802] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c02] =  Ifd35529b44c957737bf422127283c08e['h03804] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c03] =  Ifd35529b44c957737bf422127283c08e['h03806] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c04] =  Ifd35529b44c957737bf422127283c08e['h03808] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c05] =  Ifd35529b44c957737bf422127283c08e['h0380a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c06] =  Ifd35529b44c957737bf422127283c08e['h0380c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c07] =  Ifd35529b44c957737bf422127283c08e['h0380e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c08] =  Ifd35529b44c957737bf422127283c08e['h03810] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c09] =  Ifd35529b44c957737bf422127283c08e['h03812] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c0a] =  Ifd35529b44c957737bf422127283c08e['h03814] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c0b] =  Ifd35529b44c957737bf422127283c08e['h03816] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c0c] =  Ifd35529b44c957737bf422127283c08e['h03818] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c0d] =  Ifd35529b44c957737bf422127283c08e['h0381a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c0e] =  Ifd35529b44c957737bf422127283c08e['h0381c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c0f] =  Ifd35529b44c957737bf422127283c08e['h0381e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c10] =  Ifd35529b44c957737bf422127283c08e['h03820] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c11] =  Ifd35529b44c957737bf422127283c08e['h03822] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c12] =  Ifd35529b44c957737bf422127283c08e['h03824] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c13] =  Ifd35529b44c957737bf422127283c08e['h03826] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c14] =  Ifd35529b44c957737bf422127283c08e['h03828] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c15] =  Ifd35529b44c957737bf422127283c08e['h0382a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c16] =  Ifd35529b44c957737bf422127283c08e['h0382c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c17] =  Ifd35529b44c957737bf422127283c08e['h0382e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c18] =  Ifd35529b44c957737bf422127283c08e['h03830] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c19] =  Ifd35529b44c957737bf422127283c08e['h03832] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c1a] =  Ifd35529b44c957737bf422127283c08e['h03834] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c1b] =  Ifd35529b44c957737bf422127283c08e['h03836] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c1c] =  Ifd35529b44c957737bf422127283c08e['h03838] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c1d] =  Ifd35529b44c957737bf422127283c08e['h0383a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c1e] =  Ifd35529b44c957737bf422127283c08e['h0383c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c1f] =  Ifd35529b44c957737bf422127283c08e['h0383e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c20] =  Ifd35529b44c957737bf422127283c08e['h03840] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c21] =  Ifd35529b44c957737bf422127283c08e['h03842] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c22] =  Ifd35529b44c957737bf422127283c08e['h03844] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c23] =  Ifd35529b44c957737bf422127283c08e['h03846] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c24] =  Ifd35529b44c957737bf422127283c08e['h03848] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c25] =  Ifd35529b44c957737bf422127283c08e['h0384a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c26] =  Ifd35529b44c957737bf422127283c08e['h0384c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c27] =  Ifd35529b44c957737bf422127283c08e['h0384e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c28] =  Ifd35529b44c957737bf422127283c08e['h03850] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c29] =  Ifd35529b44c957737bf422127283c08e['h03852] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c2a] =  Ifd35529b44c957737bf422127283c08e['h03854] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c2b] =  Ifd35529b44c957737bf422127283c08e['h03856] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c2c] =  Ifd35529b44c957737bf422127283c08e['h03858] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c2d] =  Ifd35529b44c957737bf422127283c08e['h0385a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c2e] =  Ifd35529b44c957737bf422127283c08e['h0385c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c2f] =  Ifd35529b44c957737bf422127283c08e['h0385e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c30] =  Ifd35529b44c957737bf422127283c08e['h03860] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c31] =  Ifd35529b44c957737bf422127283c08e['h03862] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c32] =  Ifd35529b44c957737bf422127283c08e['h03864] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c33] =  Ifd35529b44c957737bf422127283c08e['h03866] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c34] =  Ifd35529b44c957737bf422127283c08e['h03868] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c35] =  Ifd35529b44c957737bf422127283c08e['h0386a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c36] =  Ifd35529b44c957737bf422127283c08e['h0386c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c37] =  Ifd35529b44c957737bf422127283c08e['h0386e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c38] =  Ifd35529b44c957737bf422127283c08e['h03870] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c39] =  Ifd35529b44c957737bf422127283c08e['h03872] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c3a] =  Ifd35529b44c957737bf422127283c08e['h03874] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c3b] =  Ifd35529b44c957737bf422127283c08e['h03876] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c3c] =  Ifd35529b44c957737bf422127283c08e['h03878] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c3d] =  Ifd35529b44c957737bf422127283c08e['h0387a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c3e] =  Ifd35529b44c957737bf422127283c08e['h0387c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c3f] =  Ifd35529b44c957737bf422127283c08e['h0387e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c40] =  Ifd35529b44c957737bf422127283c08e['h03880] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c41] =  Ifd35529b44c957737bf422127283c08e['h03882] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c42] =  Ifd35529b44c957737bf422127283c08e['h03884] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c43] =  Ifd35529b44c957737bf422127283c08e['h03886] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c44] =  Ifd35529b44c957737bf422127283c08e['h03888] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c45] =  Ifd35529b44c957737bf422127283c08e['h0388a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c46] =  Ifd35529b44c957737bf422127283c08e['h0388c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c47] =  Ifd35529b44c957737bf422127283c08e['h0388e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c48] =  Ifd35529b44c957737bf422127283c08e['h03890] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c49] =  Ifd35529b44c957737bf422127283c08e['h03892] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c4a] =  Ifd35529b44c957737bf422127283c08e['h03894] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c4b] =  Ifd35529b44c957737bf422127283c08e['h03896] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c4c] =  Ifd35529b44c957737bf422127283c08e['h03898] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c4d] =  Ifd35529b44c957737bf422127283c08e['h0389a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c4e] =  Ifd35529b44c957737bf422127283c08e['h0389c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c4f] =  Ifd35529b44c957737bf422127283c08e['h0389e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c50] =  Ifd35529b44c957737bf422127283c08e['h038a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c51] =  Ifd35529b44c957737bf422127283c08e['h038a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c52] =  Ifd35529b44c957737bf422127283c08e['h038a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c53] =  Ifd35529b44c957737bf422127283c08e['h038a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c54] =  Ifd35529b44c957737bf422127283c08e['h038a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c55] =  Ifd35529b44c957737bf422127283c08e['h038aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c56] =  Ifd35529b44c957737bf422127283c08e['h038ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c57] =  Ifd35529b44c957737bf422127283c08e['h038ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c58] =  Ifd35529b44c957737bf422127283c08e['h038b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c59] =  Ifd35529b44c957737bf422127283c08e['h038b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c5a] =  Ifd35529b44c957737bf422127283c08e['h038b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c5b] =  Ifd35529b44c957737bf422127283c08e['h038b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c5c] =  Ifd35529b44c957737bf422127283c08e['h038b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c5d] =  Ifd35529b44c957737bf422127283c08e['h038ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c5e] =  Ifd35529b44c957737bf422127283c08e['h038bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c5f] =  Ifd35529b44c957737bf422127283c08e['h038be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c60] =  Ifd35529b44c957737bf422127283c08e['h038c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c61] =  Ifd35529b44c957737bf422127283c08e['h038c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c62] =  Ifd35529b44c957737bf422127283c08e['h038c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c63] =  Ifd35529b44c957737bf422127283c08e['h038c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c64] =  Ifd35529b44c957737bf422127283c08e['h038c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c65] =  Ifd35529b44c957737bf422127283c08e['h038ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c66] =  Ifd35529b44c957737bf422127283c08e['h038cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c67] =  Ifd35529b44c957737bf422127283c08e['h038ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c68] =  Ifd35529b44c957737bf422127283c08e['h038d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c69] =  Ifd35529b44c957737bf422127283c08e['h038d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c6a] =  Ifd35529b44c957737bf422127283c08e['h038d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c6b] =  Ifd35529b44c957737bf422127283c08e['h038d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c6c] =  Ifd35529b44c957737bf422127283c08e['h038d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c6d] =  Ifd35529b44c957737bf422127283c08e['h038da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c6e] =  Ifd35529b44c957737bf422127283c08e['h038dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c6f] =  Ifd35529b44c957737bf422127283c08e['h038de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c70] =  Ifd35529b44c957737bf422127283c08e['h038e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c71] =  Ifd35529b44c957737bf422127283c08e['h038e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c72] =  Ifd35529b44c957737bf422127283c08e['h038e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c73] =  Ifd35529b44c957737bf422127283c08e['h038e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c74] =  Ifd35529b44c957737bf422127283c08e['h038e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c75] =  Ifd35529b44c957737bf422127283c08e['h038ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c76] =  Ifd35529b44c957737bf422127283c08e['h038ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c77] =  Ifd35529b44c957737bf422127283c08e['h038ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c78] =  Ifd35529b44c957737bf422127283c08e['h038f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c79] =  Ifd35529b44c957737bf422127283c08e['h038f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c7a] =  Ifd35529b44c957737bf422127283c08e['h038f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c7b] =  Ifd35529b44c957737bf422127283c08e['h038f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c7c] =  Ifd35529b44c957737bf422127283c08e['h038f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c7d] =  Ifd35529b44c957737bf422127283c08e['h038fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c7e] =  Ifd35529b44c957737bf422127283c08e['h038fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c7f] =  Ifd35529b44c957737bf422127283c08e['h038fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c80] =  Ifd35529b44c957737bf422127283c08e['h03900] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c81] =  Ifd35529b44c957737bf422127283c08e['h03902] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c82] =  Ifd35529b44c957737bf422127283c08e['h03904] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c83] =  Ifd35529b44c957737bf422127283c08e['h03906] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c84] =  Ifd35529b44c957737bf422127283c08e['h03908] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c85] =  Ifd35529b44c957737bf422127283c08e['h0390a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c86] =  Ifd35529b44c957737bf422127283c08e['h0390c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c87] =  Ifd35529b44c957737bf422127283c08e['h0390e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c88] =  Ifd35529b44c957737bf422127283c08e['h03910] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c89] =  Ifd35529b44c957737bf422127283c08e['h03912] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c8a] =  Ifd35529b44c957737bf422127283c08e['h03914] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c8b] =  Ifd35529b44c957737bf422127283c08e['h03916] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c8c] =  Ifd35529b44c957737bf422127283c08e['h03918] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c8d] =  Ifd35529b44c957737bf422127283c08e['h0391a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c8e] =  Ifd35529b44c957737bf422127283c08e['h0391c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c8f] =  Ifd35529b44c957737bf422127283c08e['h0391e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c90] =  Ifd35529b44c957737bf422127283c08e['h03920] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c91] =  Ifd35529b44c957737bf422127283c08e['h03922] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c92] =  Ifd35529b44c957737bf422127283c08e['h03924] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c93] =  Ifd35529b44c957737bf422127283c08e['h03926] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c94] =  Ifd35529b44c957737bf422127283c08e['h03928] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c95] =  Ifd35529b44c957737bf422127283c08e['h0392a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c96] =  Ifd35529b44c957737bf422127283c08e['h0392c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c97] =  Ifd35529b44c957737bf422127283c08e['h0392e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c98] =  Ifd35529b44c957737bf422127283c08e['h03930] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c99] =  Ifd35529b44c957737bf422127283c08e['h03932] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c9a] =  Ifd35529b44c957737bf422127283c08e['h03934] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c9b] =  Ifd35529b44c957737bf422127283c08e['h03936] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c9c] =  Ifd35529b44c957737bf422127283c08e['h03938] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c9d] =  Ifd35529b44c957737bf422127283c08e['h0393a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c9e] =  Ifd35529b44c957737bf422127283c08e['h0393c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01c9f] =  Ifd35529b44c957737bf422127283c08e['h0393e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ca0] =  Ifd35529b44c957737bf422127283c08e['h03940] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ca1] =  Ifd35529b44c957737bf422127283c08e['h03942] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ca2] =  Ifd35529b44c957737bf422127283c08e['h03944] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ca3] =  Ifd35529b44c957737bf422127283c08e['h03946] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ca4] =  Ifd35529b44c957737bf422127283c08e['h03948] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ca5] =  Ifd35529b44c957737bf422127283c08e['h0394a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ca6] =  Ifd35529b44c957737bf422127283c08e['h0394c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ca7] =  Ifd35529b44c957737bf422127283c08e['h0394e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ca8] =  Ifd35529b44c957737bf422127283c08e['h03950] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ca9] =  Ifd35529b44c957737bf422127283c08e['h03952] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01caa] =  Ifd35529b44c957737bf422127283c08e['h03954] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cab] =  Ifd35529b44c957737bf422127283c08e['h03956] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cac] =  Ifd35529b44c957737bf422127283c08e['h03958] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cad] =  Ifd35529b44c957737bf422127283c08e['h0395a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cae] =  Ifd35529b44c957737bf422127283c08e['h0395c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01caf] =  Ifd35529b44c957737bf422127283c08e['h0395e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cb0] =  Ifd35529b44c957737bf422127283c08e['h03960] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cb1] =  Ifd35529b44c957737bf422127283c08e['h03962] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cb2] =  Ifd35529b44c957737bf422127283c08e['h03964] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cb3] =  Ifd35529b44c957737bf422127283c08e['h03966] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cb4] =  Ifd35529b44c957737bf422127283c08e['h03968] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cb5] =  Ifd35529b44c957737bf422127283c08e['h0396a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cb6] =  Ifd35529b44c957737bf422127283c08e['h0396c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cb7] =  Ifd35529b44c957737bf422127283c08e['h0396e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cb8] =  Ifd35529b44c957737bf422127283c08e['h03970] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cb9] =  Ifd35529b44c957737bf422127283c08e['h03972] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cba] =  Ifd35529b44c957737bf422127283c08e['h03974] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cbb] =  Ifd35529b44c957737bf422127283c08e['h03976] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cbc] =  Ifd35529b44c957737bf422127283c08e['h03978] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cbd] =  Ifd35529b44c957737bf422127283c08e['h0397a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cbe] =  Ifd35529b44c957737bf422127283c08e['h0397c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cbf] =  Ifd35529b44c957737bf422127283c08e['h0397e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cc0] =  Ifd35529b44c957737bf422127283c08e['h03980] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cc1] =  Ifd35529b44c957737bf422127283c08e['h03982] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cc2] =  Ifd35529b44c957737bf422127283c08e['h03984] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cc3] =  Ifd35529b44c957737bf422127283c08e['h03986] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cc4] =  Ifd35529b44c957737bf422127283c08e['h03988] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cc5] =  Ifd35529b44c957737bf422127283c08e['h0398a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cc6] =  Ifd35529b44c957737bf422127283c08e['h0398c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cc7] =  Ifd35529b44c957737bf422127283c08e['h0398e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cc8] =  Ifd35529b44c957737bf422127283c08e['h03990] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cc9] =  Ifd35529b44c957737bf422127283c08e['h03992] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cca] =  Ifd35529b44c957737bf422127283c08e['h03994] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ccb] =  Ifd35529b44c957737bf422127283c08e['h03996] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ccc] =  Ifd35529b44c957737bf422127283c08e['h03998] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ccd] =  Ifd35529b44c957737bf422127283c08e['h0399a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cce] =  Ifd35529b44c957737bf422127283c08e['h0399c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ccf] =  Ifd35529b44c957737bf422127283c08e['h0399e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cd0] =  Ifd35529b44c957737bf422127283c08e['h039a0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cd1] =  Ifd35529b44c957737bf422127283c08e['h039a2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cd2] =  Ifd35529b44c957737bf422127283c08e['h039a4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cd3] =  Ifd35529b44c957737bf422127283c08e['h039a6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cd4] =  Ifd35529b44c957737bf422127283c08e['h039a8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cd5] =  Ifd35529b44c957737bf422127283c08e['h039aa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cd6] =  Ifd35529b44c957737bf422127283c08e['h039ac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cd7] =  Ifd35529b44c957737bf422127283c08e['h039ae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cd8] =  Ifd35529b44c957737bf422127283c08e['h039b0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cd9] =  Ifd35529b44c957737bf422127283c08e['h039b2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cda] =  Ifd35529b44c957737bf422127283c08e['h039b4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cdb] =  Ifd35529b44c957737bf422127283c08e['h039b6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cdc] =  Ifd35529b44c957737bf422127283c08e['h039b8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cdd] =  Ifd35529b44c957737bf422127283c08e['h039ba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cde] =  Ifd35529b44c957737bf422127283c08e['h039bc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cdf] =  Ifd35529b44c957737bf422127283c08e['h039be] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ce0] =  Ifd35529b44c957737bf422127283c08e['h039c0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ce1] =  Ifd35529b44c957737bf422127283c08e['h039c2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ce2] =  Ifd35529b44c957737bf422127283c08e['h039c4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ce3] =  Ifd35529b44c957737bf422127283c08e['h039c6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ce4] =  Ifd35529b44c957737bf422127283c08e['h039c8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ce5] =  Ifd35529b44c957737bf422127283c08e['h039ca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ce6] =  Ifd35529b44c957737bf422127283c08e['h039cc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ce7] =  Ifd35529b44c957737bf422127283c08e['h039ce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ce8] =  Ifd35529b44c957737bf422127283c08e['h039d0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ce9] =  Ifd35529b44c957737bf422127283c08e['h039d2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cea] =  Ifd35529b44c957737bf422127283c08e['h039d4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ceb] =  Ifd35529b44c957737bf422127283c08e['h039d6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cec] =  Ifd35529b44c957737bf422127283c08e['h039d8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ced] =  Ifd35529b44c957737bf422127283c08e['h039da] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cee] =  Ifd35529b44c957737bf422127283c08e['h039dc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cef] =  Ifd35529b44c957737bf422127283c08e['h039de] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cf0] =  Ifd35529b44c957737bf422127283c08e['h039e0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cf1] =  Ifd35529b44c957737bf422127283c08e['h039e2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cf2] =  Ifd35529b44c957737bf422127283c08e['h039e4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cf3] =  Ifd35529b44c957737bf422127283c08e['h039e6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cf4] =  Ifd35529b44c957737bf422127283c08e['h039e8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cf5] =  Ifd35529b44c957737bf422127283c08e['h039ea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cf6] =  Ifd35529b44c957737bf422127283c08e['h039ec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cf7] =  Ifd35529b44c957737bf422127283c08e['h039ee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cf8] =  Ifd35529b44c957737bf422127283c08e['h039f0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cf9] =  Ifd35529b44c957737bf422127283c08e['h039f2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cfa] =  Ifd35529b44c957737bf422127283c08e['h039f4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cfb] =  Ifd35529b44c957737bf422127283c08e['h039f6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cfc] =  Ifd35529b44c957737bf422127283c08e['h039f8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cfd] =  Ifd35529b44c957737bf422127283c08e['h039fa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cfe] =  Ifd35529b44c957737bf422127283c08e['h039fc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01cff] =  Ifd35529b44c957737bf422127283c08e['h039fe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d00] =  Ifd35529b44c957737bf422127283c08e['h03a00] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d01] =  Ifd35529b44c957737bf422127283c08e['h03a02] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d02] =  Ifd35529b44c957737bf422127283c08e['h03a04] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d03] =  Ifd35529b44c957737bf422127283c08e['h03a06] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d04] =  Ifd35529b44c957737bf422127283c08e['h03a08] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d05] =  Ifd35529b44c957737bf422127283c08e['h03a0a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d06] =  Ifd35529b44c957737bf422127283c08e['h03a0c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d07] =  Ifd35529b44c957737bf422127283c08e['h03a0e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d08] =  Ifd35529b44c957737bf422127283c08e['h03a10] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d09] =  Ifd35529b44c957737bf422127283c08e['h03a12] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d0a] =  Ifd35529b44c957737bf422127283c08e['h03a14] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d0b] =  Ifd35529b44c957737bf422127283c08e['h03a16] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d0c] =  Ifd35529b44c957737bf422127283c08e['h03a18] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d0d] =  Ifd35529b44c957737bf422127283c08e['h03a1a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d0e] =  Ifd35529b44c957737bf422127283c08e['h03a1c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d0f] =  Ifd35529b44c957737bf422127283c08e['h03a1e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d10] =  Ifd35529b44c957737bf422127283c08e['h03a20] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d11] =  Ifd35529b44c957737bf422127283c08e['h03a22] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d12] =  Ifd35529b44c957737bf422127283c08e['h03a24] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d13] =  Ifd35529b44c957737bf422127283c08e['h03a26] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d14] =  Ifd35529b44c957737bf422127283c08e['h03a28] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d15] =  Ifd35529b44c957737bf422127283c08e['h03a2a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d16] =  Ifd35529b44c957737bf422127283c08e['h03a2c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d17] =  Ifd35529b44c957737bf422127283c08e['h03a2e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d18] =  Ifd35529b44c957737bf422127283c08e['h03a30] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d19] =  Ifd35529b44c957737bf422127283c08e['h03a32] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d1a] =  Ifd35529b44c957737bf422127283c08e['h03a34] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d1b] =  Ifd35529b44c957737bf422127283c08e['h03a36] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d1c] =  Ifd35529b44c957737bf422127283c08e['h03a38] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d1d] =  Ifd35529b44c957737bf422127283c08e['h03a3a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d1e] =  Ifd35529b44c957737bf422127283c08e['h03a3c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d1f] =  Ifd35529b44c957737bf422127283c08e['h03a3e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d20] =  Ifd35529b44c957737bf422127283c08e['h03a40] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d21] =  Ifd35529b44c957737bf422127283c08e['h03a42] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d22] =  Ifd35529b44c957737bf422127283c08e['h03a44] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d23] =  Ifd35529b44c957737bf422127283c08e['h03a46] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d24] =  Ifd35529b44c957737bf422127283c08e['h03a48] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d25] =  Ifd35529b44c957737bf422127283c08e['h03a4a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d26] =  Ifd35529b44c957737bf422127283c08e['h03a4c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d27] =  Ifd35529b44c957737bf422127283c08e['h03a4e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d28] =  Ifd35529b44c957737bf422127283c08e['h03a50] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d29] =  Ifd35529b44c957737bf422127283c08e['h03a52] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d2a] =  Ifd35529b44c957737bf422127283c08e['h03a54] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d2b] =  Ifd35529b44c957737bf422127283c08e['h03a56] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d2c] =  Ifd35529b44c957737bf422127283c08e['h03a58] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d2d] =  Ifd35529b44c957737bf422127283c08e['h03a5a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d2e] =  Ifd35529b44c957737bf422127283c08e['h03a5c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d2f] =  Ifd35529b44c957737bf422127283c08e['h03a5e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d30] =  Ifd35529b44c957737bf422127283c08e['h03a60] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d31] =  Ifd35529b44c957737bf422127283c08e['h03a62] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d32] =  Ifd35529b44c957737bf422127283c08e['h03a64] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d33] =  Ifd35529b44c957737bf422127283c08e['h03a66] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d34] =  Ifd35529b44c957737bf422127283c08e['h03a68] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d35] =  Ifd35529b44c957737bf422127283c08e['h03a6a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d36] =  Ifd35529b44c957737bf422127283c08e['h03a6c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d37] =  Ifd35529b44c957737bf422127283c08e['h03a6e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d38] =  Ifd35529b44c957737bf422127283c08e['h03a70] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d39] =  Ifd35529b44c957737bf422127283c08e['h03a72] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d3a] =  Ifd35529b44c957737bf422127283c08e['h03a74] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d3b] =  Ifd35529b44c957737bf422127283c08e['h03a76] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d3c] =  Ifd35529b44c957737bf422127283c08e['h03a78] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d3d] =  Ifd35529b44c957737bf422127283c08e['h03a7a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d3e] =  Ifd35529b44c957737bf422127283c08e['h03a7c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d3f] =  Ifd35529b44c957737bf422127283c08e['h03a7e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d40] =  Ifd35529b44c957737bf422127283c08e['h03a80] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d41] =  Ifd35529b44c957737bf422127283c08e['h03a82] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d42] =  Ifd35529b44c957737bf422127283c08e['h03a84] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d43] =  Ifd35529b44c957737bf422127283c08e['h03a86] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d44] =  Ifd35529b44c957737bf422127283c08e['h03a88] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d45] =  Ifd35529b44c957737bf422127283c08e['h03a8a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d46] =  Ifd35529b44c957737bf422127283c08e['h03a8c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d47] =  Ifd35529b44c957737bf422127283c08e['h03a8e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d48] =  Ifd35529b44c957737bf422127283c08e['h03a90] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d49] =  Ifd35529b44c957737bf422127283c08e['h03a92] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d4a] =  Ifd35529b44c957737bf422127283c08e['h03a94] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d4b] =  Ifd35529b44c957737bf422127283c08e['h03a96] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d4c] =  Ifd35529b44c957737bf422127283c08e['h03a98] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d4d] =  Ifd35529b44c957737bf422127283c08e['h03a9a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d4e] =  Ifd35529b44c957737bf422127283c08e['h03a9c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d4f] =  Ifd35529b44c957737bf422127283c08e['h03a9e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d50] =  Ifd35529b44c957737bf422127283c08e['h03aa0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d51] =  Ifd35529b44c957737bf422127283c08e['h03aa2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d52] =  Ifd35529b44c957737bf422127283c08e['h03aa4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d53] =  Ifd35529b44c957737bf422127283c08e['h03aa6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d54] =  Ifd35529b44c957737bf422127283c08e['h03aa8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d55] =  Ifd35529b44c957737bf422127283c08e['h03aaa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d56] =  Ifd35529b44c957737bf422127283c08e['h03aac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d57] =  Ifd35529b44c957737bf422127283c08e['h03aae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d58] =  Ifd35529b44c957737bf422127283c08e['h03ab0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d59] =  Ifd35529b44c957737bf422127283c08e['h03ab2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d5a] =  Ifd35529b44c957737bf422127283c08e['h03ab4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d5b] =  Ifd35529b44c957737bf422127283c08e['h03ab6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d5c] =  Ifd35529b44c957737bf422127283c08e['h03ab8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d5d] =  Ifd35529b44c957737bf422127283c08e['h03aba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d5e] =  Ifd35529b44c957737bf422127283c08e['h03abc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d5f] =  Ifd35529b44c957737bf422127283c08e['h03abe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d60] =  Ifd35529b44c957737bf422127283c08e['h03ac0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d61] =  Ifd35529b44c957737bf422127283c08e['h03ac2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d62] =  Ifd35529b44c957737bf422127283c08e['h03ac4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d63] =  Ifd35529b44c957737bf422127283c08e['h03ac6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d64] =  Ifd35529b44c957737bf422127283c08e['h03ac8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d65] =  Ifd35529b44c957737bf422127283c08e['h03aca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d66] =  Ifd35529b44c957737bf422127283c08e['h03acc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d67] =  Ifd35529b44c957737bf422127283c08e['h03ace] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d68] =  Ifd35529b44c957737bf422127283c08e['h03ad0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d69] =  Ifd35529b44c957737bf422127283c08e['h03ad2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d6a] =  Ifd35529b44c957737bf422127283c08e['h03ad4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d6b] =  Ifd35529b44c957737bf422127283c08e['h03ad6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d6c] =  Ifd35529b44c957737bf422127283c08e['h03ad8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d6d] =  Ifd35529b44c957737bf422127283c08e['h03ada] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d6e] =  Ifd35529b44c957737bf422127283c08e['h03adc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d6f] =  Ifd35529b44c957737bf422127283c08e['h03ade] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d70] =  Ifd35529b44c957737bf422127283c08e['h03ae0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d71] =  Ifd35529b44c957737bf422127283c08e['h03ae2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d72] =  Ifd35529b44c957737bf422127283c08e['h03ae4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d73] =  Ifd35529b44c957737bf422127283c08e['h03ae6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d74] =  Ifd35529b44c957737bf422127283c08e['h03ae8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d75] =  Ifd35529b44c957737bf422127283c08e['h03aea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d76] =  Ifd35529b44c957737bf422127283c08e['h03aec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d77] =  Ifd35529b44c957737bf422127283c08e['h03aee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d78] =  Ifd35529b44c957737bf422127283c08e['h03af0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d79] =  Ifd35529b44c957737bf422127283c08e['h03af2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d7a] =  Ifd35529b44c957737bf422127283c08e['h03af4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d7b] =  Ifd35529b44c957737bf422127283c08e['h03af6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d7c] =  Ifd35529b44c957737bf422127283c08e['h03af8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d7d] =  Ifd35529b44c957737bf422127283c08e['h03afa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d7e] =  Ifd35529b44c957737bf422127283c08e['h03afc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d7f] =  Ifd35529b44c957737bf422127283c08e['h03afe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d80] =  Ifd35529b44c957737bf422127283c08e['h03b00] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d81] =  Ifd35529b44c957737bf422127283c08e['h03b02] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d82] =  Ifd35529b44c957737bf422127283c08e['h03b04] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d83] =  Ifd35529b44c957737bf422127283c08e['h03b06] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d84] =  Ifd35529b44c957737bf422127283c08e['h03b08] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d85] =  Ifd35529b44c957737bf422127283c08e['h03b0a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d86] =  Ifd35529b44c957737bf422127283c08e['h03b0c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d87] =  Ifd35529b44c957737bf422127283c08e['h03b0e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d88] =  Ifd35529b44c957737bf422127283c08e['h03b10] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d89] =  Ifd35529b44c957737bf422127283c08e['h03b12] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d8a] =  Ifd35529b44c957737bf422127283c08e['h03b14] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d8b] =  Ifd35529b44c957737bf422127283c08e['h03b16] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d8c] =  Ifd35529b44c957737bf422127283c08e['h03b18] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d8d] =  Ifd35529b44c957737bf422127283c08e['h03b1a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d8e] =  Ifd35529b44c957737bf422127283c08e['h03b1c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d8f] =  Ifd35529b44c957737bf422127283c08e['h03b1e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d90] =  Ifd35529b44c957737bf422127283c08e['h03b20] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d91] =  Ifd35529b44c957737bf422127283c08e['h03b22] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d92] =  Ifd35529b44c957737bf422127283c08e['h03b24] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d93] =  Ifd35529b44c957737bf422127283c08e['h03b26] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d94] =  Ifd35529b44c957737bf422127283c08e['h03b28] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d95] =  Ifd35529b44c957737bf422127283c08e['h03b2a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d96] =  Ifd35529b44c957737bf422127283c08e['h03b2c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d97] =  Ifd35529b44c957737bf422127283c08e['h03b2e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d98] =  Ifd35529b44c957737bf422127283c08e['h03b30] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d99] =  Ifd35529b44c957737bf422127283c08e['h03b32] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d9a] =  Ifd35529b44c957737bf422127283c08e['h03b34] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d9b] =  Ifd35529b44c957737bf422127283c08e['h03b36] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d9c] =  Ifd35529b44c957737bf422127283c08e['h03b38] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d9d] =  Ifd35529b44c957737bf422127283c08e['h03b3a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d9e] =  Ifd35529b44c957737bf422127283c08e['h03b3c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01d9f] =  Ifd35529b44c957737bf422127283c08e['h03b3e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01da0] =  Ifd35529b44c957737bf422127283c08e['h03b40] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01da1] =  Ifd35529b44c957737bf422127283c08e['h03b42] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01da2] =  Ifd35529b44c957737bf422127283c08e['h03b44] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01da3] =  Ifd35529b44c957737bf422127283c08e['h03b46] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01da4] =  Ifd35529b44c957737bf422127283c08e['h03b48] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01da5] =  Ifd35529b44c957737bf422127283c08e['h03b4a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01da6] =  Ifd35529b44c957737bf422127283c08e['h03b4c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01da7] =  Ifd35529b44c957737bf422127283c08e['h03b4e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01da8] =  Ifd35529b44c957737bf422127283c08e['h03b50] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01da9] =  Ifd35529b44c957737bf422127283c08e['h03b52] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01daa] =  Ifd35529b44c957737bf422127283c08e['h03b54] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dab] =  Ifd35529b44c957737bf422127283c08e['h03b56] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dac] =  Ifd35529b44c957737bf422127283c08e['h03b58] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dad] =  Ifd35529b44c957737bf422127283c08e['h03b5a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dae] =  Ifd35529b44c957737bf422127283c08e['h03b5c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01daf] =  Ifd35529b44c957737bf422127283c08e['h03b5e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01db0] =  Ifd35529b44c957737bf422127283c08e['h03b60] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01db1] =  Ifd35529b44c957737bf422127283c08e['h03b62] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01db2] =  Ifd35529b44c957737bf422127283c08e['h03b64] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01db3] =  Ifd35529b44c957737bf422127283c08e['h03b66] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01db4] =  Ifd35529b44c957737bf422127283c08e['h03b68] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01db5] =  Ifd35529b44c957737bf422127283c08e['h03b6a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01db6] =  Ifd35529b44c957737bf422127283c08e['h03b6c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01db7] =  Ifd35529b44c957737bf422127283c08e['h03b6e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01db8] =  Ifd35529b44c957737bf422127283c08e['h03b70] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01db9] =  Ifd35529b44c957737bf422127283c08e['h03b72] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dba] =  Ifd35529b44c957737bf422127283c08e['h03b74] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dbb] =  Ifd35529b44c957737bf422127283c08e['h03b76] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dbc] =  Ifd35529b44c957737bf422127283c08e['h03b78] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dbd] =  Ifd35529b44c957737bf422127283c08e['h03b7a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dbe] =  Ifd35529b44c957737bf422127283c08e['h03b7c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dbf] =  Ifd35529b44c957737bf422127283c08e['h03b7e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dc0] =  Ifd35529b44c957737bf422127283c08e['h03b80] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dc1] =  Ifd35529b44c957737bf422127283c08e['h03b82] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dc2] =  Ifd35529b44c957737bf422127283c08e['h03b84] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dc3] =  Ifd35529b44c957737bf422127283c08e['h03b86] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dc4] =  Ifd35529b44c957737bf422127283c08e['h03b88] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dc5] =  Ifd35529b44c957737bf422127283c08e['h03b8a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dc6] =  Ifd35529b44c957737bf422127283c08e['h03b8c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dc7] =  Ifd35529b44c957737bf422127283c08e['h03b8e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dc8] =  Ifd35529b44c957737bf422127283c08e['h03b90] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dc9] =  Ifd35529b44c957737bf422127283c08e['h03b92] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dca] =  Ifd35529b44c957737bf422127283c08e['h03b94] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dcb] =  Ifd35529b44c957737bf422127283c08e['h03b96] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dcc] =  Ifd35529b44c957737bf422127283c08e['h03b98] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dcd] =  Ifd35529b44c957737bf422127283c08e['h03b9a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dce] =  Ifd35529b44c957737bf422127283c08e['h03b9c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dcf] =  Ifd35529b44c957737bf422127283c08e['h03b9e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dd0] =  Ifd35529b44c957737bf422127283c08e['h03ba0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dd1] =  Ifd35529b44c957737bf422127283c08e['h03ba2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dd2] =  Ifd35529b44c957737bf422127283c08e['h03ba4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dd3] =  Ifd35529b44c957737bf422127283c08e['h03ba6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dd4] =  Ifd35529b44c957737bf422127283c08e['h03ba8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dd5] =  Ifd35529b44c957737bf422127283c08e['h03baa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dd6] =  Ifd35529b44c957737bf422127283c08e['h03bac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dd7] =  Ifd35529b44c957737bf422127283c08e['h03bae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dd8] =  Ifd35529b44c957737bf422127283c08e['h03bb0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dd9] =  Ifd35529b44c957737bf422127283c08e['h03bb2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dda] =  Ifd35529b44c957737bf422127283c08e['h03bb4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ddb] =  Ifd35529b44c957737bf422127283c08e['h03bb6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ddc] =  Ifd35529b44c957737bf422127283c08e['h03bb8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ddd] =  Ifd35529b44c957737bf422127283c08e['h03bba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dde] =  Ifd35529b44c957737bf422127283c08e['h03bbc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ddf] =  Ifd35529b44c957737bf422127283c08e['h03bbe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01de0] =  Ifd35529b44c957737bf422127283c08e['h03bc0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01de1] =  Ifd35529b44c957737bf422127283c08e['h03bc2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01de2] =  Ifd35529b44c957737bf422127283c08e['h03bc4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01de3] =  Ifd35529b44c957737bf422127283c08e['h03bc6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01de4] =  Ifd35529b44c957737bf422127283c08e['h03bc8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01de5] =  Ifd35529b44c957737bf422127283c08e['h03bca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01de6] =  Ifd35529b44c957737bf422127283c08e['h03bcc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01de7] =  Ifd35529b44c957737bf422127283c08e['h03bce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01de8] =  Ifd35529b44c957737bf422127283c08e['h03bd0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01de9] =  Ifd35529b44c957737bf422127283c08e['h03bd2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dea] =  Ifd35529b44c957737bf422127283c08e['h03bd4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01deb] =  Ifd35529b44c957737bf422127283c08e['h03bd6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dec] =  Ifd35529b44c957737bf422127283c08e['h03bd8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ded] =  Ifd35529b44c957737bf422127283c08e['h03bda] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dee] =  Ifd35529b44c957737bf422127283c08e['h03bdc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01def] =  Ifd35529b44c957737bf422127283c08e['h03bde] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01df0] =  Ifd35529b44c957737bf422127283c08e['h03be0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01df1] =  Ifd35529b44c957737bf422127283c08e['h03be2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01df2] =  Ifd35529b44c957737bf422127283c08e['h03be4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01df3] =  Ifd35529b44c957737bf422127283c08e['h03be6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01df4] =  Ifd35529b44c957737bf422127283c08e['h03be8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01df5] =  Ifd35529b44c957737bf422127283c08e['h03bea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01df6] =  Ifd35529b44c957737bf422127283c08e['h03bec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01df7] =  Ifd35529b44c957737bf422127283c08e['h03bee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01df8] =  Ifd35529b44c957737bf422127283c08e['h03bf0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01df9] =  Ifd35529b44c957737bf422127283c08e['h03bf2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dfa] =  Ifd35529b44c957737bf422127283c08e['h03bf4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dfb] =  Ifd35529b44c957737bf422127283c08e['h03bf6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dfc] =  Ifd35529b44c957737bf422127283c08e['h03bf8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dfd] =  Ifd35529b44c957737bf422127283c08e['h03bfa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dfe] =  Ifd35529b44c957737bf422127283c08e['h03bfc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01dff] =  Ifd35529b44c957737bf422127283c08e['h03bfe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e00] =  Ifd35529b44c957737bf422127283c08e['h03c00] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e01] =  Ifd35529b44c957737bf422127283c08e['h03c02] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e02] =  Ifd35529b44c957737bf422127283c08e['h03c04] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e03] =  Ifd35529b44c957737bf422127283c08e['h03c06] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e04] =  Ifd35529b44c957737bf422127283c08e['h03c08] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e05] =  Ifd35529b44c957737bf422127283c08e['h03c0a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e06] =  Ifd35529b44c957737bf422127283c08e['h03c0c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e07] =  Ifd35529b44c957737bf422127283c08e['h03c0e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e08] =  Ifd35529b44c957737bf422127283c08e['h03c10] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e09] =  Ifd35529b44c957737bf422127283c08e['h03c12] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e0a] =  Ifd35529b44c957737bf422127283c08e['h03c14] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e0b] =  Ifd35529b44c957737bf422127283c08e['h03c16] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e0c] =  Ifd35529b44c957737bf422127283c08e['h03c18] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e0d] =  Ifd35529b44c957737bf422127283c08e['h03c1a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e0e] =  Ifd35529b44c957737bf422127283c08e['h03c1c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e0f] =  Ifd35529b44c957737bf422127283c08e['h03c1e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e10] =  Ifd35529b44c957737bf422127283c08e['h03c20] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e11] =  Ifd35529b44c957737bf422127283c08e['h03c22] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e12] =  Ifd35529b44c957737bf422127283c08e['h03c24] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e13] =  Ifd35529b44c957737bf422127283c08e['h03c26] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e14] =  Ifd35529b44c957737bf422127283c08e['h03c28] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e15] =  Ifd35529b44c957737bf422127283c08e['h03c2a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e16] =  Ifd35529b44c957737bf422127283c08e['h03c2c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e17] =  Ifd35529b44c957737bf422127283c08e['h03c2e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e18] =  Ifd35529b44c957737bf422127283c08e['h03c30] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e19] =  Ifd35529b44c957737bf422127283c08e['h03c32] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e1a] =  Ifd35529b44c957737bf422127283c08e['h03c34] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e1b] =  Ifd35529b44c957737bf422127283c08e['h03c36] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e1c] =  Ifd35529b44c957737bf422127283c08e['h03c38] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e1d] =  Ifd35529b44c957737bf422127283c08e['h03c3a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e1e] =  Ifd35529b44c957737bf422127283c08e['h03c3c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e1f] =  Ifd35529b44c957737bf422127283c08e['h03c3e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e20] =  Ifd35529b44c957737bf422127283c08e['h03c40] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e21] =  Ifd35529b44c957737bf422127283c08e['h03c42] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e22] =  Ifd35529b44c957737bf422127283c08e['h03c44] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e23] =  Ifd35529b44c957737bf422127283c08e['h03c46] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e24] =  Ifd35529b44c957737bf422127283c08e['h03c48] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e25] =  Ifd35529b44c957737bf422127283c08e['h03c4a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e26] =  Ifd35529b44c957737bf422127283c08e['h03c4c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e27] =  Ifd35529b44c957737bf422127283c08e['h03c4e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e28] =  Ifd35529b44c957737bf422127283c08e['h03c50] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e29] =  Ifd35529b44c957737bf422127283c08e['h03c52] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e2a] =  Ifd35529b44c957737bf422127283c08e['h03c54] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e2b] =  Ifd35529b44c957737bf422127283c08e['h03c56] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e2c] =  Ifd35529b44c957737bf422127283c08e['h03c58] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e2d] =  Ifd35529b44c957737bf422127283c08e['h03c5a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e2e] =  Ifd35529b44c957737bf422127283c08e['h03c5c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e2f] =  Ifd35529b44c957737bf422127283c08e['h03c5e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e30] =  Ifd35529b44c957737bf422127283c08e['h03c60] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e31] =  Ifd35529b44c957737bf422127283c08e['h03c62] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e32] =  Ifd35529b44c957737bf422127283c08e['h03c64] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e33] =  Ifd35529b44c957737bf422127283c08e['h03c66] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e34] =  Ifd35529b44c957737bf422127283c08e['h03c68] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e35] =  Ifd35529b44c957737bf422127283c08e['h03c6a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e36] =  Ifd35529b44c957737bf422127283c08e['h03c6c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e37] =  Ifd35529b44c957737bf422127283c08e['h03c6e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e38] =  Ifd35529b44c957737bf422127283c08e['h03c70] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e39] =  Ifd35529b44c957737bf422127283c08e['h03c72] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e3a] =  Ifd35529b44c957737bf422127283c08e['h03c74] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e3b] =  Ifd35529b44c957737bf422127283c08e['h03c76] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e3c] =  Ifd35529b44c957737bf422127283c08e['h03c78] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e3d] =  Ifd35529b44c957737bf422127283c08e['h03c7a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e3e] =  Ifd35529b44c957737bf422127283c08e['h03c7c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e3f] =  Ifd35529b44c957737bf422127283c08e['h03c7e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e40] =  Ifd35529b44c957737bf422127283c08e['h03c80] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e41] =  Ifd35529b44c957737bf422127283c08e['h03c82] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e42] =  Ifd35529b44c957737bf422127283c08e['h03c84] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e43] =  Ifd35529b44c957737bf422127283c08e['h03c86] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e44] =  Ifd35529b44c957737bf422127283c08e['h03c88] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e45] =  Ifd35529b44c957737bf422127283c08e['h03c8a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e46] =  Ifd35529b44c957737bf422127283c08e['h03c8c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e47] =  Ifd35529b44c957737bf422127283c08e['h03c8e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e48] =  Ifd35529b44c957737bf422127283c08e['h03c90] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e49] =  Ifd35529b44c957737bf422127283c08e['h03c92] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e4a] =  Ifd35529b44c957737bf422127283c08e['h03c94] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e4b] =  Ifd35529b44c957737bf422127283c08e['h03c96] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e4c] =  Ifd35529b44c957737bf422127283c08e['h03c98] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e4d] =  Ifd35529b44c957737bf422127283c08e['h03c9a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e4e] =  Ifd35529b44c957737bf422127283c08e['h03c9c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e4f] =  Ifd35529b44c957737bf422127283c08e['h03c9e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e50] =  Ifd35529b44c957737bf422127283c08e['h03ca0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e51] =  Ifd35529b44c957737bf422127283c08e['h03ca2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e52] =  Ifd35529b44c957737bf422127283c08e['h03ca4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e53] =  Ifd35529b44c957737bf422127283c08e['h03ca6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e54] =  Ifd35529b44c957737bf422127283c08e['h03ca8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e55] =  Ifd35529b44c957737bf422127283c08e['h03caa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e56] =  Ifd35529b44c957737bf422127283c08e['h03cac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e57] =  Ifd35529b44c957737bf422127283c08e['h03cae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e58] =  Ifd35529b44c957737bf422127283c08e['h03cb0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e59] =  Ifd35529b44c957737bf422127283c08e['h03cb2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e5a] =  Ifd35529b44c957737bf422127283c08e['h03cb4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e5b] =  Ifd35529b44c957737bf422127283c08e['h03cb6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e5c] =  Ifd35529b44c957737bf422127283c08e['h03cb8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e5d] =  Ifd35529b44c957737bf422127283c08e['h03cba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e5e] =  Ifd35529b44c957737bf422127283c08e['h03cbc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e5f] =  Ifd35529b44c957737bf422127283c08e['h03cbe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e60] =  Ifd35529b44c957737bf422127283c08e['h03cc0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e61] =  Ifd35529b44c957737bf422127283c08e['h03cc2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e62] =  Ifd35529b44c957737bf422127283c08e['h03cc4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e63] =  Ifd35529b44c957737bf422127283c08e['h03cc6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e64] =  Ifd35529b44c957737bf422127283c08e['h03cc8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e65] =  Ifd35529b44c957737bf422127283c08e['h03cca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e66] =  Ifd35529b44c957737bf422127283c08e['h03ccc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e67] =  Ifd35529b44c957737bf422127283c08e['h03cce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e68] =  Ifd35529b44c957737bf422127283c08e['h03cd0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e69] =  Ifd35529b44c957737bf422127283c08e['h03cd2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e6a] =  Ifd35529b44c957737bf422127283c08e['h03cd4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e6b] =  Ifd35529b44c957737bf422127283c08e['h03cd6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e6c] =  Ifd35529b44c957737bf422127283c08e['h03cd8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e6d] =  Ifd35529b44c957737bf422127283c08e['h03cda] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e6e] =  Ifd35529b44c957737bf422127283c08e['h03cdc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e6f] =  Ifd35529b44c957737bf422127283c08e['h03cde] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e70] =  Ifd35529b44c957737bf422127283c08e['h03ce0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e71] =  Ifd35529b44c957737bf422127283c08e['h03ce2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e72] =  Ifd35529b44c957737bf422127283c08e['h03ce4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e73] =  Ifd35529b44c957737bf422127283c08e['h03ce6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e74] =  Ifd35529b44c957737bf422127283c08e['h03ce8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e75] =  Ifd35529b44c957737bf422127283c08e['h03cea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e76] =  Ifd35529b44c957737bf422127283c08e['h03cec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e77] =  Ifd35529b44c957737bf422127283c08e['h03cee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e78] =  Ifd35529b44c957737bf422127283c08e['h03cf0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e79] =  Ifd35529b44c957737bf422127283c08e['h03cf2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e7a] =  Ifd35529b44c957737bf422127283c08e['h03cf4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e7b] =  Ifd35529b44c957737bf422127283c08e['h03cf6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e7c] =  Ifd35529b44c957737bf422127283c08e['h03cf8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e7d] =  Ifd35529b44c957737bf422127283c08e['h03cfa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e7e] =  Ifd35529b44c957737bf422127283c08e['h03cfc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e7f] =  Ifd35529b44c957737bf422127283c08e['h03cfe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e80] =  Ifd35529b44c957737bf422127283c08e['h03d00] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e81] =  Ifd35529b44c957737bf422127283c08e['h03d02] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e82] =  Ifd35529b44c957737bf422127283c08e['h03d04] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e83] =  Ifd35529b44c957737bf422127283c08e['h03d06] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e84] =  Ifd35529b44c957737bf422127283c08e['h03d08] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e85] =  Ifd35529b44c957737bf422127283c08e['h03d0a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e86] =  Ifd35529b44c957737bf422127283c08e['h03d0c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e87] =  Ifd35529b44c957737bf422127283c08e['h03d0e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e88] =  Ifd35529b44c957737bf422127283c08e['h03d10] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e89] =  Ifd35529b44c957737bf422127283c08e['h03d12] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e8a] =  Ifd35529b44c957737bf422127283c08e['h03d14] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e8b] =  Ifd35529b44c957737bf422127283c08e['h03d16] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e8c] =  Ifd35529b44c957737bf422127283c08e['h03d18] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e8d] =  Ifd35529b44c957737bf422127283c08e['h03d1a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e8e] =  Ifd35529b44c957737bf422127283c08e['h03d1c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e8f] =  Ifd35529b44c957737bf422127283c08e['h03d1e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e90] =  Ifd35529b44c957737bf422127283c08e['h03d20] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e91] =  Ifd35529b44c957737bf422127283c08e['h03d22] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e92] =  Ifd35529b44c957737bf422127283c08e['h03d24] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e93] =  Ifd35529b44c957737bf422127283c08e['h03d26] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e94] =  Ifd35529b44c957737bf422127283c08e['h03d28] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e95] =  Ifd35529b44c957737bf422127283c08e['h03d2a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e96] =  Ifd35529b44c957737bf422127283c08e['h03d2c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e97] =  Ifd35529b44c957737bf422127283c08e['h03d2e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e98] =  Ifd35529b44c957737bf422127283c08e['h03d30] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e99] =  Ifd35529b44c957737bf422127283c08e['h03d32] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e9a] =  Ifd35529b44c957737bf422127283c08e['h03d34] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e9b] =  Ifd35529b44c957737bf422127283c08e['h03d36] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e9c] =  Ifd35529b44c957737bf422127283c08e['h03d38] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e9d] =  Ifd35529b44c957737bf422127283c08e['h03d3a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e9e] =  Ifd35529b44c957737bf422127283c08e['h03d3c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01e9f] =  Ifd35529b44c957737bf422127283c08e['h03d3e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ea0] =  Ifd35529b44c957737bf422127283c08e['h03d40] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ea1] =  Ifd35529b44c957737bf422127283c08e['h03d42] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ea2] =  Ifd35529b44c957737bf422127283c08e['h03d44] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ea3] =  Ifd35529b44c957737bf422127283c08e['h03d46] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ea4] =  Ifd35529b44c957737bf422127283c08e['h03d48] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ea5] =  Ifd35529b44c957737bf422127283c08e['h03d4a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ea6] =  Ifd35529b44c957737bf422127283c08e['h03d4c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ea7] =  Ifd35529b44c957737bf422127283c08e['h03d4e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ea8] =  Ifd35529b44c957737bf422127283c08e['h03d50] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ea9] =  Ifd35529b44c957737bf422127283c08e['h03d52] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01eaa] =  Ifd35529b44c957737bf422127283c08e['h03d54] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01eab] =  Ifd35529b44c957737bf422127283c08e['h03d56] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01eac] =  Ifd35529b44c957737bf422127283c08e['h03d58] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ead] =  Ifd35529b44c957737bf422127283c08e['h03d5a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01eae] =  Ifd35529b44c957737bf422127283c08e['h03d5c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01eaf] =  Ifd35529b44c957737bf422127283c08e['h03d5e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01eb0] =  Ifd35529b44c957737bf422127283c08e['h03d60] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01eb1] =  Ifd35529b44c957737bf422127283c08e['h03d62] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01eb2] =  Ifd35529b44c957737bf422127283c08e['h03d64] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01eb3] =  Ifd35529b44c957737bf422127283c08e['h03d66] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01eb4] =  Ifd35529b44c957737bf422127283c08e['h03d68] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01eb5] =  Ifd35529b44c957737bf422127283c08e['h03d6a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01eb6] =  Ifd35529b44c957737bf422127283c08e['h03d6c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01eb7] =  Ifd35529b44c957737bf422127283c08e['h03d6e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01eb8] =  Ifd35529b44c957737bf422127283c08e['h03d70] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01eb9] =  Ifd35529b44c957737bf422127283c08e['h03d72] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01eba] =  Ifd35529b44c957737bf422127283c08e['h03d74] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ebb] =  Ifd35529b44c957737bf422127283c08e['h03d76] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ebc] =  Ifd35529b44c957737bf422127283c08e['h03d78] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ebd] =  Ifd35529b44c957737bf422127283c08e['h03d7a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ebe] =  Ifd35529b44c957737bf422127283c08e['h03d7c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ebf] =  Ifd35529b44c957737bf422127283c08e['h03d7e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ec0] =  Ifd35529b44c957737bf422127283c08e['h03d80] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ec1] =  Ifd35529b44c957737bf422127283c08e['h03d82] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ec2] =  Ifd35529b44c957737bf422127283c08e['h03d84] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ec3] =  Ifd35529b44c957737bf422127283c08e['h03d86] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ec4] =  Ifd35529b44c957737bf422127283c08e['h03d88] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ec5] =  Ifd35529b44c957737bf422127283c08e['h03d8a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ec6] =  Ifd35529b44c957737bf422127283c08e['h03d8c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ec7] =  Ifd35529b44c957737bf422127283c08e['h03d8e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ec8] =  Ifd35529b44c957737bf422127283c08e['h03d90] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ec9] =  Ifd35529b44c957737bf422127283c08e['h03d92] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01eca] =  Ifd35529b44c957737bf422127283c08e['h03d94] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ecb] =  Ifd35529b44c957737bf422127283c08e['h03d96] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ecc] =  Ifd35529b44c957737bf422127283c08e['h03d98] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ecd] =  Ifd35529b44c957737bf422127283c08e['h03d9a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ece] =  Ifd35529b44c957737bf422127283c08e['h03d9c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ecf] =  Ifd35529b44c957737bf422127283c08e['h03d9e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ed0] =  Ifd35529b44c957737bf422127283c08e['h03da0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ed1] =  Ifd35529b44c957737bf422127283c08e['h03da2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ed2] =  Ifd35529b44c957737bf422127283c08e['h03da4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ed3] =  Ifd35529b44c957737bf422127283c08e['h03da6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ed4] =  Ifd35529b44c957737bf422127283c08e['h03da8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ed5] =  Ifd35529b44c957737bf422127283c08e['h03daa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ed6] =  Ifd35529b44c957737bf422127283c08e['h03dac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ed7] =  Ifd35529b44c957737bf422127283c08e['h03dae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ed8] =  Ifd35529b44c957737bf422127283c08e['h03db0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ed9] =  Ifd35529b44c957737bf422127283c08e['h03db2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01eda] =  Ifd35529b44c957737bf422127283c08e['h03db4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01edb] =  Ifd35529b44c957737bf422127283c08e['h03db6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01edc] =  Ifd35529b44c957737bf422127283c08e['h03db8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01edd] =  Ifd35529b44c957737bf422127283c08e['h03dba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ede] =  Ifd35529b44c957737bf422127283c08e['h03dbc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01edf] =  Ifd35529b44c957737bf422127283c08e['h03dbe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ee0] =  Ifd35529b44c957737bf422127283c08e['h03dc0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ee1] =  Ifd35529b44c957737bf422127283c08e['h03dc2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ee2] =  Ifd35529b44c957737bf422127283c08e['h03dc4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ee3] =  Ifd35529b44c957737bf422127283c08e['h03dc6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ee4] =  Ifd35529b44c957737bf422127283c08e['h03dc8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ee5] =  Ifd35529b44c957737bf422127283c08e['h03dca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ee6] =  Ifd35529b44c957737bf422127283c08e['h03dcc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ee7] =  Ifd35529b44c957737bf422127283c08e['h03dce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ee8] =  Ifd35529b44c957737bf422127283c08e['h03dd0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ee9] =  Ifd35529b44c957737bf422127283c08e['h03dd2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01eea] =  Ifd35529b44c957737bf422127283c08e['h03dd4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01eeb] =  Ifd35529b44c957737bf422127283c08e['h03dd6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01eec] =  Ifd35529b44c957737bf422127283c08e['h03dd8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01eed] =  Ifd35529b44c957737bf422127283c08e['h03dda] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01eee] =  Ifd35529b44c957737bf422127283c08e['h03ddc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01eef] =  Ifd35529b44c957737bf422127283c08e['h03dde] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ef0] =  Ifd35529b44c957737bf422127283c08e['h03de0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ef1] =  Ifd35529b44c957737bf422127283c08e['h03de2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ef2] =  Ifd35529b44c957737bf422127283c08e['h03de4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ef3] =  Ifd35529b44c957737bf422127283c08e['h03de6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ef4] =  Ifd35529b44c957737bf422127283c08e['h03de8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ef5] =  Ifd35529b44c957737bf422127283c08e['h03dea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ef6] =  Ifd35529b44c957737bf422127283c08e['h03dec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ef7] =  Ifd35529b44c957737bf422127283c08e['h03dee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ef8] =  Ifd35529b44c957737bf422127283c08e['h03df0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ef9] =  Ifd35529b44c957737bf422127283c08e['h03df2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01efa] =  Ifd35529b44c957737bf422127283c08e['h03df4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01efb] =  Ifd35529b44c957737bf422127283c08e['h03df6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01efc] =  Ifd35529b44c957737bf422127283c08e['h03df8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01efd] =  Ifd35529b44c957737bf422127283c08e['h03dfa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01efe] =  Ifd35529b44c957737bf422127283c08e['h03dfc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01eff] =  Ifd35529b44c957737bf422127283c08e['h03dfe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f00] =  Ifd35529b44c957737bf422127283c08e['h03e00] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f01] =  Ifd35529b44c957737bf422127283c08e['h03e02] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f02] =  Ifd35529b44c957737bf422127283c08e['h03e04] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f03] =  Ifd35529b44c957737bf422127283c08e['h03e06] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f04] =  Ifd35529b44c957737bf422127283c08e['h03e08] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f05] =  Ifd35529b44c957737bf422127283c08e['h03e0a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f06] =  Ifd35529b44c957737bf422127283c08e['h03e0c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f07] =  Ifd35529b44c957737bf422127283c08e['h03e0e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f08] =  Ifd35529b44c957737bf422127283c08e['h03e10] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f09] =  Ifd35529b44c957737bf422127283c08e['h03e12] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f0a] =  Ifd35529b44c957737bf422127283c08e['h03e14] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f0b] =  Ifd35529b44c957737bf422127283c08e['h03e16] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f0c] =  Ifd35529b44c957737bf422127283c08e['h03e18] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f0d] =  Ifd35529b44c957737bf422127283c08e['h03e1a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f0e] =  Ifd35529b44c957737bf422127283c08e['h03e1c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f0f] =  Ifd35529b44c957737bf422127283c08e['h03e1e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f10] =  Ifd35529b44c957737bf422127283c08e['h03e20] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f11] =  Ifd35529b44c957737bf422127283c08e['h03e22] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f12] =  Ifd35529b44c957737bf422127283c08e['h03e24] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f13] =  Ifd35529b44c957737bf422127283c08e['h03e26] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f14] =  Ifd35529b44c957737bf422127283c08e['h03e28] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f15] =  Ifd35529b44c957737bf422127283c08e['h03e2a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f16] =  Ifd35529b44c957737bf422127283c08e['h03e2c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f17] =  Ifd35529b44c957737bf422127283c08e['h03e2e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f18] =  Ifd35529b44c957737bf422127283c08e['h03e30] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f19] =  Ifd35529b44c957737bf422127283c08e['h03e32] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f1a] =  Ifd35529b44c957737bf422127283c08e['h03e34] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f1b] =  Ifd35529b44c957737bf422127283c08e['h03e36] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f1c] =  Ifd35529b44c957737bf422127283c08e['h03e38] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f1d] =  Ifd35529b44c957737bf422127283c08e['h03e3a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f1e] =  Ifd35529b44c957737bf422127283c08e['h03e3c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f1f] =  Ifd35529b44c957737bf422127283c08e['h03e3e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f20] =  Ifd35529b44c957737bf422127283c08e['h03e40] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f21] =  Ifd35529b44c957737bf422127283c08e['h03e42] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f22] =  Ifd35529b44c957737bf422127283c08e['h03e44] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f23] =  Ifd35529b44c957737bf422127283c08e['h03e46] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f24] =  Ifd35529b44c957737bf422127283c08e['h03e48] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f25] =  Ifd35529b44c957737bf422127283c08e['h03e4a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f26] =  Ifd35529b44c957737bf422127283c08e['h03e4c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f27] =  Ifd35529b44c957737bf422127283c08e['h03e4e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f28] =  Ifd35529b44c957737bf422127283c08e['h03e50] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f29] =  Ifd35529b44c957737bf422127283c08e['h03e52] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f2a] =  Ifd35529b44c957737bf422127283c08e['h03e54] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f2b] =  Ifd35529b44c957737bf422127283c08e['h03e56] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f2c] =  Ifd35529b44c957737bf422127283c08e['h03e58] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f2d] =  Ifd35529b44c957737bf422127283c08e['h03e5a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f2e] =  Ifd35529b44c957737bf422127283c08e['h03e5c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f2f] =  Ifd35529b44c957737bf422127283c08e['h03e5e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f30] =  Ifd35529b44c957737bf422127283c08e['h03e60] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f31] =  Ifd35529b44c957737bf422127283c08e['h03e62] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f32] =  Ifd35529b44c957737bf422127283c08e['h03e64] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f33] =  Ifd35529b44c957737bf422127283c08e['h03e66] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f34] =  Ifd35529b44c957737bf422127283c08e['h03e68] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f35] =  Ifd35529b44c957737bf422127283c08e['h03e6a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f36] =  Ifd35529b44c957737bf422127283c08e['h03e6c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f37] =  Ifd35529b44c957737bf422127283c08e['h03e6e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f38] =  Ifd35529b44c957737bf422127283c08e['h03e70] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f39] =  Ifd35529b44c957737bf422127283c08e['h03e72] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f3a] =  Ifd35529b44c957737bf422127283c08e['h03e74] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f3b] =  Ifd35529b44c957737bf422127283c08e['h03e76] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f3c] =  Ifd35529b44c957737bf422127283c08e['h03e78] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f3d] =  Ifd35529b44c957737bf422127283c08e['h03e7a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f3e] =  Ifd35529b44c957737bf422127283c08e['h03e7c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f3f] =  Ifd35529b44c957737bf422127283c08e['h03e7e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f40] =  Ifd35529b44c957737bf422127283c08e['h03e80] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f41] =  Ifd35529b44c957737bf422127283c08e['h03e82] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f42] =  Ifd35529b44c957737bf422127283c08e['h03e84] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f43] =  Ifd35529b44c957737bf422127283c08e['h03e86] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f44] =  Ifd35529b44c957737bf422127283c08e['h03e88] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f45] =  Ifd35529b44c957737bf422127283c08e['h03e8a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f46] =  Ifd35529b44c957737bf422127283c08e['h03e8c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f47] =  Ifd35529b44c957737bf422127283c08e['h03e8e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f48] =  Ifd35529b44c957737bf422127283c08e['h03e90] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f49] =  Ifd35529b44c957737bf422127283c08e['h03e92] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f4a] =  Ifd35529b44c957737bf422127283c08e['h03e94] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f4b] =  Ifd35529b44c957737bf422127283c08e['h03e96] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f4c] =  Ifd35529b44c957737bf422127283c08e['h03e98] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f4d] =  Ifd35529b44c957737bf422127283c08e['h03e9a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f4e] =  Ifd35529b44c957737bf422127283c08e['h03e9c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f4f] =  Ifd35529b44c957737bf422127283c08e['h03e9e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f50] =  Ifd35529b44c957737bf422127283c08e['h03ea0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f51] =  Ifd35529b44c957737bf422127283c08e['h03ea2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f52] =  Ifd35529b44c957737bf422127283c08e['h03ea4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f53] =  Ifd35529b44c957737bf422127283c08e['h03ea6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f54] =  Ifd35529b44c957737bf422127283c08e['h03ea8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f55] =  Ifd35529b44c957737bf422127283c08e['h03eaa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f56] =  Ifd35529b44c957737bf422127283c08e['h03eac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f57] =  Ifd35529b44c957737bf422127283c08e['h03eae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f58] =  Ifd35529b44c957737bf422127283c08e['h03eb0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f59] =  Ifd35529b44c957737bf422127283c08e['h03eb2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f5a] =  Ifd35529b44c957737bf422127283c08e['h03eb4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f5b] =  Ifd35529b44c957737bf422127283c08e['h03eb6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f5c] =  Ifd35529b44c957737bf422127283c08e['h03eb8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f5d] =  Ifd35529b44c957737bf422127283c08e['h03eba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f5e] =  Ifd35529b44c957737bf422127283c08e['h03ebc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f5f] =  Ifd35529b44c957737bf422127283c08e['h03ebe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f60] =  Ifd35529b44c957737bf422127283c08e['h03ec0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f61] =  Ifd35529b44c957737bf422127283c08e['h03ec2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f62] =  Ifd35529b44c957737bf422127283c08e['h03ec4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f63] =  Ifd35529b44c957737bf422127283c08e['h03ec6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f64] =  Ifd35529b44c957737bf422127283c08e['h03ec8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f65] =  Ifd35529b44c957737bf422127283c08e['h03eca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f66] =  Ifd35529b44c957737bf422127283c08e['h03ecc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f67] =  Ifd35529b44c957737bf422127283c08e['h03ece] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f68] =  Ifd35529b44c957737bf422127283c08e['h03ed0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f69] =  Ifd35529b44c957737bf422127283c08e['h03ed2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f6a] =  Ifd35529b44c957737bf422127283c08e['h03ed4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f6b] =  Ifd35529b44c957737bf422127283c08e['h03ed6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f6c] =  Ifd35529b44c957737bf422127283c08e['h03ed8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f6d] =  Ifd35529b44c957737bf422127283c08e['h03eda] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f6e] =  Ifd35529b44c957737bf422127283c08e['h03edc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f6f] =  Ifd35529b44c957737bf422127283c08e['h03ede] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f70] =  Ifd35529b44c957737bf422127283c08e['h03ee0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f71] =  Ifd35529b44c957737bf422127283c08e['h03ee2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f72] =  Ifd35529b44c957737bf422127283c08e['h03ee4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f73] =  Ifd35529b44c957737bf422127283c08e['h03ee6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f74] =  Ifd35529b44c957737bf422127283c08e['h03ee8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f75] =  Ifd35529b44c957737bf422127283c08e['h03eea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f76] =  Ifd35529b44c957737bf422127283c08e['h03eec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f77] =  Ifd35529b44c957737bf422127283c08e['h03eee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f78] =  Ifd35529b44c957737bf422127283c08e['h03ef0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f79] =  Ifd35529b44c957737bf422127283c08e['h03ef2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f7a] =  Ifd35529b44c957737bf422127283c08e['h03ef4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f7b] =  Ifd35529b44c957737bf422127283c08e['h03ef6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f7c] =  Ifd35529b44c957737bf422127283c08e['h03ef8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f7d] =  Ifd35529b44c957737bf422127283c08e['h03efa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f7e] =  Ifd35529b44c957737bf422127283c08e['h03efc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f7f] =  Ifd35529b44c957737bf422127283c08e['h03efe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f80] =  Ifd35529b44c957737bf422127283c08e['h03f00] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f81] =  Ifd35529b44c957737bf422127283c08e['h03f02] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f82] =  Ifd35529b44c957737bf422127283c08e['h03f04] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f83] =  Ifd35529b44c957737bf422127283c08e['h03f06] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f84] =  Ifd35529b44c957737bf422127283c08e['h03f08] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f85] =  Ifd35529b44c957737bf422127283c08e['h03f0a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f86] =  Ifd35529b44c957737bf422127283c08e['h03f0c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f87] =  Ifd35529b44c957737bf422127283c08e['h03f0e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f88] =  Ifd35529b44c957737bf422127283c08e['h03f10] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f89] =  Ifd35529b44c957737bf422127283c08e['h03f12] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f8a] =  Ifd35529b44c957737bf422127283c08e['h03f14] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f8b] =  Ifd35529b44c957737bf422127283c08e['h03f16] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f8c] =  Ifd35529b44c957737bf422127283c08e['h03f18] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f8d] =  Ifd35529b44c957737bf422127283c08e['h03f1a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f8e] =  Ifd35529b44c957737bf422127283c08e['h03f1c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f8f] =  Ifd35529b44c957737bf422127283c08e['h03f1e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f90] =  Ifd35529b44c957737bf422127283c08e['h03f20] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f91] =  Ifd35529b44c957737bf422127283c08e['h03f22] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f92] =  Ifd35529b44c957737bf422127283c08e['h03f24] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f93] =  Ifd35529b44c957737bf422127283c08e['h03f26] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f94] =  Ifd35529b44c957737bf422127283c08e['h03f28] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f95] =  Ifd35529b44c957737bf422127283c08e['h03f2a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f96] =  Ifd35529b44c957737bf422127283c08e['h03f2c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f97] =  Ifd35529b44c957737bf422127283c08e['h03f2e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f98] =  Ifd35529b44c957737bf422127283c08e['h03f30] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f99] =  Ifd35529b44c957737bf422127283c08e['h03f32] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f9a] =  Ifd35529b44c957737bf422127283c08e['h03f34] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f9b] =  Ifd35529b44c957737bf422127283c08e['h03f36] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f9c] =  Ifd35529b44c957737bf422127283c08e['h03f38] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f9d] =  Ifd35529b44c957737bf422127283c08e['h03f3a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f9e] =  Ifd35529b44c957737bf422127283c08e['h03f3c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01f9f] =  Ifd35529b44c957737bf422127283c08e['h03f3e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fa0] =  Ifd35529b44c957737bf422127283c08e['h03f40] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fa1] =  Ifd35529b44c957737bf422127283c08e['h03f42] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fa2] =  Ifd35529b44c957737bf422127283c08e['h03f44] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fa3] =  Ifd35529b44c957737bf422127283c08e['h03f46] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fa4] =  Ifd35529b44c957737bf422127283c08e['h03f48] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fa5] =  Ifd35529b44c957737bf422127283c08e['h03f4a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fa6] =  Ifd35529b44c957737bf422127283c08e['h03f4c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fa7] =  Ifd35529b44c957737bf422127283c08e['h03f4e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fa8] =  Ifd35529b44c957737bf422127283c08e['h03f50] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fa9] =  Ifd35529b44c957737bf422127283c08e['h03f52] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01faa] =  Ifd35529b44c957737bf422127283c08e['h03f54] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fab] =  Ifd35529b44c957737bf422127283c08e['h03f56] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fac] =  Ifd35529b44c957737bf422127283c08e['h03f58] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fad] =  Ifd35529b44c957737bf422127283c08e['h03f5a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fae] =  Ifd35529b44c957737bf422127283c08e['h03f5c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01faf] =  Ifd35529b44c957737bf422127283c08e['h03f5e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fb0] =  Ifd35529b44c957737bf422127283c08e['h03f60] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fb1] =  Ifd35529b44c957737bf422127283c08e['h03f62] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fb2] =  Ifd35529b44c957737bf422127283c08e['h03f64] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fb3] =  Ifd35529b44c957737bf422127283c08e['h03f66] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fb4] =  Ifd35529b44c957737bf422127283c08e['h03f68] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fb5] =  Ifd35529b44c957737bf422127283c08e['h03f6a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fb6] =  Ifd35529b44c957737bf422127283c08e['h03f6c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fb7] =  Ifd35529b44c957737bf422127283c08e['h03f6e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fb8] =  Ifd35529b44c957737bf422127283c08e['h03f70] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fb9] =  Ifd35529b44c957737bf422127283c08e['h03f72] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fba] =  Ifd35529b44c957737bf422127283c08e['h03f74] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fbb] =  Ifd35529b44c957737bf422127283c08e['h03f76] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fbc] =  Ifd35529b44c957737bf422127283c08e['h03f78] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fbd] =  Ifd35529b44c957737bf422127283c08e['h03f7a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fbe] =  Ifd35529b44c957737bf422127283c08e['h03f7c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fbf] =  Ifd35529b44c957737bf422127283c08e['h03f7e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fc0] =  Ifd35529b44c957737bf422127283c08e['h03f80] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fc1] =  Ifd35529b44c957737bf422127283c08e['h03f82] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fc2] =  Ifd35529b44c957737bf422127283c08e['h03f84] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fc3] =  Ifd35529b44c957737bf422127283c08e['h03f86] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fc4] =  Ifd35529b44c957737bf422127283c08e['h03f88] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fc5] =  Ifd35529b44c957737bf422127283c08e['h03f8a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fc6] =  Ifd35529b44c957737bf422127283c08e['h03f8c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fc7] =  Ifd35529b44c957737bf422127283c08e['h03f8e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fc8] =  Ifd35529b44c957737bf422127283c08e['h03f90] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fc9] =  Ifd35529b44c957737bf422127283c08e['h03f92] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fca] =  Ifd35529b44c957737bf422127283c08e['h03f94] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fcb] =  Ifd35529b44c957737bf422127283c08e['h03f96] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fcc] =  Ifd35529b44c957737bf422127283c08e['h03f98] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fcd] =  Ifd35529b44c957737bf422127283c08e['h03f9a] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fce] =  Ifd35529b44c957737bf422127283c08e['h03f9c] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fcf] =  Ifd35529b44c957737bf422127283c08e['h03f9e] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fd0] =  Ifd35529b44c957737bf422127283c08e['h03fa0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fd1] =  Ifd35529b44c957737bf422127283c08e['h03fa2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fd2] =  Ifd35529b44c957737bf422127283c08e['h03fa4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fd3] =  Ifd35529b44c957737bf422127283c08e['h03fa6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fd4] =  Ifd35529b44c957737bf422127283c08e['h03fa8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fd5] =  Ifd35529b44c957737bf422127283c08e['h03faa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fd6] =  Ifd35529b44c957737bf422127283c08e['h03fac] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fd7] =  Ifd35529b44c957737bf422127283c08e['h03fae] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fd8] =  Ifd35529b44c957737bf422127283c08e['h03fb0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fd9] =  Ifd35529b44c957737bf422127283c08e['h03fb2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fda] =  Ifd35529b44c957737bf422127283c08e['h03fb4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fdb] =  Ifd35529b44c957737bf422127283c08e['h03fb6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fdc] =  Ifd35529b44c957737bf422127283c08e['h03fb8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fdd] =  Ifd35529b44c957737bf422127283c08e['h03fba] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fde] =  Ifd35529b44c957737bf422127283c08e['h03fbc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fdf] =  Ifd35529b44c957737bf422127283c08e['h03fbe] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fe0] =  Ifd35529b44c957737bf422127283c08e['h03fc0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fe1] =  Ifd35529b44c957737bf422127283c08e['h03fc2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fe2] =  Ifd35529b44c957737bf422127283c08e['h03fc4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fe3] =  Ifd35529b44c957737bf422127283c08e['h03fc6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fe4] =  Ifd35529b44c957737bf422127283c08e['h03fc8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fe5] =  Ifd35529b44c957737bf422127283c08e['h03fca] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fe6] =  Ifd35529b44c957737bf422127283c08e['h03fcc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fe7] =  Ifd35529b44c957737bf422127283c08e['h03fce] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fe8] =  Ifd35529b44c957737bf422127283c08e['h03fd0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fe9] =  Ifd35529b44c957737bf422127283c08e['h03fd2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fea] =  Ifd35529b44c957737bf422127283c08e['h03fd4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01feb] =  Ifd35529b44c957737bf422127283c08e['h03fd6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fec] =  Ifd35529b44c957737bf422127283c08e['h03fd8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fed] =  Ifd35529b44c957737bf422127283c08e['h03fda] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fee] =  Ifd35529b44c957737bf422127283c08e['h03fdc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fef] =  Ifd35529b44c957737bf422127283c08e['h03fde] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ff0] =  Ifd35529b44c957737bf422127283c08e['h03fe0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ff1] =  Ifd35529b44c957737bf422127283c08e['h03fe2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ff2] =  Ifd35529b44c957737bf422127283c08e['h03fe4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ff3] =  Ifd35529b44c957737bf422127283c08e['h03fe6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ff4] =  Ifd35529b44c957737bf422127283c08e['h03fe8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ff5] =  Ifd35529b44c957737bf422127283c08e['h03fea] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ff6] =  Ifd35529b44c957737bf422127283c08e['h03fec] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ff7] =  Ifd35529b44c957737bf422127283c08e['h03fee] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ff8] =  Ifd35529b44c957737bf422127283c08e['h03ff0] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ff9] =  Ifd35529b44c957737bf422127283c08e['h03ff2] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ffa] =  Ifd35529b44c957737bf422127283c08e['h03ff4] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ffb] =  Ifd35529b44c957737bf422127283c08e['h03ff6] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ffc] =  Ifd35529b44c957737bf422127283c08e['h03ff8] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ffd] =  Ifd35529b44c957737bf422127283c08e['h03ffa] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01ffe] =  Ifd35529b44c957737bf422127283c08e['h03ffc] ;
//end
//always_comb begin // 
               If409768b648a33a7ed878a070d4f6251['h01fff] =  Ifd35529b44c957737bf422127283c08e['h03ffe] ;
//end
