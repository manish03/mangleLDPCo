reg [flogtanh_WDTH -1:0] I5615abbd072d30da52163f16f1980957, I148a2b6bf6253f900182125f4f086010;
reg [flogtanh_WDTH -1:0] Ie7e694e2f86689b06efbd2eb66c5ffd8, I23d8325c203e2a9e4118ea94210effa0;
reg [flogtanh_WDTH -1:0] Id0287bb263a65d5eea34cbd5be2cfe3d, I9cdc23307c28dd846a7981b6a1b8552e;
reg [flogtanh_WDTH -1:0] Ic223bac65f3241d30afc2e21178eebfc, I2b9e2a2b9bea3cdd0c7b48f864254aa8;
reg [flogtanh_WDTH -1:0] I22794d7d1503d8cf477ad8b189d53ace, I0da340314517b5042829528ed7621d8f;
reg [flogtanh_WDTH -1:0] I8ccd9901d0629218945ab24f6eea34a3, I4edefd1be2348543f0e11dbce5623271;
reg [flogtanh_WDTH -1:0] Ifdeb82639682ca4a87f76e40a181bf79, I8315a1e97dcb0458031c17b029afac99;
reg [flogtanh_WDTH -1:0] Ib1879574e569ce9d6787132cc87e8de4, I2b91900229ffbdfcd6ff7f127546ea17;
reg [flogtanh_WDTH -1:0] Ifbb918c9c8ed9c0de0d1fd1e02eccd4d, I551b47851eee1b096612760b461e8207;
reg [flogtanh_WDTH -1:0] Ib230198837d881f6349f181cf4b3c4c8, I273b2b9c28034900d30631a61f1aecc7;
reg [flogtanh_WDTH -1:0] I1a07a0d5e3768a4ecf4c56f6698fef63, I641d4634620bb210a64564be02fa920f;
reg [flogtanh_WDTH -1:0] I55ff759485b4e816fac06d20ac5b2790, Ib0f8bb863f94f35f2c880323f8793565;
reg I317f33f435342ed704cee1defacfb4d6 ;
always @(posedge clk or negedge rstn)
if (!rstn) begin
 I148a2b6bf6253f900182125f4f086010 <= 'h0;
 I23d8325c203e2a9e4118ea94210effa0 <= 'h0;
 I9cdc23307c28dd846a7981b6a1b8552e <= 'h0;
 I2b9e2a2b9bea3cdd0c7b48f864254aa8 <= 'h0;
 I0da340314517b5042829528ed7621d8f <= 'h0;
 I4edefd1be2348543f0e11dbce5623271 <= 'h0;
 I8315a1e97dcb0458031c17b029afac99 <= 'h0;
 I2b91900229ffbdfcd6ff7f127546ea17 <= 'h0;
 I551b47851eee1b096612760b461e8207 <= 'h0;
 I273b2b9c28034900d30631a61f1aecc7 <= 'h0;
 I641d4634620bb210a64564be02fa920f <= 'h0;
 Ib0f8bb863f94f35f2c880323f8793565 <= 'h0;
 I317f33f435342ed704cee1defacfb4d6 <= 'h0;
end
else
begin
 I148a2b6bf6253f900182125f4f086010 <=  I5615abbd072d30da52163f16f1980957;
 I23d8325c203e2a9e4118ea94210effa0 <=  Ie7e694e2f86689b06efbd2eb66c5ffd8;
 I9cdc23307c28dd846a7981b6a1b8552e <=  Id0287bb263a65d5eea34cbd5be2cfe3d;
 I2b9e2a2b9bea3cdd0c7b48f864254aa8 <=  Ic223bac65f3241d30afc2e21178eebfc;
 I0da340314517b5042829528ed7621d8f <=  I22794d7d1503d8cf477ad8b189d53ace;
 I4edefd1be2348543f0e11dbce5623271 <=  I8ccd9901d0629218945ab24f6eea34a3;
 I8315a1e97dcb0458031c17b029afac99 <=  Ifdeb82639682ca4a87f76e40a181bf79;
 I2b91900229ffbdfcd6ff7f127546ea17 <=  Ib1879574e569ce9d6787132cc87e8de4;
 I551b47851eee1b096612760b461e8207 <=  Ifbb918c9c8ed9c0de0d1fd1e02eccd4d;
 I273b2b9c28034900d30631a61f1aecc7 <=  Ib230198837d881f6349f181cf4b3c4c8;
 I641d4634620bb210a64564be02fa920f <=  I1a07a0d5e3768a4ecf4c56f6698fef63;
 Ib0f8bb863f94f35f2c880323f8793565 <=  I55ff759485b4e816fac06d20ac5b2790;
 I317f33f435342ed704cee1defacfb4d6 <=  I5a0cb346d513664787453b72c079d980;
end
