 parameter fgallag_WDTH =  20 ;
 reg  [fgallag_WDTH -1 :0] fgallag_sel ;
 reg  ['h7ffff:0] [$clog2('h7000+1)-1:0] I2921115a104a4c6799b85673837b12992d6251292ee3f5f63bf7126c12eac61b ;
