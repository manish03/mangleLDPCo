`include "fgallag/GF2_LDPC_fgallag_0x00000_assign.sv.1"
`include "fgallag/GF2_LDPC_fgallag_0x00000_assign.sv.2"
