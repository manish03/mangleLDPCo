//#;; Ic23fa9996925b610710d93e28c59a3e2 I10df3d67626099df882920ba6552f16d I93762d802eed04b3e1c59d1d46b35248 Ic9f869114804f0a61ce9b03def9d71f5 I9fc5887c030f7a3e19821ebec457e719
/*I816842ff6f8526885b6ad2d49236bc84*/
////////////////////////////////////////////////////////////////////////////////
//# Copyright (c) 2018 Secantec
//# No Permission to modify and distribute this program
//# even if this copyright message remains unaltered.
//#
//# Author: Secantec 27 April, 2018
//# $Id: $//#
//# Revision History
//#       MM      17  April, 2018    Initial release
//#
////////////////////////////////////////////////////////////////////////////////

// /Ic1111bd512b29e821b120b86446026b8/Id67f249b90615ca158b1258712c3a9fc -Ibea2f3fe6ec7414cdf0bf233abba7ef0 *I66986ae1d2ec0253762b97e22f881595* *If4ed727b4ff4652b44f0b32f7198402e* ; If83a0aa1f9ca0f7dd5994445ba7d9e80 I21f66e7dd81ae29064c26b66d9b3e967.I288404204e3d452229308317344a285d -If83a0aa1f9ca0f7dd5994445ba7d9e80 Ic4c7fcc09295dba6fc1fd0469d7e92e1.1.sv > Ic4c7fcc09295dba6fc1fd0469d7e92e1.1.I21f66e7dd81ae29064c26b66d9b3e967.sv ; Id6bfe3ce1bf5714887f4ffbb7b94feab -I958fb7ed1fb6d4960d15ffd3254be634 -Ie1e1d3d40573127e9ee0480caf1283d6 -Ia823f97963868b5794f5a36e4dbe5dec Ic4c7fcc09295dba6fc1fd0469d7e92e1.1.I21f66e7dd81ae29064c26b66d9b3e967.sv -I2db95e8e1a9267b7a1188556b2013b33 Ic4c7fcc09295dba6fc1fd0469d7e92e1.1.I21f66e7dd81ae29064c26b66d9b3e967.sv.Idc1d71bbb5c4d2a5e936db79ef10c19f

 /*I816842ff6f8526885b6ad2d49236bc84*/

/* I0c35fcd8aa6b70a1e6a2f67174222bd1 Ifaf61c215f3a90fcc150ac387f759daf I54a78636e8c6bd0efb73150b779d5eb5 */

module  sntc_ldpc_decoder#(
// I67ec42122b652ab9b7e9a4810f9f0db0/I58d53a433022417c56e36facb426c2b8.sv
parameter MM   = 'h 000a8 ,
// parameter MM =  'h  000a8  , 
parameter NN   = 'h 000d0 ,
// parameter NN =  'h  000d0  , 
parameter cmax = 'h 00017 ,
// parameter cmax =  'h  00017  , 
parameter rmax = 'h 0000a ,
// parameter rmax =  'h  0000a  , 


parameter SUM_NN         = $clog2(NN+1), // 8 : I307afb7f348272492f3cca58ef2f95d8
parameter SUM_MM         = $clog2(MM+1), // 8 : If78618843e4df2223e60ec190987c019
parameter LEN            = MM,
parameter SUM_NN_WDTH    = $clog2(SUM_NN+2),
parameter SUM_MM_WDTH    = $clog2(SUM_MM+2),
`include "NR_2_0_4/sntc_LDPC_dec_param.sv"
parameter MAX_SUM_WDTH_LONG = MAX_SUM_WDTH +8 +1,
parameter SIGN_MAX_SUM_WDTH_LONG = MAX_SUM_WDTH_LONG - 2,
parameter SUM_LEN= 32
) (

input wire [NN-1:0]                  q0_0,
input wire [NN-1:0]                  q0_1,
output wire [NN-1:0]                 final_y_nr_dec,

input wire [MM-1:0]                  exp_syn,
input wire [MM-1:0]                  cur_syndrome,
input wire [31:0]                    percent_probability_int,


input wire  [SUM_LEN-1:0]            HamDist_sum_mm,
input wire  [SUM_LEN-1:0]            HamDist_loop,
input wire  [SUM_LEN-1:0]            HamDist_loop_max,
input wire  [SUM_LEN-1:0]            HamDist_loop_percentage,

output reg                           converged_loops_ended,
output reg                           converged_pass_fail,

output reg                           HamDist_cntr_inc_converged_valid,

input wire  [SUM_LEN-1:0]            HamDist_iir1,
input wire  [SUM_LEN-1:0]            HamDist_iir2,
input wire  [SUM_LEN-1:0]            HamDist_iir3,

input wire                           start_dec,
input wire                           iter_start_int,
output reg                           hamming_code_calc_out,
/* I0c35fcd8aa6b70a1e6a2f67174222bd1 Ifaf61c215f3a90fcc150ac387f759daf I3bc180bd00be2c60a3a5a68e0dd49503 */
input wire                           clr,
/* I0c35fcd8aa6b70a1e6a2f67174222bd1 I18c0d99dcef0c6b3cc1cadd623fdbf9f I3bc180bd00be2c60a3a5a68e0dd49503 */
input wire                           rstn,
input wire                           clk

);

wire [NN-1:0]           tmp_bit;
assign final_y_nr_dec = tmp_bit;
`ifdef ENCRYPT
`endif

reg [MAX_SUM_WDTH_LONG-1:0]                  Ifeb14203f4daf31c7701a6a742be57cc;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic188ebb37ff178022c61400613f4f3dc;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib581c19864deecf01268595049268b19;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3f80921fd94cff373648fa34fcadd4d2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I661d84af541e30828bcbd962d72baba3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I229f7430f590d86a323b48806beec48c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1c6928cccb4bf7ea7dfd74e425b9624d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I26fa0a5f87600d9535e8f83fa1a11136;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6eabc5c074fb1e2183a5f1ecee87a518;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id87360986474c9bfa5266a90b59a9a8b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0107769bbd7c239685b4818731334437;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id63daaeb52208682533b5f136480a29c;
reg [MAX_SUM_WDTH_LONG-1:0]                  If723180430080198d18a08d6775ab208;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1e9d5c2338b6f89e43c30c0ad71f675c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I44abc734d6acf92a8e8209186d7a1676;
reg [MAX_SUM_WDTH_LONG-1:0]                  I11cce7dd119eb0e3acafc12dbc6d3536;
reg [MAX_SUM_WDTH_LONG-1:0]                  I72aa55988d58c664f3291b5786fc8ceb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I934b111c08439d3797cb8928c7238f23;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie69528583db8155917ab3d32a446de04;
reg [MAX_SUM_WDTH_LONG-1:0]                  I508cb12fa71441b216fd7c1899d00e24;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib22b47d95b72871e74069fe80a191680;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic69c6ea6b4f360efae87611c00b00fdb;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id9451e945bd26b8dcb4cb83ab4ade73b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifccbe59b7ebe3f692f5b7e7564ca50ba;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iba4627d3d3ef91f168068ed128c04113;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifd7275bc534fe9da81b12b25ed218e91;
reg [MAX_SUM_WDTH_LONG-1:0]                  I39bef4d462b0a3f88ce1485a58d66da0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I01a99ac2a3f919f4fc1680edb11c576b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib95e457d5ae9fc89e197c249414abbcd;
reg [MAX_SUM_WDTH_LONG-1:0]                  I322b3879383d75c43c55535f01fdfdd6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2be28be47a38e9ca9d3b9167327d3d59;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1adc689464e0b81fa165eb17e71310fa;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2ee6154b613d0d86c2354604e93a9a57;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2bdc0908c3d365d25f8026263dc4a258;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia7479d4940b575cf918cb8421f041e44;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icf6c6fcfa42c48f16a1b30cd325c139f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3c5b1cddd608ad869e0182ad68bd0494;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ife8337f33629521c096d4dcfde96e879;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic4425ae997c479e05e12347a803213dd;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8afa93d48ae589bb90cc74897defe4de;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3a0518d0d382758ae579acd7e6cd634a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I56d0b4df55f7f4181a51f58187d399e4;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifd28c1cd286b7a483891bdd094b70db1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8ae9260d2a5dd6c2ed4b6157946e38d4;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iadf7734be049c645819d9d023b58c4dc;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie405c3459c9caf16c0a257a059a9fa96;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5f23af0d0853ea6de084ccf77702b78d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie76a46f18cbb52a93a4fad65462da3e8;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic5c99c42e9ebe5dded369ac78a1bedb5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0445dbe40692ef21353aacc7b4f7a4c9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4f2498bec0e96802b82f0419d97c527f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie3be0f770c8ddbdf301ae23881499e9d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icaf86e0abee612aa972388c0b6f90763;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3a4d175e3b015a17f7a49cc6bacbd12f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I478c4f13c05651605a2045bb5fd6b60d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id85473220f4909f9182711939cf6a978;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ide67911b52687d67ef0c25f2aadf14c5;
reg [MAX_SUM_WDTH_LONG-1:0]                  If77ecdb29d692c01752be0908c4f4392;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie9e7630af25f39a0e820181918edd029;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia188482ea4a2696f188f637912aa6f3b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0e1f07f30cfe36f189e9dcb4e713b5c8;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibd0c9231ee029200ca39013c839bc4ae;
reg [MAX_SUM_WDTH_LONG-1:0]                  I31cee5e2a93635987776b0ea477e6211;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0fed2eb07a75f701ff7b7ca9dbcddb81;
reg [MAX_SUM_WDTH_LONG-1:0]                  I84721f2bc5ae10db78d2e7e07cc28d94;
reg [MAX_SUM_WDTH_LONG-1:0]                  I96140f2ad00cb9a1249b5135ea251bc8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6c6d057e910da53aa47441566f95153e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I34fecbd6c558b25e7f8d08fb10b224f4;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iecbf70768fbaaab8da98eaa9a2b956ee;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8df49bd85a846a4c4c32af63798f3e0e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I71b8492d70b423e95938995c07395def;
reg [MAX_SUM_WDTH_LONG-1:0]                  I05be7b5c657867c4331ed3df72a1aec5;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iae469bcbba9598bb46aa7ccf9fa06a37;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id47eecb4e17f799da48d80451cb47b5d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie2e854376f4b6509ec41507401173269;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iedabb8b1ffd46b983fd74b9f6010dcca;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7b1401c3c2c389d9bf05658c88ff6b40;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib032a08190a75ceb242a9dc8272b4a02;
reg [MAX_SUM_WDTH_LONG-1:0]                  I88ee95aeb6c744eca0e127e8497b5dc9;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia870db84a0411e463b6e15f502323810;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5573e18ade3430ef3eff5e6d960e44eb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8105600a0847cabdb96310074840bdb7;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id6260fa8a9be077673e82344c736b1c4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7d6591184fd95d3f288f481734e85c02;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic052eadb342350c52d89e73d5fea80bb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I69c3d2866b040d67900eeb991b7c2981;
reg [MAX_SUM_WDTH_LONG-1:0]                  I98b8d024432fc54ebf2f15d99968f2e0;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ice61d34abe5e2a9593bfb911da54e959;
reg [MAX_SUM_WDTH_LONG-1:0]                  I98f54ab8454940141a484332f2a05369;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7dfe4eb1588a68b8a35dec39978d06eb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9d94ad2da06ac1fef4da7dcc56abffca;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ica59cc444ecf8f8700bf1ce16a254b89;
reg [MAX_SUM_WDTH_LONG-1:0]                  I51262e3abe460148e3c2d2b74989c2b8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0d69f1eb92a8b30d86ffbe0c153197f2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I560583680bb2f5a0b5ede42ceaafcf8b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5a48ea253b357c8e6441be01918bc57c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I389f83346ffaffe8186fb0074d71f43c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic3c81f609bf98f2ded891b55bacbd453;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie89c2a1b3943d12197bb972bd12595b0;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie38b3f5ad91f2c983d519c9b1200559c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic7be56919976a2d1088114c21c3c1ffb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1e5e2679a0e75104cc0be107ecadd01c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icb5dab0df062ab46bd3d1a73e85ef4c2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I903e174feff2be7109cdb19fa15a63ec;
reg [MAX_SUM_WDTH_LONG-1:0]                  I27a568cfc2df13cf689d366a25e5d05f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6893d09bc4fca46b4ad33c42d1950790;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia6688964078f1ea87b742352877aac45;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4ec84e063fb84d278ae90b84751b1bcc;
reg [MAX_SUM_WDTH_LONG-1:0]                  I180deab4fe0d03104cf2ee035f6a9b8c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I33998829023b087dbfa2e568d77291b3;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iff6cd034bb64d13c21910c11bd92266e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5bc68432bc0a9ea8cd024d7fc3d3fdc8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7c34057a77f2bdda93c422506959818d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib84e5271ffa3584148ce87dcf2a4f2a2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7ff7d3fd63fa67cd72d1591c1a373180;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib633998a5fd0df508b47ba9c2f7c390a;
reg [MAX_SUM_WDTH_LONG-1:0]                  If910e75bf10cf02a5b414cbb4fad1304;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie36cfd3519810d325d5cdc5150380fe0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I266697a6eca2b73a76fd375a0ad72a05;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6ac3755ff9de4d43d0493891b2a5758d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iba188abd7715fcbdad3b1f3d985c6fc3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5f0212d2ffe8f85614891882390bbc25;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic60c640562e3e45c89a1de78af509b6a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1e009fcbec9031954637f055cb9cfe01;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0456494b33e4ec852c123cb3003b9886;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia6caeb0fcc8e7486e4d55b72a0d499a5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2ed7c217fe3e21fcb27e04f68b95dd6b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I631e31da7dccd5b9311a4fa73e6a0227;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifda5780b42bf451a7ce834f17b3fdd20;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib152eea9af905931ab45c4f9d89fa50b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iadca92fd39d1fd6032feb8415ca5246f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I94118c50e80e5fed4294d16358d41579;
reg [MAX_SUM_WDTH_LONG-1:0]                  I613453382f19dd7eb9bdf51e945a33b0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1269d97f8ab4f5dddc002acf38b4a189;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ideafa683e6a3a38848fb8bee22eba11b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I89a793ddaf4887ddb8dbaaba13225d08;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie4226e7e17c7971f07aaf0cfaeae495a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2b4fe952791866aecbbbcf01257d527b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifbbfa268bd4c31c7eed45cd43fe6a405;
reg [MAX_SUM_WDTH_LONG-1:0]                  I797321bb9e3c2d7d3727af9a4cf5418b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib2d99d95f7a31e4745211c5ff96f851c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5eeb78b1511aa7b76765d82328323a4c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I692c0a91b415b400a3640e2d9a40edad;
reg [MAX_SUM_WDTH_LONG-1:0]                  I55f8232fcfcb929a35717f724f44eb4c;
reg [MAX_SUM_WDTH_LONG-1:0]                  If8c4dc70212e8873167e1cad8e8e5692;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7a7705607e93fca1cf1e7b1c92c4e3cc;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib2f75e91bf9e1d32a3f170fc85244139;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7e2e0ffb2b5622ba6e03a47755a9a1dc;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3606dc61f24567cb1ace443cea62a43b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5f50e835526833015a2087dbdb77686e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie402c9f793b7306323efb8fe23533250;
reg [MAX_SUM_WDTH_LONG-1:0]                  I98f32439ec64d796ebb157815b259aa2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I54652565023310e2eccfc4cb87c56b43;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id59ca1b1cff93a8544c54c6d4ee22b2f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I616b7a5987edbc001e0ae1b638f25a39;
reg [MAX_SUM_WDTH_LONG-1:0]                  I726538434626c5202d53d29faedddd56;
reg [MAX_SUM_WDTH_LONG-1:0]                  I06604bac478ee906b3fe8ff307cdf046;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8ea236c734f7b96620a37750134d3872;
reg [MAX_SUM_WDTH_LONG-1:0]                  I135dd8a85aca863db660f2ad4f80ca2e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I259d7244226dbcbd1d02df5ca164afdc;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8715d73b58270dfa33b903e9cfb50be8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I086375f289b769938edfc8b9b5146714;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7f60cb59895af6d314f5d0f401c80350;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icb82f8092f14511d62f7cbe821af9faf;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3e25e6e9de5ee9242a472ce957056762;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7e8df00362c29bd3924ecbe3dd1db23c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4c5f36517aaf872e7f05de2f7f76a6ce;
reg [MAX_SUM_WDTH_LONG-1:0]                  If1014cbbd6e267aaacbcf3c8ba33a98b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0e993e6f98616632f17835a2994f45e3;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iae4dfe3ede67923e8b740dd575b216b6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I281f996740b16568b9d29ca41a3fa50d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iccfddf46ea48242ca751b5d53f98d270;
reg [MAX_SUM_WDTH_LONG-1:0]                  I55bbb73d68871d9dbce4d590c029aeab;
reg [MAX_SUM_WDTH_LONG-1:0]                  I804705ac9a613b4107c8ceaac4127386;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ida491561008f4984480d1b0f09d2fa77;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8f40972503fbfdab92676a32f351dfe6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I624e237f248d292c0417ff85056857b0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8fc9ec077c7c6ce5e2660a4530a234ae;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic7c1fd79ba76dbb254c6183017f40b3e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3e3bf3c2155f584784863ae41cb73c7d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I546d683af76dc209a5205c6274abe908;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9cc24d95a0ddbe4145d144003778eebc;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7b4bb785489c5bb22c84d9778192fe44;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib9b96de1e217660c2ac9f7815249c6a2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifc6af7d7aeb7162d554b8604a44f3361;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2cc498e11d3d487d1e8319df8521ff6d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5b650c4c3291670b480a7f1095093dfb;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iae3d8158d13c8179719cbe12fdd7f9ab;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2f5f88cb5e5e4723bd8a83c5fa80cc4c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ieadf1b0e427ecddd261297ae4054a0bd;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic174b361182c98486e65b7f87b073274;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8dbe4e03db655e1f691254835fb58798;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7ba2f7201745258dbf224de087a25233;
reg [MAX_SUM_WDTH_LONG-1:0]                  I14b22818be28bc385f91920399012555;
reg [MAX_SUM_WDTH_LONG-1:0]                  I131a4bd335fc23ee10f7ccb1881ab9cd;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id2878a17128a23eee2272c7e39743bd3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I90cb3e06b42f25956b788a792eef371f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3701d2d2e74c43b3ae347902c0efff20;
reg [MAX_SUM_WDTH_LONG-1:0]                  I56302770a8d56932e7bb5dcff56c71e2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id6487b559b7ebad725aa43382f09bab3;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id3b8c058b3838c388eb5ddcb31dfc799;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib6ea830665d44628aef5041b2fa46328;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7ca8ce63dfb821d10304958bada71737;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia6181e1acc2ea46a85626a22983e2662;
reg [MAX_SUM_WDTH_LONG-1:0]                  I06ad44414b45d262f9542015d2dead8d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8b38fb1f95f036393933d07e0a60b875;
reg [MAX_SUM_WDTH_LONG-1:0]                  I833ef4acfed17e4699d65cbaa3e7dbd5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I33d76ad1185bbf80de5e8ff0ad52b15f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia77e3db939408af719e0a8555dcb68ed;
reg [MAX_SUM_WDTH_LONG-1:0]                  If2c522a90684b77b18f0058d1d2b14d8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I57ab4999187992eda55a82bf0f09b31f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I869e040de179572cdfd9373a4de8b31c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I21f7b5402ae8e8954d99931bd5108250;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3fb8890ee1f1cb30ecdf50d69e4ac0fa;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3627708869b47d460182bc5040092f9a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6b60e2478c009889776de20209929ee0;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifd88f0f0abd1c037434dc16e34550d2a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie6b559c2f0bd388d072b660341eebe31;
reg [MAX_SUM_WDTH_LONG-1:0]                  I27eec53da48406e7e1202345a0810e08;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia46aa3a3e6a01d4690dfe0e7f1eab548;
reg [MAX_SUM_WDTH_LONG-1:0]                  I682d42afaaf103550ce4fbdba6192c88;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idb7244908662bcd97fe8fe0db4b1abdc;
reg [MAX_SUM_WDTH_LONG-1:0]                  If225534847db8723768941c3819ed7c0;
reg [MAX_SUM_WDTH_LONG-1:0]                  If570b3495ea5b3f250cf4873f5dd0bb9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I43a91b2232a47d1f6731bafc15ced5db;
reg [MAX_SUM_WDTH_LONG-1:0]                  I50bbcccc40af5e9700b97e682953c8c9;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic54026604afd19b0c7c71ea1ac0f1c4e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5422f11a7e0b646dd4fa254602f91b34;
reg [MAX_SUM_WDTH_LONG-1:0]                  I218bd69f079aa21f0dda241ae6e387ad;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic5c34f86b03fffdcf723ff4116822e3f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iaaacca4d06ad0f202d839fd7674f1829;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2ebd72fb063702a7c36b4b546f4b94b8;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iecddac410bb2121da0df2d73c2d23cb8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6328eca7325eea20ccf30adf8b928edb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1aabc0c0b7b602297ad592ae48b23452;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ica13fd6daec896ddb0fa6be797edf6bb;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ida3aaf7237b1383cfe95eeccf3971a8e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I970c832cf68b5178f3d8111c9fed3b5a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idd2a8ed39edf6697b0988ee4eb4f2d95;
reg [MAX_SUM_WDTH_LONG-1:0]                  I65f78ccc122f96f97fee54955d370288;
reg [MAX_SUM_WDTH_LONG-1:0]                  I735c660d5232e03dd8fb129e2ca4b445;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5f77d7804a3e4adb641908be74f3ea19;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia04d6065987df3f007658614406cbc28;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9263e4ab78ca05f93ff921c4fd9ff787;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7aeddde5b60828ac7f8b6c2addaf220b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6f8f253cfb1fe1c2254e557f732a9b22;
reg [MAX_SUM_WDTH_LONG-1:0]                  I150c28296847348d69cce123f20656c3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3f247e74edd47e346d3bbb5dc3408844;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib94d38d19b3791fa2d1b42fdfde8435e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie0b33e2c1def11ccdaaae4ed2b042df6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I94865622898b2e481e86a244f7aa2759;
reg [MAX_SUM_WDTH_LONG-1:0]                  I39448514454c92ce93c3b0bc1d0e5d50;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1a4a432e735367f515ca747cef7d7d04;
reg [MAX_SUM_WDTH_LONG-1:0]                  I677e9047c3ede581db9512b4fe072ea9;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib3a2b744d8f38671a63da6f8f8f1a6a1;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ief6fbe6927f26b7a037f8e0bcb7751d8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I87716ad5a64592abb812ffe041ccc163;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie1e5c12afad8f2d8c2abef26473b7d9c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I71b259faefbea7ce8f47e0ffb556a0be;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic8f2ae80147ee27c548de195dfefa382;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2161b2ff3514dbdbb79d25da87eeec2b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I533eb0729cc85339e2fcd1847930adc9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I860a3c9fca8d240c68ce3825192353b0;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic68fd0a9ea4b641913aadb7fe011d8ab;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie4eb18c7e906c9a25c12e9980a9f61cb;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ica1f13759a67176573842e56bcdf09bd;
reg [MAX_SUM_WDTH_LONG-1:0]                  I20a24846a74af76fa4470d6350546a9a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifed30886099cbeb5da64d1d0696bb5de;
reg [MAX_SUM_WDTH_LONG-1:0]                  I90d40f6e9721a7d075512b8b81907453;
reg [MAX_SUM_WDTH_LONG-1:0]                  I317b34a0f6e16550b4a3e887cdd0c250;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifc4525a25f38affb399004b057d1318c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I39fa2bacef89a2f523f91b1e7f3cbe90;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icc93649a2050b9ded1e625be936b411f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id01272140c18ae29a8c75e493cf01268;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibcc30c960ae0f29c4efb1266c9e490ac;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4d981fbbadbaa97ef98429ac12ca6710;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3b2ffa79fd2227a24c6468a89f2bd989;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2a1672224d3a3c513f2f04bb4dc123e0;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib489a11dfdd8a2b3ad561c965b3d7d2a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I364afb3546858e133a2bb541798e7886;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifa51cf9f9d3d1b91c72387f5daf05c79;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9908671d65856b8714d43d83f0811a17;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifda20d77c574c8f13816620c56fff950;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3e3f06cade9b6c8ea10e45996449e405;
reg [MAX_SUM_WDTH_LONG-1:0]                  I03ce0915d3a170429959221b6c8cd16c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9525b42d4dc80c42608cfa0ea10b8b2d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9c2da511df8277b7e61cf8611d04dd32;
reg [MAX_SUM_WDTH_LONG-1:0]                  I94361c7eb9f16c4b20dfcdb7b8ad8cf3;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib8c628f3d97ffdf8a8b5db0fe90bbfa8;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idc043493a919ec50417594df96f4d669;
reg [MAX_SUM_WDTH_LONG-1:0]                  I42e0e42ae26723497a1da5e86e855499;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9e051ecfe79c36a913b15a0c7fe27f4d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id7e44a94fcaa2ca22ac9eb6756ecb830;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5479857f4f724aaea25ba124c9edb232;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie91db5e628b828dfaa8c1bd7d614d986;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id2ed64cae3cb1e0ada8e3fb4ebb2dc78;
reg [MAX_SUM_WDTH_LONG-1:0]                  I683ebfd7677d9e175d7a86479a5b42c6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I16b9849d3f2edd7f9ed7accb138d2c02;
reg [MAX_SUM_WDTH_LONG-1:0]                  I11090ba16ce17a70438618b474837c33;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibcfe38455aa7aa33ae950172fb915dc5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I845dd61995152e9d39cea7f0370b5a4d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic9d9832294a3707b4041b2c4d8f92615;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia3e4dff8c98b38b6aebec9094ed26421;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3ef9641c53e7aa6a588481b57b865aa3;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id69a54dc4854348a482f052c64a736ca;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie838f76c6fc041e4fa66441094ae477c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0f56c52253603ac01a22f3b942429262;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ice9f8149ed08f537da5e146b417085e0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I718f82404f82fe0e822ee20d33ad20a2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I71f6bd2fe34731aab306cfb89a3335ca;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6c86073aaa32b64a43d06eb1a2d9fba8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5dd57cfd0d7ce83fcbdb3f560ac713fb;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie0c8e27167e6ba97a83dd238086f45e6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I239498228bdcb1c2a8b2cbef48e850a6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6bb5e8ee16a2bc0c3b77c882cfb659e7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I82fc4233a3d2840670eb9b9adf6c9215;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ieef625ad664ddadc849be46d1c083748;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ieb08f6a94aa827632606608d014e26d3;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ice91b069200a91b2ad48fbf87bb2e766;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifdbb9947713ac574738236fcb5c6ae07;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9d4c7c85b4da5f7003ff05ed3a240a2e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia737ee8f2c01feba1db87fe3e1a2388c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia8f1616f8a65025446a5ab4cc1624f9b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5d8e065dba640832d9d8db3e4338fbb5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I29848deb21ad480cdf155d849dc7bd48;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3b3e36ffb1cff2c07bc9a61afdde10c1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1ae69988f89b200bd0e48f640211321c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2c8137e5ee04a1067858d7bb8d09d65b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7ddcc3c9f4d21aacc07d8eb285dee83e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I38eb22d29ad9f4192499980fc17898b4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I28f7cf50ea7ac81667ff1353e0e121bd;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib714941df0aaca40e7573e030d97b3f1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I09b7dd699ae0c4d34a7d1588efc90452;
reg [MAX_SUM_WDTH_LONG-1:0]                  I47bcab5b082a8ce6312244224c162d39;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic937101cc53e67403e56ac85011aa9ba;
reg [MAX_SUM_WDTH_LONG-1:0]                  I68ded74f52dbd02ceb1da62a79d619d2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib42b03d2f76b8939ff3183008b17a969;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iaa113fd5f1e0c51d9f47240fe81b5604;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4b99f00b1c2cdcee6bf4f1d2e8199ee4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I907bf413f65fad54303751c054687b29;
reg [MAX_SUM_WDTH_LONG-1:0]                  I01e153b020e1349eb66b47de581408df;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7b727f2e9454f90d4fa4ef2cf69ddf23;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8ca1a48206ed8f1dc7ca57d77d0331a2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6fc1f37134064dd7514b46ce7d27ceaa;
reg [MAX_SUM_WDTH_LONG-1:0]                  I40e8430f50206db37e500c22f461b0c7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7856585e0374651fc5f9921f69706a0b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I521128b7d945e025ded04037494c850a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I79b1967c2128c611ee4fe0d14bced1f4;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic24dbb1a30bb9a32c1992afcba90d4fb;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib8aeaf62789d1d7a5a23d7492ff551b2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I06cc903106b42e397fa7c4bc6c5edea4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9a8e8c3ce2c6323acee0877d445a2268;
reg [MAX_SUM_WDTH_LONG-1:0]                  I765dff22de01d419a6626919d23850f2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I701a3c05ad8e6ac5cea30b78707e77d1;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie9538b63a057a50371de2d17898d3ad7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I75fefd09122859510021931c16051262;
reg [MAX_SUM_WDTH_LONG-1:0]                  If93a5596528db9017b8783fa0cf1dbc2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2779af0ff280ea511af850df795d1fb6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I68016caaf170fbe2734c5b6aaf089894;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2eb84b0b6b12b9269bb791ae03e5094d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I169b0fac6d01a713986b636bf8dfc3fb;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie42cb87efb2b87d88eed6139132bb23e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iddb14d68b464d04fe9e0b4e62789601a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id2e2722999e300df1bc7ea89dbf5689d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie5b71f77beb734a6ab7f7be6c6f9c252;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2b7e1a65c52821f3f7e194a443b0117d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I59f9fa0b81ca88915c338ece1d1e08d5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8b31aa4edbc800c99628c5851cad8770;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4f27922ccb21b65dcfe2dc0fcc97cdf3;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id40d461c28ecc2017d9b7d2eadf5ea44;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idd7ae55ba748fb36e49684037212936d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4b8f58440e6848610f2e7e06efbc64fe;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib8da505d1572487e814e7b0682e6dfa9;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ica1d5cc8dc277e91787ec1bf0f2ed65c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idedb59a6fa2f6ad049f81ac652c645d8;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie5d481ac7a371e1fd3c48c5cf9649a67;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7d50b49718ab2007accda67ac77a65d0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9786bf468ba8540d7e75d762fc832709;
reg [MAX_SUM_WDTH_LONG-1:0]                  I27e0600689451a7475a36143f0eb1079;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib093fabefab0a1b46d2199c1c948abc8;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iba6724b61ecb74552b9bb3cab96480c6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9b53bbb22003297175c6c4655ef83c93;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0abb44bd896fbc695e880fee67fb0c42;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9df2a441fadba7dc49effc5eecf4b0e8;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifd714548110aa979e735cc6e13d3ef57;
reg [MAX_SUM_WDTH_LONG-1:0]                  I102372ac8a06119e5d827d83f172bbd2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ieeb6c7cdf1379ee3d2933d81bc812dbc;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5cad4cd564b0956b08f22cd42d594b01;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id682af5250edce8e3811d418ecf2dd10;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id685ced1c37d97c75b49b2f790dbabad;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1d02127e28fb2e9aaf352815627960e7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I219e400c87948e7b2bf715745a4b152c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibee34260749dc92b8523e83cd64d6a40;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3372567dacc350adf991928753209605;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie9a2a59c7b3571194198dca0c679c5f6;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibf50476ac553bceaedcb121b28093394;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie4b5a941feb385e88498a98e5f8ddc01;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5d20fcccde5844e36b83d7fd7034c413;
reg [MAX_SUM_WDTH_LONG-1:0]                  I30b2b34a0cecfdbdeecba5f286befccd;
reg [MAX_SUM_WDTH_LONG-1:0]                  I47e720341773b3a11f4c71b4e9644525;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8ce739ddc344cacb2de7f2c88a882170;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0251d8ecec82a24878ce494f0b417ce3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8b00260bb93e928e66e9d4aaeb0d9b55;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibeef795b2235c98439628da8d7c094e0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9c1ca916654bad308af37d040b486cf8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I61769f7c08a0b9cf78068455410b6bb2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I05749703a8a131453c563ed2264680a7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I77fe52c685b1075c294ac3c0a5b0d63a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4b76fe5f9863a41733b76decf9867d16;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia688029a35b4a62417906c9aa1cd7719;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2805bb16fd574a64de548b39a532cd8a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifaaab2c6f368b133936a7295eeb9b45d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ide6a696c06f17f455d56bb28cad98bd0;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifbe064ac0a5f4bbf6caae486064a983d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I39bce1f71ede4663c187ddfd6501eda1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I439ac39c831e0ca87a40f49e439ce24f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id0e769bee61ae0a90c167fab061f5965;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5c616021ebd98fc8e0fcf5b19732175c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I83e03af8657a4a237641a9da7922e502;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id3a6c8114a92efaf5f6c280f897bef71;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7565e071282ca6e77bb469afc522f1a2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I854d4e2867b459da2e2fc06c438e6077;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5d0dc5d40385ab67bc7f540f212b6a97;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3b334e8064cbfe97e70a0f4055496f04;
reg [MAX_SUM_WDTH_LONG-1:0]                  I548cac395730b8386670cc4c7a64319a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iff92d12470884efa033800c88e1983e3;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic6d9bbbfb7890540edd10aa5758b0c4b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3d167f5af41902dc0a6477d55cf0abfd;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7beb1f915a881a302f93c869d81417d1;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iaa7edba3767735cad1ec76479b5548b0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5fc389bbc1ce31f7b326da719dc576d4;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifaa7aff0fb2af9d3e04b2641b13cf884;
reg [MAX_SUM_WDTH_LONG-1:0]                  I922e6f05f7c6e0f6f0b1a5c9548df238;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia78b9e9a1faddb38b4a1472f5eea3939;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8c6bb234a1ca3deba637adf746672194;
reg [MAX_SUM_WDTH_LONG-1:0]                  I367d25430d8ec417123931f9534f3eba;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ide24ebd7423d4c4f43577b019f2e30e4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I38a19bd51c6ee4fcb38493d869b7808a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifc412122eab7560c9021a17d7f8700c4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0fe662c7d5cce9cf3cac56b6125852ff;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia5a56ed2c6b98e72002c6c5f946e7264;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6867bb41ee0a7f4c6ae0071e7975526d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia888ed8885f66084b777f66e25cef1e7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I74d3dc7b6116f47b27dbfd112d7afd5d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I248229aecef00b87a70ce88920e407f5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I13440021cb8441969d3242de4fc6a0b5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3d162a0ec918f220a7d5f4efdf89cb58;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id3c71879c307df1390bbc60c55a5f249;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1ca0372f60e48f2f803778c9017023c0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2e1fa8e49bf48184e6a669d18f5c8ced;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ieb9693d54f0808b0ba463fd3c316a80e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibc9c9339a0bcbc6addcce833051a8cd0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I63da03315d7e51fcacb0bc0298e506ed;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2c0a2ad9eef6e84c60d1a6503aa836db;
reg [MAX_SUM_WDTH_LONG-1:0]                  I918f5a12e96bb96941f019940f27a5be;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3b06c3a23b2068e8f45870524c4af870;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib4fb115f442ff544fa3d21b4e9d3f075;
reg [MAX_SUM_WDTH_LONG-1:0]                  I87d44c01b261e9c13add415e6b3cc5ba;
reg [MAX_SUM_WDTH_LONG-1:0]                  I387403482432a3196109484d1120d584;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifc15e0dd91741676f23cc20fc542ec14;
reg [MAX_SUM_WDTH_LONG-1:0]                  I619af17eaa4a56726d6ab322a74dd0a4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I50fdfffb4e2dbcf33282b3653f595ad0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7a67ed3bb370520d0d25ce407ab8cd8b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4e9786ec39d388cdce110c86bb436ae3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7629b35ca548190a81021a2c13d8919b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I47cb30eb341ae7ce99042a16cd109f26;
reg [MAX_SUM_WDTH_LONG-1:0]                  I004851d3828f135ebe4d2e6ab83936bf;
reg [MAX_SUM_WDTH_LONG-1:0]                  If004fa1c4e6bbe1f458c2d2a4f1f6e03;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0e2c382b2e62ed43b76697230e34b719;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7c9910ade59c54e170c4f10822b5aff4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I36dac27d10701db70fb2b5996a3f038f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I98939499dd98e583a4788cacc66c7fc4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I51d62ebd160eb0d073a7efb64d20079a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic530781e13180026815873e12550e405;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib3545a88d68631af1c94ca2cb1f379af;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iba43927cdbcb6a80953fced163686073;
reg [MAX_SUM_WDTH_LONG-1:0]                  I81ad7b044118734f4dc32a1a4e8eba31;
reg [MAX_SUM_WDTH_LONG-1:0]                  I29aefee3f95a7d2838ec5068515f69b0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5ad8c235d46349b6d310d0f175f84288;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib964c4dd0a0ce2553766251b73018699;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibc00920378e2427df2a63a47dc3eaded;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifd870cf74e7e3e5b348ad55af7242c27;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic5195bbaa69d95059cca6e152dc9f705;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic4ba744721cdd747affca302b2b926d4;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia01f20e0bcf35c2ee4963e9c392c1004;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id381e35622a3ac2c549a8c9b702ec020;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9f6f48fea88d1cd73ef2b24c7e819964;
reg [MAX_SUM_WDTH_LONG-1:0]                  If49e3943165e2782c928a7da86847145;
reg [MAX_SUM_WDTH_LONG-1:0]                  I847feea780cc8a06caea2d2ea79ad281;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie4d85aa4951d1a918d698c9e411b1ab2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7ef6f4aeda7fd6775839c068c681f9bc;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iff6a8d4bc8f5f37d0ccc2d41f469ca86;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0645e741da20a4957747188273a655b1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6bed9b6e8b499c11d719f869467d2322;
reg [MAX_SUM_WDTH_LONG-1:0]                  I71125dffdd2d37e44dbb46143c1e8d9a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id1db54a136ab42fe675fa77b2b7fd2de;
reg [MAX_SUM_WDTH_LONG-1:0]                  I50c166f958b22ce866cd40334918274c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia6ed9442d22d3228ce14749ffdacfab2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icd225144fd331b870847044b4d02bed0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I32e0c22a86e88cadc6a956c213ff992c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5e876482090ce6007c2a2f2101c24654;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1b0dcddcb3e0a398857f038d3a52e719;
reg [MAX_SUM_WDTH_LONG-1:0]                  I026ded06f56d9ca93f47fd85aec4f7ad;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8c6bcabb8814607901102aca5f820293;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iec596e94ec168a564bccbbaa7df833c9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I731089de22b5becf3621097ed7a81b7e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib514e01c261e43a725582a10596eed32;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifb3674681315fa8cf6739996b823a7aa;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic19a62cdecb2329370f7e11c48d3738d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2d5ef5bf9c28065a2a4ab718fbc8ba3e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib2f5691baa59adfbaad62f6ffc71fb05;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7c5f9c301a0bdbf642f7b3f33e9bfc66;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9bdfaca6112385deb86e24ad7e45bbaa;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7bde3bcef8556c1b1e4c7d2192196e00;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0e647bb8351cfe7828423e7099525585;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id13f3a39b334d8a80b7c8286b09bd1e1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I185b758fb3e50bcfb1464fe2ab593cfe;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie6443f42260e0a2983927d0940c82a06;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie25e944f9e3100c39b69bb38dffca177;
reg [MAX_SUM_WDTH_LONG-1:0]                  I43003b2ef41b34363169f004a6668a59;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8e77032a54376578b3d16799e30c97f7;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic385923d90d69cd387eb9fb5f62fd9ba;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4cd2a7f8f8ec378200b00d03e447ac92;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2f642acd0cb0bd30177bc0d65751ed99;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1b3c55aca0da232cf3f81d6d0914729f;
reg [MAX_SUM_WDTH_LONG-1:0]                  If1064670adff5b00cbf7809e2621cfd5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I34c76f1a126120c4474e750e9b51e034;
reg [MAX_SUM_WDTH_LONG-1:0]                  I72311a2c7557be2b6cb95b3bc6f511a5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0edb624c344787066a2267757052196b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I79ee4c7277f713aa710ae8cf7c470aa1;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia8443f199838742595ac114f35c00143;
reg [MAX_SUM_WDTH_LONG-1:0]                  I32bfef7a7ecaa533e3bf92fb560e657b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib25b8a538c9d64880e114bf4a80ca42e;
reg [MAX_SUM_WDTH_LONG-1:0]                  If4a6b6a8b44d2c55c93b111d20525ec6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I25f6a3d7bb869082e4dbbd0ee8574c95;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7d41f27ff64d549b7e5df6b172969d8a;
reg [MAX_SUM_WDTH_LONG-1:0]                  If96057023747a1538d9f06966af48bc2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie3a2d4d85d4e4ac011887cbd329bd9b7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I199e995390462e06853b1f5cdbd46e0a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3bc9fcec69ab6a1efb2d86e03804415c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iec6325d585ddd0a9f86bb5cd0229960d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9ee16e46a399d1445fcdf251757a5e43;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4be1ccfec148a522fbf5b8375245cbb3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I45cf986a60a429a68051f76beb8188fb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I074386ff6a3d8d644f4b2501c69f26c7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4e48461fcd58a133a09d856852887a4f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I83b378e5534c553b57beb22c5178a3ce;
reg [MAX_SUM_WDTH_LONG-1:0]                  I901714025da5b89ee929ea2859f3e6c7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I14f79d67f75af6a495d6eb2986210cda;
reg [MAX_SUM_WDTH_LONG-1:0]                  I976786b0539b07b056dad0f050eeb53f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iacd805413ec1eb001b3083554f187554;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8e1ad4f44dcac3e770dd862413b25a4e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3e61e09fcc81a0011a79f5c5ce77bc46;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iaf5caa6558f0a98b91fb72db734bbec4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6e6cbb7dba8eb3c02b5b4e4469e23cea;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7b37d3b1b23f09c6ac46a94cf2c4ead7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8b25822c33f7d506ef69216af3fdab44;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ief8b577d924f257ae5e1dd47009b0db2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I06fd642cbc8aa2f65197801d7459cfa2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie59366fcd6132a48f3e9be1bb5b600c6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I22202e6c3de9b06c04ce9514af28933e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I273c1e28c3ed897b7d0f6b36a3a8def9;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib991cdbb91133cb82e154c575e00a174;
reg [MAX_SUM_WDTH_LONG-1:0]                  I64b507fe58b933919d0766631985a74e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5590364df6874420e169aa444ab520b9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7c0376cbc3660f3d82a5da22806ef5e3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I43a9e393037fb4aa84741dca22648459;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3884d561185660e7e0f461b3487fdfd4;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibb4d8301d90c66fdfac92b3fbc53c019;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4b991f90354e3f74d105a64929a97d6f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibae217fa4b808e4accbeb8f4a9a976ab;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9534939768f7d2532ca4e6757dfafb72;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia8bd7a3594f7084a57e64da023bf784c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I090228a60e5919fa88d842b1638ee296;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3ce4b9d41f5472bf60ed2802a2ab10eb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8994d511d611a3c1b7a8122cd3d2825e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I93ec9bc6fbd056e7e52496546493e727;
reg [MAX_SUM_WDTH_LONG-1:0]                  I43d14ec8853bfd211aa6b887c7ebdd5a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2374b90dde1cf481baa40af31e1a43e3;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icd810cceba64ffbb087600155338911c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0cee595f488a909ade8a3b4c90dbb0c7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I33ddd4cdef0a0704f204f4fdb14fd859;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iba4c3d91d492b000ab1de7add9f171a9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0c87f78f08ac77246d7b3b8604dfd700;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2b4152aa4c51cc1c1ffabac78cea267c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I54745c58c61eba829e4717cd842d519d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie4c3dd5c191aff00a6d62006223c2b76;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9e278d7b6cccaa39163d0867427709ed;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie4c0ba9510f9b924999bb5f432137271;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3e5d8af6fed6b47aebf2eef7010afa8b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5bad544a17b384973d5672acbe0ac0d5;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie96538fd32c8f8d7a3144012d10b29a5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I231bfb8e19e1d9c4bbd29a0bd75c1ed3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I050a226112c903de442358e2d5be8274;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1ecf87e33de04d02db9e64590bcaffde;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4df410c6a7eea67fd73cc33c791e7aa0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I60c97bf58193f004e3fcfdbd6a03ce6e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id7e318f124e0534c8e0538f99616ed01;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib71065a3fe70d3ab5f05b0c393278631;
reg [MAX_SUM_WDTH_LONG-1:0]                  I66ba7e48a07f5fdfe16d23b0dc243514;
reg [MAX_SUM_WDTH_LONG-1:0]                  I984074a5c77445ad266463e20d77899e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I62e6e8be411f12cd5c4d63f1825521f3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I50bb40691aa09c42e0b64a076b50a971;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2f94d5aad80c081124e3efa3804af183;
reg [MAX_SUM_WDTH_LONG-1:0]                  I753bff437b6c563f5fddf19685405504;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7a91b23716bf81bea4956eafb467c96a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I21f2ec69bcc507756e2a5f85d3ead3e8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I17572136bb435e84505c016523a6ec88;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iddec4486996054e475499d370016a685;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9b0ac56afa21022e8bc69f5d20d17b66;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3d3edd06f8907f4369b825062348da87;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id9468cba18d4c67a84cb2b16d2cf495e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I72467ef10ecced8395a6870a39525787;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2bda0265c40a5cedc359dee75fb15b4c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9b74b672f55e7bf7560ba4dd2d0c79fd;
reg [MAX_SUM_WDTH_LONG-1:0]                  I318ebdf91ab8e83b80a880395879fc77;
reg [MAX_SUM_WDTH_LONG-1:0]                  I285b012d2fb5e2279a79cf8edca24ac8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8ac8dbc25a20c0c27e09240a5cd1bfd2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8faf911a7d1ea8b0abe54f6688068ca0;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id8c4e5d6318622bd8ec2974684f542b6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3dca974bf2d5631a47ebf8b945efab20;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8df19e0871c18890419c593410596b59;
reg [MAX_SUM_WDTH_LONG-1:0]                  I12141c45d147b058a9e392f3b7d7d06e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifb977d4c5bac50b9d7f2f814a500f0f2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia527c96e30b782f837bc6206961400e4;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id9a1f5bd846dc7d093ed9392722317be;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6adbdb64422a08be9bf9e538db97463b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic886ecf946cd5c297012444cb34980ab;
reg [MAX_SUM_WDTH_LONG-1:0]                  I958cdf5367c7b0bd58b70b763d3af8aa;
reg [MAX_SUM_WDTH_LONG-1:0]                  I37085a233f195dce1a76d05b0157fcac;
reg [MAX_SUM_WDTH_LONG-1:0]                  I91b7b8e8887b5dd9853297463c55b78d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia2812d1ba8ca6831a2f059eb23384b38;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6162978f0c57958ad0403246fb0530dd;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id176f2681568337762559e78cde29ba6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I508142e70fd04513977130556aa574ef;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia0c4e9942a4b08f69c2a027a712c9e39;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2afab673e4b803ffd888f187de47fa49;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2da299005fed6f2b710e25acd48ebe91;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7a56f81596920126a9ea2c9fb3a19285;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia1038e3b807e16a30f6f4564509ddd30;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic6252de2c819f2243476ddf82e22d137;
reg [MAX_SUM_WDTH_LONG-1:0]                  I25d94516522c19c0e53b5f52f4480216;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ieea8672b2f23711c6ba893de5c5d8bc2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4b96be53e3d059113bb74b27ffe30179;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3a4dbdf517b8f9c93b567f91870e6160;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic091d8daff9f609c53cb191ed6b6ddeb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4731ee7a0e08c69e2bd2a8bcea0838c2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2468caeaf9733c8bc6a485542b6b263f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1b6cbbcf01a65cd1c2f1e241f849c904;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6611d1fa58dd253fe6344a41584d7e22;
reg [MAX_SUM_WDTH_LONG-1:0]                  I663aee79f824c854f57c19e87207529b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8afb33eced17e8675a8e2bd90d16030b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I34ff7299c9d83affa4512b7da302c199;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idac55755226133905d3250273b1eccb8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I70ca6c9d0a5c99e0036479f7b5dd760a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4cd564459b8d65976195b2994e7d44f2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I835bb7345787eaadc41816858e0a71a1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2280162ee1c08ccc9f0c17d1ca0e3628;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3c7f6fdd0e9cc7426df76027912d1ccb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I28b3ba64175358f277427fd790a9228b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9ff512085174a7720705d0fb37c4ec34;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6c03138440f9bd0cb2cfe12abf619c10;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6a69cdf2bae1ea68c9be56dcc4e76a59;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib3709eb9dfc3a594d38ea5a0ef0cd444;
reg [MAX_SUM_WDTH_LONG-1:0]                  I855ddead34ac131137ba644afbfea2b7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I44cf5ba18d7d029df13f446f09191b2c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib1a463388daf270eb0ce698d7b5ded4b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6aa1e5acf0c2b01c94438bd1cff484c6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I74e4bb7530c02073f9b15a6389659d4b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia23629f3881e4119c36576f7da58ceaa;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6721b13abeddc76139bdc7380434cc2a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2f12d1fa0b815564cefafc28ceb3de82;
reg [MAX_SUM_WDTH_LONG-1:0]                  I84fba239c5705bcd92096e204cc9438c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib09ac099bcf61b09922b353403b29987;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4d46e4d50176768fda897949545e2125;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3c2b6da8e286d0a7b628ba1071f29424;
reg [MAX_SUM_WDTH_LONG-1:0]                  I57086cfab3b163c3911c3cf7bfb3141a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I550630b507ceec38b960ab2a86a57f1a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ice174debd5dc911fdf5d5756cff8d731;
reg [MAX_SUM_WDTH_LONG-1:0]                  I795c1c91cb6b7870b7efb07d67085be1;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie369670edc5b602d305904f3a4a4381f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I531b70d12349f3bc67e6a3ec53368d97;
reg [MAX_SUM_WDTH_LONG-1:0]                  I41f66f79339962ef42fab3b88e571170;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id8a109043bc922b718c203bd5d60a999;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5cbd2fad4d90bd77ba3d2448a37ac60f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic126109499ee1dc2787ab05b404e7ae2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id86a2869148e2885633d9e277f7041c3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1cd8ba53b876e2436901749e355f354b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifb7b585189db23efabfb522c9b45bede;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4e8ff51a6f70f8ca6a17a1dea8caf0a9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7763f0d28d8065d8c94ef8df96b2ab06;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic1a27480c9acc1684f3fed116d74cb5f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I115ba88588187c7115977e95bd26ee5a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0df7a888610865486aa1aaa2703dd041;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6e7f2bdd0c8231a3689893ef4877fdba;
reg [MAX_SUM_WDTH_LONG-1:0]                  If6448c72403a3d0bd904beac87f8aa96;
reg [MAX_SUM_WDTH_LONG-1:0]                  I546c513d5357ac1a6fe669888dfaf717;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iecf45496b391208d62e88544b5d2ca49;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib3e12c614471912d0b276cb9f0382b1b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib0fd0a839c85f3da5ae7b221f6e623d6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7187a2499e3319da90b6d6fc64411b46;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie045750c9289c899860823f90a306f3c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9b46582473bb4dd5541a35ac708486f4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1627b19e0ca42f9c264b626809fb37b7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I929796fe327ee9c8a05e6bb683ae5d7c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic9593f3fe23f258c2ab4ddcadaa8ca4c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib6638da8b69373c2026d3f5305825cde;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idc0085a6595a7de7e2bc87c789b7d935;
reg [MAX_SUM_WDTH_LONG-1:0]                  I28c26bf4cf9693d1807818b2ca7883ac;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id029b4c310acea870263d3715689e729;
reg [MAX_SUM_WDTH_LONG-1:0]                  I291fc4eef4b80d1020c96488b869727e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iec123ddb8d1e623d03d85a667c97ef31;
reg [MAX_SUM_WDTH_LONG-1:0]                  I53006ed50f6211439681aa7659647e35;
reg [MAX_SUM_WDTH_LONG-1:0]                  I89f0b0713e165a454e187fa51e89c642;
reg [MAX_SUM_WDTH_LONG-1:0]                  I47fe32973727237ae0cd4c306c7efbfb;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id812cf3919ed50a5e3897d129eeb4b8d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic3e0c7d71f13a56a9a63e158c7f2cfa8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2d65b5115be2a22ed1e29426be3f0d15;
reg [MAX_SUM_WDTH_LONG-1:0]                  If383f241447cbea4e18f4f79fcdbf144;
reg [MAX_SUM_WDTH_LONG-1:0]                  I47c8671569e2c5c2a21f27aff2d1f4b8;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia05354d3b4f61299d5897832639df2c2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iaf2144dab2167cd2629067e40bea3053;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9faec40665477e8b3237773d606af2f0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4c2b80e4bbbd4c5e8d0da28c5d0f681e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id231ab3133d4bed02aad7e5f560ee5f0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6300fbbd385ad9280c751076bc68d70c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I13616c8c7be221cf4d2c13ae87c38bed;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iea078843b3c5139a395997c54462850a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8793bc728a4d423fb96a88c83bb9746f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I654debf65019f2748e631a051f3b17ca;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2fb6af0f152232550a3cadd55656df20;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1e88b57c19a1ddfc1c1f0e168b60f814;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5144918fcd4ce1a061644240730fc52a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibaf7ab7333434b0d7e76e436ee40a406;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1821eb21cdf8208ff6c2f28d963f7bd6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1af14572832bd6d6b5890b8340b79ec7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I80471575b1d4b69ef073056f798394ea;
reg [MAX_SUM_WDTH_LONG-1:0]                  I652d3ed935b39f8fda8d84296456d633;
reg [MAX_SUM_WDTH_LONG-1:0]                  I890bf9b72cc3c71351547178d72796e5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5e33cad360aae934f418852541f5f2bd;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icc9d28b84fa91028ae96cc9b8bae7555;
reg [MAX_SUM_WDTH_LONG-1:0]                  If950e448e3cba7cc9aa7aff7718775f7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0b0d167c415f8c14594bd61907d46d80;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9adf8836419a1c85b146e5e36de68af5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9577d49a74520355e53a1818f479db0e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0f2bcdf124dff4219fd1a35ed1db7937;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie6e888d582ba9e600e91b119e2804642;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iae82e5de28b12f962bd7c5e221317ac2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iccfac3d489b4b110d6b6e005a5ba45d8;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia7b3cb9de8e18f41561c2a46dda8696a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I69a67481ca8fd01dc5400dbe887b4f83;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id0119672c8b017bce6fdba53d4dccf8b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1f36f045becec7f0528f4a935d3da2ff;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4aaef2f654ba03b1dc05719c81d5da69;
reg [MAX_SUM_WDTH_LONG-1:0]                  I530fe7720e3bcda35e940aa4973a7da4;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia6355e548635a4107a11c7952aa8b3d9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I03069dda9fa863172d8747408800eeba;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0bd950eee6abde9d1eaaabbe902fff5d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie7f36ee89f2b092555fbf8031d2347d9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I93caf487f67a2adce04a7b2cd7fff358;
reg [MAX_SUM_WDTH_LONG-1:0]                  I18af7980562b28c537be3bea8dc5252b;
reg [MAX_SUM_WDTH_LONG-1:0]                  If68a9cc5609ea7d87062bad2ebddb1a8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I22ec20f9396d28ed39c5fc4bf060c44a;
reg [MAX_SUM_WDTH_LONG-1:0]                  If201a7afedfd1c329b55048e6bbad629;
reg [MAX_SUM_WDTH_LONG-1:0]                  I105eac4e38f4661c7c7ca32161e42baa;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1f8936599ead5ce1cd85132e382533f1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5030734bfa54065cbef20c1350cd647d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I37eb148270af62adba8341c83411f9f2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ieccf25e3abd6bae7dcf08baf815f3439;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie4729048b95fede1806dbd006de01338;
reg [MAX_SUM_WDTH_LONG-1:0]                  I600c21fca7901299f8e95e8fa0ea0eb0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I02330d212434a6e8c303db2c3d36a3e5;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic4363dfd133124dd45ec2211499d0788;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id89498cf205e0cdef4886afd878c48f6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7c0bc779c09847e3beb0a139e8826511;
reg [MAX_SUM_WDTH_LONG-1:0]                  I547ae5055196f12eeeb36d69c325b84d;
reg [MAX_SUM_WDTH_LONG-1:0]                  If64db4386bf8f7d07292f14e3b313520;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4871ccbe2f182791243b7bdcc9b8e286;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibf51e537b992c4b4c0539dda9948f45c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I12fd829f22ba908180290432320a3660;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9f83063bdc3c352024f702cb9dc71ce8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8f967710d03870e026564db0df46d146;
reg [MAX_SUM_WDTH_LONG-1:0]                  I72127f6d422ec68dcd47126b87b3d3b1;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia347d80a70a49605c51d19bc2e696aef;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0b4a1b48d110b820d8d87f6e94d32988;
reg [MAX_SUM_WDTH_LONG-1:0]                  I730db85d3d11d8327c6d48b8b87a00a4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2e3aeede695007fabe0d6247a93ed403;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5c6a3ec08cb17d6646bb3e63411a9698;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8c5ea3dc59fdcdea1c5f503dde1e815f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7b5baeec7b11eca457dcd9d2b2b64ac5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I873c4dbe95220e40d7388870520261bd;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic4c7a9d491c560d7b6c410d8216f59bf;
reg [MAX_SUM_WDTH_LONG-1:0]                  I561fa67a9bfbedffcb04e7a4d6b76a64;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2151735079b41a7f8cbfe2b93f1b7470;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia55752d6c4f20378ff570a661ab31d9a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia69e34af60619fa04e8478e2d04768bb;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia13307be43e9155ed0333df62ccc8bf2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7f9984597d0e7bcda92f13fbb8805687;
reg [MAX_SUM_WDTH_LONG-1:0]                  I07b3d1451487a55fbbedda48b0cb6c73;
reg [MAX_SUM_WDTH_LONG-1:0]                  I342ef25fefdb6a326dac80d76052bbd9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9f8cf1a6cd0182fba35a49bd232f062a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id1414254ab35ee805c4010432eb24243;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie2e488a8589559deeec8598cf6726f1f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8db7cc6cb4bf55131bee6b00e76baf46;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9118ee5ff8c9ba9b125e5baa07bf52e0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I355aec2468fa96e2f32c8c324c48c5f5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I13b894057e2deae2c00787385de252a8;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic45ea6e09fd20a2285b7e6e2507910f4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7797a3ea5b97b514a797243cf9fe890a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I288b192ad6d04370df8084511c7f44ce;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3af78697aacc410108d0be7fd13c686b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4d589e9479ee494636d90a910e530863;
reg [MAX_SUM_WDTH_LONG-1:0]                  I871cb63247618a543b444aa3f888fffe;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib8fcb6e6569d34c67145861431ad5334;
reg [MAX_SUM_WDTH_LONG-1:0]                  I124404013f8fc6b302661900b9ad8ed8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5405b3c646988338f12191bb8cb02205;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8e413271c9d13748a1aa2d1a018ff28f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I371946ff4a809b62ceed2334a9656787;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4d799e93b4dfcabd69977ddb25634a69;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6d5be8ddd471c1ddf781949169bd9807;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1487f0027b7d16f4bc85bb00e537cbaf;
reg [MAX_SUM_WDTH_LONG-1:0]                  I499f6bbf3456d23378ff02b6f65a5ae4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1a5cdaa10022adf0ffbbc0f58b3e690a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0c81821914371a777679053e2aa5a55e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I98246759d003e9bc6676ceb2d093a06b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ief591e9d4759a4b1059574bb624e4ce6;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia3c2dfb3c4a45091be7cfecfad11f3ec;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie40648c85ed87c979a54dfc1f85d1cc8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I74cda651bcb24472a7697ba017f831a4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I36956634f94d6053aa455b29bc0b7a0f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id7ba55b14ac0f471142011dc2d57cc4b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I05a652e83a9b8c2c38de64de6a70f8bc;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5890643c88c4255a0e5efd45f8af3ee2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iaefa87388884b85eed690e9917bc9d5b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4f53e4955e9e506a7169ae810da5dde6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I98836c38732b8da439946aa5fcbbd963;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifc7c1ea337b122fb720767f1890f1a6a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8ff116e234a1007cc47989f3fdcf88d6;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id40d6f3a8dd09678b25b3e579dd5fb68;
reg [MAX_SUM_WDTH_LONG-1:0]                  I53dfee31709f8eca30897d6bf1618418;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7002830b0a5f40ba2a2fe7a00c7b6d58;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3ac389b6b81baf93095cc3e9e9c3d8ef;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3f377e8994959ef8182a08538e393d9a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ief52e91e9170809b980aa881bf76957a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I71bf29f3519e3238cec112ef97ce0579;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iebf813928bcad8ee3b6911057c59752b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iaa4bc2f51984f383479b597e6cd4c873;
reg [MAX_SUM_WDTH_LONG-1:0]                  I57ae0d331753595cd56d45a28cd5c790;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9066a5cf776f80ebf89bdac1f2edb4ac;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibd173152b9400b4c8011451d68b07e4c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7319203d7231bebb6d6e52422cce5ed2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idc21b018b7b6f2e0bc627e8968e06eda;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4e8309976fd6011d78728cef935dc3c1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I783423950d0e0229826b2249f5cfdf5c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5ed502118c175d5bdb4607973554a3a3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6b8fc6d29fb4549e3f191f913bccff9e;
reg [MAX_SUM_WDTH_LONG-1:0]                  If457f80b3d29b60b840f886fa928297c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idc98380b110c22495027a7cdb6f2029d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7e0f785ec7554540c9a4a413a3afa75f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ieb72df81e325eda4d80a237454fa9dbd;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id3662bbe1b5191995d1656045fe6b6a6;
reg [MAX_SUM_WDTH_LONG-1:0]                  If70e7ed8d4989cd75d37af1dc5d185ed;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idf922fab93bc2357ac1f66f73f3ead0b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifc99661bc592c2c43bae53db10c8d472;
reg [MAX_SUM_WDTH_LONG-1:0]                  I780371393ef898aa144c5bc36e74c654;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic8860cc8d323e5a4c68233109ed70512;
reg [MAX_SUM_WDTH_LONG-1:0]                  I79696cd10cffa4c0181a2089da6b3262;
reg [MAX_SUM_WDTH_LONG-1:0]                  I439288f09536ca87fa0feb5f6436716e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I073155ab0359a13b77f730653dcfc08d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I66c4beb8fe2d9f363c8e153a12f216ca;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1b44f781d81438654f69bb7fbdb94011;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib2a96d55b1f7bf9b89286de32e59fad3;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id68f1a0ec8ff80da3190fe517bd935e3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3028dabd706c9e5768eac56c66463955;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3704464d41956032b779eebe27511815;
reg [MAX_SUM_WDTH_LONG-1:0]                  I265f3da3571d2ddb786b98ba3959823b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie6756ee9631791940ffc6fddb223b4d0;
reg [MAX_SUM_WDTH_LONG-1:0]                  If8d81c152d863660081339144b37a052;
reg [MAX_SUM_WDTH_LONG-1:0]                  I085151dfc2e773a7a485f5ef1b7cd6bd;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie9cba6422546d378655d0ef98ef974fb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2654e83fff153df7760c341f59a23396;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iaddf6de71a6329eb536f54e3d18d43d6;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iee3eec7a9d7a3a5c22281545ec143e50;
reg [MAX_SUM_WDTH_LONG-1:0]                  I280ed7bf157554fcad915f0e7fa12653;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ied2b9ca07a6d498abada30fb0726df24;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0ca797b233dcdac8e390e1e41d99b196;
reg [MAX_SUM_WDTH_LONG-1:0]                  If95315702519e7a08386a870e599aab0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I150792edd72cc07cf8242d787cb52056;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1091064aef7d915ba8fb6cbded069102;
reg [MAX_SUM_WDTH_LONG-1:0]                  I186c13747ff5a1ee6e562ad9e5faabd9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I40685c7d2c8be12698f734ec6213b5b4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6fb8240f8c68b71cafe4c2c43ac7db33;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icc7775fe34c162006b93662530fd4944;
reg [MAX_SUM_WDTH_LONG-1:0]                  I166f5cab59c2a66117f2287d2b11c096;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2e6f1a5695ad23b8ca282b344832ee8e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie896986a747c1cd8ccad7117125c6e0d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I016ce894bebdaa7e56af9deb1ccfb3f5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0c829f14ef188ff7ae1417e28903f2b3;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iad2dd0815c1107160992e5070632f76c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3591d4f320f8401ef8ad8f92d2d89bf6;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iefaba2acd282081b9a0a98ed057ca85e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3816895f23a1381e42aaeb64dd158fda;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id4ef94eb8d5db8810bca4c9d669f0b7f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic9c34a36b2fde9649064680904ec9150;
reg [MAX_SUM_WDTH_LONG-1:0]                  I04e845e6a5ed71978b636593dd749b12;
reg [MAX_SUM_WDTH_LONG-1:0]                  If7eb75eccc5a6384c80d99b64d534fca;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0b2760b437be2cb79382f8d6a7b8969e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib788a897a1d1b86b2c16caade11846ee;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1b0fdaeebe5fee6fbb2e13aac5e233a1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6a5fec9dad124f6d8c5574bcc2643ede;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iee872d17e4a28075be0ad7086c3acc91;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3936f324b08bea1bc5f8bcd12437b161;
reg [MAX_SUM_WDTH_LONG-1:0]                  I87656ddd4ef8f1ae36c7566d5e7892d8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1a59337d4da3e3ad1a738a9c3b56ef8c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I865cd0535644db7f17db1180c85f1744;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic3e3b4cba05d80c0ceaa6e25a906a602;
reg [MAX_SUM_WDTH_LONG-1:0]                  I71d46741fa94df65e1bdf6abff53d2ba;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ife0830e12b8bbb5aa0b8c2c0e4191e59;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic223d7941250d739ce9bb0ae5013646e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I95eaa4ac5199ebbb06f780d1376062ec;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1ef9b548b943a1f2012b91c7e0b445f2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib40ccfdb9ea28f333a7cc67f2446c923;
reg [MAX_SUM_WDTH_LONG-1:0]                  I88b6d7894d82ff394e89c7471c80dd5b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I507515355429e697cd5496809aa03cfb;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia5fc7e1f991f30042b848888a546534b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6bcc3a323e67f95eb4bf28a0704d3c50;
reg [MAX_SUM_WDTH_LONG-1:0]                  If699df4c8261ebce5c5d1aebe062cd61;
reg [MAX_SUM_WDTH_LONG-1:0]                  I55e3a2566ef3ac257021a294376be634;
reg [MAX_SUM_WDTH_LONG-1:0]                  I19338369553e96bb2476d80fe84dec3e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I40f10dc3289ea8a59f593f62066aaff8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9844ff02042cbc04dd5f4179908bbb2d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ieeabde5600d81208346ebd50d4a95d83;
reg [MAX_SUM_WDTH_LONG-1:0]                  I89cc6a060b714985b24f724adc782e7b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibb9220dcdd6d7fc2b6d6ca5f4cc93a8b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I39d94ce7fbe37a74404e0043060441ed;
reg [MAX_SUM_WDTH_LONG-1:0]                  I05a3aebc90966144a6809e460d6ceda1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0a1c9a8d59dbcffd6847f3a65107c407;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7e3150622eb318e94f99b36016ac7d2f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2328556c467a9e639f2b6ba1d0cb99b7;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifb146b2073d447377a1b21fe21baa4da;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5c9d75d6431d69db1abe412e591000a7;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifa5048ac43025e9cdf3f3436c37bb835;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8dc3dcdefc85b6ff8ecfa09cfc7e69fa;
reg [MAX_SUM_WDTH_LONG-1:0]                  I837ba4049e4973924e51d642f7f481ad;
reg [MAX_SUM_WDTH_LONG-1:0]                  I69f6c909ea6b207c200b154e00e13a05;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2910e5e74ca008b7e5502d787cb88a6d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id365c9f8f7f97c777bd5da0ce9490511;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia24816d601e29172628cad0c364b47e9;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idf0206d2ad2bdef7db1d30a2d715cc6a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8f99af880f329241cfc9616ff9859091;
reg [MAX_SUM_WDTH_LONG-1:0]                  I07d1c54431eed887554a136f15f86d22;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iea7c2970a7d80c55c1a6d6933c6c81c9;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic16809a3c82787ed88819fc9e9613f85;
reg [MAX_SUM_WDTH_LONG-1:0]                  I75a12697a4ee6de46fc098b0f02b8349;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1613ae89442495e703a52e65b8a0bf9f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I623d1f0b6829caf5dc0f0eab0ca47f74;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6089da825af433e847c0b1bb9ff7d373;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ieabf207f10f7df1e9059f1e953d7b399;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6aa7fccf4e225fa70063fd24dab74e6b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1399b55530e343bd85606e7c7529d453;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibe2a5f680405f233256b6fd806b72ae5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I39ee898ed8a8af64552e1aa145437310;
reg [MAX_SUM_WDTH_LONG-1:0]                  I662d408ffd8fb9f249e531a167161429;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0af241f9f65af3bff2bb0d69977bb0c6;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie95b8a5c2da6c0877d49c646c194f5b7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9de68705b5430023d2eb5554370bb188;
reg [MAX_SUM_WDTH_LONG-1:0]                  If940f33461f5e297e158db54f6aad610;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icdf7ba01c4813abe3cfa760f2d8d5c84;
reg [MAX_SUM_WDTH_LONG-1:0]                  I54aa9d4c6333d94970eae97aeb3603fa;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia6b995eb6bbaad8a638c80d587d45ab9;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib82fc62720e6346e1c05cc33d596447e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I75c2987dcebc9cdca578aeebec96fccc;
reg [MAX_SUM_WDTH_LONG-1:0]                  I24873624848b61f313865e10e77e35c6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6fab90e9a0f606d7c26346c89c6f1d47;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icc3915d8325c22fc172f731553798fef;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iab2f70a1d3093b3194e9047a8fe8e487;
reg [MAX_SUM_WDTH_LONG-1:0]                  I93b9837e63103431a0fdaf319a465c90;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic84b6224be8eb8eefc9ad9bcc2280291;
reg [MAX_SUM_WDTH_LONG-1:0]                  I91237af3aa2af551dbbc626bb701215e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I64a0e60fdcc93d84606774196b2b7598;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib254d9701567f642d3586641edf85128;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iaa6a4f3826d87e43dd3213dc5083184b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I25c50067a62d2b3599d15f12f89d384e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I94fd5b790a9dceab1b4b3f1b5e30a0d9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I238be7f0e4a209a6b4201a024c8aed82;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9c8c1d22021bbe798b1863ae1dfc3965;
reg [MAX_SUM_WDTH_LONG-1:0]                  I233f5ddadd45c0df2108ea6c1d634f3c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I870366e9c3b29c1683a7528f4b5d5329;
reg [MAX_SUM_WDTH_LONG-1:0]                  I87a320ddaa1478146ff6e519dc65c40a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I066db3b79f8b4581f96567d943a7e7db;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibf03d6940c0a38bef038a28b6a7b625d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iabd6f58c4760c939dfd58e4f426bcab9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I90942470e2057e50ce4f5745ed68b81c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia3505661cb9b7eacbd47774346d12f5b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I77fbc3f3b65962b610e39f4b085ecb7e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4e7245fc882e3e284d8c152c8998b028;
reg [MAX_SUM_WDTH_LONG-1:0]                  I701845efaf1b02aefa381d4f6b45c401;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibe962754759204890883a6de0993a64b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id446ddfd713c6e1592c562cfb123ea8b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id2ef1e193163adc702763541f37fec4d;
reg [MAX_SUM_WDTH_LONG-1:0]                  If4f752779d27392e7536565d425bce25;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8a925721cf106d4e6ca1f69bbc2f53d4;
reg [MAX_SUM_WDTH_LONG-1:0]                  If112169057d6293326a56443ac3cf517;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib97671e4daa1b606aa01c5e8f753a9e8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I78f727f8d85b5d7f0ffa57f02538f939;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icdd0962fd06355a7dcbb491543eb9cb6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I01ec629f60c17c2251f977205234cd44;
reg [MAX_SUM_WDTH_LONG-1:0]                  I003f9dc1b83f386f070b0a2e8c7ce4f4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I23f774adb64807c0edaa9941c75651b6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I66e8ad34c764833f038cff700a237fcb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2361ef4fd70e4c05b25289d0845564c4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I614bddda696787a552e28cfaa81a3aa3;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic3067b434ca17be7bad595e1f9b822c5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I38c22e6b7c066be10ec1f8929dbf88f9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3546ddbae9c9db4517802db56cee35f0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I245816ec4a0392af2cfa4b44a4e93610;
reg [MAX_SUM_WDTH_LONG-1:0]                  I35e91092ed503831ed818f36a1ce1537;
reg [MAX_SUM_WDTH_LONG-1:0]                  I83253182662d56779685c9742f55789f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I973f185cf29e13193abf0108d4faa9d1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I963a4391dba3d12756b89dda1e962c3f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iee58b0442a6cccf0990ebb551b47fa92;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie959690f46f82cbb15ae0cee69f3135f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2cb3207a5c1b25386ac7eb532955f260;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic475c578935fa69db2b1c834539750af;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icd4f07bc30c66f7f5b431ed97e7ac7b6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4f9bc0f2aeafb89fbaa0d0af7dbda06a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifec6f3a1e10144acb320d5d502ed1ea3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I393fa73117dcbf1fb1b74ea1fc7e6c99;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic87bff64a597e6d02583041b552328ee;
reg [MAX_SUM_WDTH_LONG-1:0]                  I95836c571386b3b6de07c9195932fe22;
reg [MAX_SUM_WDTH_LONG-1:0]                  I489f21ef8243ef8caa1c29f034c3e2ac;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6dd6f9abc962974c292d22f17a21a936;
reg [MAX_SUM_WDTH_LONG-1:0]                  I773901563077961acada85962209d68a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9f9e6bc8d2cc6e41813d42ffcd5cff01;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifbd176fe3e78bc2dc2e0e77ba3ccd2d0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2ba75ccf97b5caf5aa676a9e3c42a366;
reg [MAX_SUM_WDTH_LONG-1:0]                  I53f68a4cb81c71ee7bd6f61171b7478d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I006699f0e016e7022b2706751965c42c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7568ec59f1359bedce86dbc6af50df71;
reg [MAX_SUM_WDTH_LONG-1:0]                  I66d5992f4f39337782cfbbb9fec3b2c8;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id2bf82d6bf0a201f80a58357038a0992;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie5f503c91ddf6eff2b9645e6e3c22b2e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I22442354ca2b77306f25839ce6124699;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ieb7e6a2425e93a2b96a94f0e2c4442c3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I71a5c2876a07d8edd001ef2d108e59c1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4a0483f2d2585cd44fe35191d7cd88b1;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iaf333aa6b135927cf1ad1f76298ccd63;
reg [MAX_SUM_WDTH_LONG-1:0]                  I00e8b3cde14889fcb0b40dc5582a58f9;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia71cfd8cf9bea4e600ea204e41271c7d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib53dbb62231f729a278d2afa3acffdbf;
reg [MAX_SUM_WDTH_LONG-1:0]                  I164b032929ac2b8cf1a6672859639a30;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5503d6011d58dfa4e1ec524eb1875c7d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2ef0447f5c64fd5c65e23c16069a62ef;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id86fbda00d923c29c99b4a9fe52d513a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ide7008ee7f1fba156dc6145b3505e553;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3ba6e9f7d7fa98ad776299f8cd8a8363;
reg [MAX_SUM_WDTH_LONG-1:0]                  I129a7ced6bc6f48f20fa552e2519925c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I67b512efbaf9c063a4ac75cb97a8abdb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I67123cf825352e52cf0158060ad69a13;
reg [MAX_SUM_WDTH_LONG-1:0]                  If5f5eecf512463544c8b2419c0a58779;
reg [MAX_SUM_WDTH_LONG-1:0]                  I09923d784a9f9625a37221f639537941;
reg [MAX_SUM_WDTH_LONG-1:0]                  I81cdc8b54bc7f98798713985e8f4553e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5947be93fdb18bf0ad341fb826c9e6d7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I35bb2eb0cb589f694001ba1509cbf7f8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I08621ee033cd49702ad08af4d31eb999;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3bf8f19c98c78f8e1c315e75a533bb1c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id5eca60b22d3835119571fe4b1a03479;
reg [MAX_SUM_WDTH_LONG-1:0]                  I71cbdcd6e3a873851e9084bc9dcd99bd;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7267ba2b9cb511a48a3a7044e854f7da;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iebad2e3d84bae3d4807badae823aec52;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5893fa21ec8bbdcea9677cc12fc4057a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I054f07cdf6a44100034c7e2fb438055f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I564896fe01ec799a0fbe790473753559;
reg [MAX_SUM_WDTH_LONG-1:0]                  If3b82307d1ad78e262f76ba9b711e1a6;
reg [MAX_SUM_WDTH_LONG-1:0]                  If279ab7c515c4039c8272b913c2fa107;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0f40c8301521c136b3ede2cc9e8352a3;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib61705ff5820f531eb17c40ed05f6ec3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3615a34cbf1646a7cd0f1da43d62faa5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I50149e5de41ca2998c4e8cc4b19e166b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0bbd697ad8d3877570ab9e200e66164a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id40cac3272643f3f91b73c6aa1740f3b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I298f7389a7fd8e927b7e3354f0d32344;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic63eee2d700493c41ee2d186ff7111b9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9960d39fce3c5b9945965dedac46dfed;
reg [MAX_SUM_WDTH_LONG-1:0]                  I51de42598e0df4a76cf7b02c61ae9550;
reg [MAX_SUM_WDTH_LONG-1:0]                  I02f48e93599dc91bb24a144a0ef1a933;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia89a1a58f6327ee3c105cae860942171;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7e31af1959a0374af6c2767e4837c566;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib149a5872e31cd5df77b66298b4aad12;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8d18e2ecaf2bda4a0ba47d9782e9917a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iaa16c14572ad0442eb3c58a97bef5ada;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id0a13655f967dfd3000b8dcf4a57f555;
reg [MAX_SUM_WDTH_LONG-1:0]                  I88d5d48e05b1c9a6d8060f58917e3834;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibf384c0b998b5a5f7808c54292c6b844;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4269e18c2df4d39c683ffb7d01a08322;
reg [MAX_SUM_WDTH_LONG-1:0]                  I58b8202ae510e96b4f6ae334f3b282c6;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia29017fa9327fdaa7c10b2797f8aa6ec;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icbc75d6e4d0bcc42cdf813529b017e0e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia142ac799256541fe33f898a6a31dd71;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6fa1835a8e7f8ea435c4515b1c059cc9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4c039794243933a9bb7ad6db7eda6a87;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id3984a3dd1009c9c76347b9843f27b25;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0debb3ed4f9540c162cd525588e0ae3f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id5fd757abdc0b2e1b1d4c5dab96ee08a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I681eed68ee814fb18fd794207d9266e1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I98ab1b82b2991b4cb3bec530711bdc43;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic260784b8910f5a0483afee9b68efb31;
reg [MAX_SUM_WDTH_LONG-1:0]                  I610d0ed6f55a4906aac1be5823358392;
reg [MAX_SUM_WDTH_LONG-1:0]                  I22cd2d30a7684002cacca4deae4c95a0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2ed0ad73f73f9f4e1b7ec38af320ee4d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I136b4136d582f9fad21f90297cfafea3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3dfc4dd447cd1f4e40506f516c106861;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id8d6be9677d3b0ceca26b3b671757c2c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idfeea354b3f9ca8c671851fd90f4e1bc;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6a93f928c104ea211dcc8a461506327d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I415d8306edb869fc838eb518aad75168;
reg [MAX_SUM_WDTH_LONG-1:0]                  I240da147648bec33195a5f5c273fc6f4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1dc6b2aef1bb326c3d5c19f97a2e1d4f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I55494d0e8454e3cbb4158559e0d29984;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie2f47a06ca4b6d5823cbbe099f5de0f0;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ied3cc579b3cf126081acf8e1117007cf;
reg [MAX_SUM_WDTH_LONG-1:0]                  I55b7a58384e50ade254c3c8934c290f6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I76140bdc374dd6031097575fd231b468;
reg [MAX_SUM_WDTH_LONG-1:0]                  I53bf5dca5911aec50866be5a720d4aa2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I650345d21e5c2e7a9bf1810630161089;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie57f78d4c002e69e0e92b25bad752d3f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie852635f073dc918e7b1075ffad46f24;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2ac511a908c9973254672fd38cabccd3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9ec80c14eb5f0f305e1a9e6107a6001e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8f06d78dd2e6be736f4e4f41fadf130d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I80ba56447ab19b33610c23105b0b1637;
reg [MAX_SUM_WDTH_LONG-1:0]                  I65450e396e33720967b7a6271e3a70e1;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib9132d9fa7180c3fcbacb7c570d6b0f2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I876c6361d2164d03cad2ffc8bf920ac0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I01621f113f636a9caf9b5ca0bb20ef77;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id3b8e1157a3e9eea4d210f466740f673;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3eeddb549c6e1f07469c0e0dca68be92;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6973de59fb6014d7c4bf5b982cddc4d8;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibe664dd203ed4162abcd36eb8d57bfa6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I26cb99c4cc37be5f52dfeeca60d5d102;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia66176893fe306ecfb415d948c50486d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie9835b1d512d9c9c4f2801956fbf13cb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8bd4210dcbfc1956381b460fd9ef789b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I89057e4e979b903ae1f10f9dd2f196fe;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1ba6328ea9cb7cebcce47d5407d0eae7;
reg [MAX_SUM_WDTH_LONG-1:0]                  If1299e6b34cd1f2239d64ade23f33f01;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9e79c17bd782bb7981b4a3623baf96a1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3f106ef1876021bb3cc5866d2b5698f4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7c6f64d73ff9c6e7f2ed69713e056a2b;
reg [MAX_SUM_WDTH_LONG-1:0]                  If6cb9fec3dc380f1c4894bccfa35b33c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I00b962a9bf04b62244591051d2dfdbbd;
reg [MAX_SUM_WDTH_LONG-1:0]                  I313980f8406e9f26d5eaa53270a23b9e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3a660b57588325989319701026f658e6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I792b5aea212da69a9c18f5723e820432;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibae27cccf3f64e8653c1e244e940e421;
reg [MAX_SUM_WDTH_LONG-1:0]                  I98f245ec9b667dc065c9494c00ecdf88;
reg [MAX_SUM_WDTH_LONG-1:0]                  I27b89a5001312b2aa48fe385d8a52063;
reg [MAX_SUM_WDTH_LONG-1:0]                  I15254b39b6e136520a9497d8684f9d94;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic6a7476db711a812d146331c562ca7c9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6c8312a9d655f143a0b65d91907ce533;
reg [MAX_SUM_WDTH_LONG-1:0]                  I01ca07fe91b5f1edf87300b3583e77c5;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie6df2f89b05947f6be3b64e3b4f23df3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6da707fd74249175d1f68dccb66390c0;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia71232b0b468b729fa1262957cbe9faa;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0ae62aae426b75b06d95c46baf33f08e;
reg [MAX_SUM_WDTH_LONG-1:0]                  If75d8d882c6afc3df62096486b8e5b80;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iec512b5870f295a50921e7e0289a7d35;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7ed551b891500784c827992eb53f9ef9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3aac84acd9d78070472b1cbc745c80a7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5b5a24fd7116acd8ad2161513848c6a2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibbb900f56de318bf6e65b49791835ef4;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id7055f4e578533dbd25d0505f8e47f34;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2c2ac1e722fba72c759f1d37b88a9a10;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9c78f3a2aa3986718caf8e70d4d939d4;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ida0a18f1b79aff4ddf0e8f7e27794674;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2def789e23f8ea0edee6f58200144096;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9f2029db42c5a968b370587c958c8929;
reg [MAX_SUM_WDTH_LONG-1:0]                  I319c2cb3a815a6347511f0c398876a3c;
reg [MAX_SUM_WDTH_LONG-1:0]                  If5755f4f61a89d91a91188c17ff5dc5a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0603434655e30a66d4e00b2bc2c878c0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4419d97c3174ee4610eb6ee9c06cb256;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia6f16190b83b661f68a7a217bb356bdc;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia964f83676273055e20a2f63c8fffa0d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I68fc61dbee0900bd66be7c7f5aaf8825;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iab4fbc811e87df1d1f5821ea732b6a93;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4ddd7ecf84b4ee4a4b6290f3d362f190;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4fbefbb10724b0844c95e85495d4a87f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8e60b67eb6a187737de2717ebb95cf6c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I717217d0b5a526f04c7f5ab0835dd5c7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7e17264500cb48d228c20542c40169cb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I235937b643e8f2848116dc76c43f47a7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6bddfc7b277ff042899fb2acd5625c5e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7481f17d659cce5b4c72a68a9f6be67f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6daafbc7b14e2736b2a4e29c5f6fc5ff;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5715c21c80992a61bff8aabc3f80415b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I29df797d4c3ebd64fb088660bf89e922;
reg [MAX_SUM_WDTH_LONG-1:0]                  I434e3216a615eb46be5c26ef914b9cd2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9418cc6766916bf1afc1f8a01feaad4e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I918326ac0a744d234d74e2c08cf41eb4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I90e1a5b43e93c02512a76c5cab15c5ad;
reg [MAX_SUM_WDTH_LONG-1:0]                  I966706d314f4c0a7ec842dd699d34926;
reg [MAX_SUM_WDTH_LONG-1:0]                  I26977fe4cdb2f9714fae2f12ca4a809b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5a7d246d88ef12e999f4bdee40e5a585;
reg [MAX_SUM_WDTH_LONG-1:0]                  I59775b68e199902c38d62e28cff01393;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic2dfaf65c4e17a8dcd55f766c314d6ef;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9470ef82dad13754d8d061b5fd00a667;
reg [MAX_SUM_WDTH_LONG-1:0]                  I151831ba6bd0e162275c84815e3c0f12;
reg [MAX_SUM_WDTH_LONG-1:0]                  I62eb7a176351be84d086ce3c463214e8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5a8f1675234ebed14d719344b530bbd7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I106eb0d8f9ea92cda7bec4fe4aed6409;
reg [MAX_SUM_WDTH_LONG-1:0]                  I95dce76a8d0e729d40fb3f573cfc06ad;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id0c12bc1a2139e57ea40c3254f30de7b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6c26c7918254426c18f2e747c91438c5;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib809a6099992799ce0235f22ce798c9a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0414ead2472e42da8a271cb0bd1debf4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1a9be3897e044e9b24ac330ef3a20419;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic6a6f5090470a76ddb7315c022ddc104;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6e87b3400b7ddab94faf11c3910fa534;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2a00ee56a5aa639f45eb3b1bdcffe81c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I51e0ff0f52ca609663781545174b763d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibceb2b824cd4bc10bb06ee8adc693bd1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5c523df1fb2161ab4efd1c9b3e6b7aef;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia8b9f373fe68ac4cbca35e04376e3cca;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia307e5901694783f7761cdf724b767d0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5d1a89e85f6609b469e73e15aeffcbc4;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia47164e8ba831b85e696e30ff59ceab1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I677fe06bad241bc8dd6a65a97f6db520;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic217af0cb9728801034fdcb273a577fc;
reg [MAX_SUM_WDTH_LONG-1:0]                  If3c0f892fd71eb0ed8d1f70b4b33450b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id5c8ea61025914f6e5a9b5eab9269261;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic65f0f75f56bf85122a89cdf07e98152;
reg [MAX_SUM_WDTH_LONG-1:0]                  I924ef8499a83579e3449bbac0994775e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I41d22bafaf58e4a6de04640864653a16;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia8da4833c93e9ef6188709e7082092de;
reg [MAX_SUM_WDTH_LONG-1:0]                  I06a46b86f6edede0f5f72658a19910b7;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icd8516e6bf231bce29ebefbc7c97bff7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8591d0399594adacfeb006c5195c2c71;
reg [MAX_SUM_WDTH_LONG-1:0]                  I76c6762c515d0c9de1d777c0868b20af;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id90588b5f82cd32e801fbea04d24e4a5;
reg [MAX_SUM_WDTH_LONG-1:0]                  If5da296bcf91d370f8341fc402eed6df;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib642d757fae818cd6d713ffb6ce18fc1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I64673b4b013682f9ce54925853c06ca4;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id76bff2a12cf792e52ccc463647334c0;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iabfccf7b60f9be4e3714ad753cd8922a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I92ffa890ed6d83d4fc543504e4d421c1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I73ab1f85232818929b1b2e9d343584a3;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifc4a65edeaf630b3d29437bcd6c20121;
reg [MAX_SUM_WDTH_LONG-1:0]                  I06f989f65e614903ffba3594e8112235;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id57a11f56fc223501a9b68b8b05ebd3e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0391247480cb6bd6bda2c59dcf8f7607;
reg [MAX_SUM_WDTH_LONG-1:0]                  I522ba8bfc1949337e8befe82cc1e86e6;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iee114a92d2238e4b8fcdfa79c4c99d6a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7153e27c44ebbc2f04e9ba03cf09b5e1;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ida429b8e252b80b45435af1c6522f783;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id15e4b4f186ec863f12a54acd8ef8963;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id3849d43e39d78fd2428109bf9677e0d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I95c77eec7575cd7aa93a36f31ea635a2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5e51799e585f3dbef5e64908bcfc3e7a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3c8114dbe0658cc2889c787f1366abfa;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6d12e4545b8befb8d09545ea00c8ea96;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ieacf971e9e10fb73c7df9f1da8372f30;
reg [MAX_SUM_WDTH_LONG-1:0]                  I98d04e6bae91796784a864c5bed637cb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I35de1b03ea865f2c6381ce73e03dc220;
reg [MAX_SUM_WDTH_LONG-1:0]                  I83b3247bed67d1e2ed488d5b7812851d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idec12e02904ea98c7580919584f2dba1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I868021f44830a9d81c4ba3dad804f889;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia370c83631a2c1bbf39c7264deafafb5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I685e59e3865058f29978a8cc2f1b6c7c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I05b4a07dfc0d2695eae34bea4c1c6565;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5a76dd9f4a2078dee81102a9f205ca53;
reg [MAX_SUM_WDTH_LONG-1:0]                  If1ecdc27e3419dd1434e403f237c2b58;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ice3bd7a4bbf0705a3dc1f89c5ceca084;
reg [MAX_SUM_WDTH_LONG-1:0]                  I039c552777d0fb40bebcdd2d4a3394c2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5f741a3213cecdf58440120c2ea78e87;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iaa52fb63184514b6d754bcc896235150;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idad89ade7f96091abfea876b3af0d5b4;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ied9781e625c1fa8741853dd6b8b3a9e7;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie0ab4b7c79196195db0971e7c7a85adb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I767272262e9d2e85dba1aa93f578f25c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0093585d710940feaa8ebdc5fb000806;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib3b4cd6d8ab17869a2278552c02635c8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I76a0b74bb633743ac56cf4a0d52f80c0;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie7a5cb2ecb3fce35825785b9bca6b3bd;
reg [MAX_SUM_WDTH_LONG-1:0]                  I11931fd13219c1ae615d164a8f4130f9;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib9a0f8efd3dad427f247ce90fdfb94a4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6de7a344ae1574e551c7c10a1773d880;
reg [MAX_SUM_WDTH_LONG-1:0]                  I69a221a1bd95a588aa74b9bed0357762;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4920b0740cb56988ba4fc10b86195cdd;
reg [MAX_SUM_WDTH_LONG-1:0]                  I64f125cf2ca6a6da8a9cdae9e246c24a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I37d27fda03770ad37a1fbad835c076c3;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifac9dd60dd6c543aa94b39c599f0819a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib868fcb71300c09a49719e0b0459ca06;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icf062382a1e462571569ccee75b0a3ee;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2c67e89b58d7f998c43c68d857fa2381;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ieed8b94295bed265961c4f52c3379914;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idb770d9fc630f77beca27c3182279001;
reg [MAX_SUM_WDTH_LONG-1:0]                  I165eabcdde76821fdc308ff7a8c6d2ea;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6ab74c183d97a5df7a336c6c66c66e2e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8b3542a6d64d6a7ebba4124bc6702f3e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic4fc6d6a69dccb796d208aba87ec002c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7b68afec199be705d766c169f1ece981;
reg [MAX_SUM_WDTH_LONG-1:0]                  I450cd05f0109ad62ae4ca7f540ac7505;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4b6c8226ef2bc20dbd31d242bdb98b8c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia6f1bdee90a01ee3f3e59eec00689d50;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic3b4a86f22caf5b6103d52b6c9d2a991;
reg [MAX_SUM_WDTH_LONG-1:0]                  I33193403a8d72dcd02e87ae03b668e09;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia37592b207086f63e2d94e3d7d26c740;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5208f3202b32a30c4abaca4c617d3b3b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id0d786026e3ab0ddbffbc20e4d409857;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib607167c806dd831aaed4a42b9cf4349;
reg [MAX_SUM_WDTH_LONG-1:0]                  I333837f976cfc7f90ab0a6dcd8c1ce79;
reg [MAX_SUM_WDTH_LONG-1:0]                  I42b87e52c168abb775c1e1e5ddfc1958;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id115b4708a49dcfd167e79ef6993e371;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifc4e50801a1606717efd57bd5ac6f41f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I666da645400344644e848ee6f7592d3c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5e7282e9a35cead2f4d1d9860d45852c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibafeadd691eee03f855ed657c01022c9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8503b90594f3d4b492cca9cf154fc3d3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I10ec5c43a3fb65273053063001307280;
reg [MAX_SUM_WDTH_LONG-1:0]                  I95010cdf08c373916ab02e3794afa77a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I05c778eb3588bdaccf714ba456f534c2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I832fdc71e665ad2acac2576188e0d65b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icd11e8d97a6ac6c0a73e8adee1f98c4e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic21a6f1abcecf14acaf2aa23b7dcdb6b;
reg [MAX_SUM_WDTH_LONG-1:0]                  If07c2223d4262e22cca9b77c3ed5ee01;
reg [MAX_SUM_WDTH_LONG-1:0]                  I49847c8c979d9ed82be80f62552e97bf;
reg [MAX_SUM_WDTH_LONG-1:0]                  If0c8ce0ff66fe2806448f1c819d58ec8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7a2bfe5efbe1d0dc222bff675c621485;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iccdc2371dfd9fda3e506adc2b1681ba3;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie0d874ce4b0713de7d087396a1879c54;
reg [MAX_SUM_WDTH_LONG-1:0]                  I26e61dca9d045c4661b97afe346152c8;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iaf4c12394552f42e476b70f6c75003d7;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id488d650b86f5def0668f4a1ef841b6a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I64d7f4a0df87ce07ce49350610122f79;
reg [MAX_SUM_WDTH_LONG-1:0]                  I479365266255d2228ecd86c350e8d38b;
reg [MAX_SUM_WDTH_LONG-1:0]                  If51795ea140bec96fdefbc52291801b5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I08d9c488fd85db45344e649699196263;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib0a0f80cb818018b2fe0fd4597325bb4;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icde86d0ead44385b07e9a29057417417;
reg [MAX_SUM_WDTH_LONG-1:0]                  If01a65e097f026a816133c34d73ccff1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I21feecd24d912ef3d0aec0e375958f3f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ida9ed61c543afde2257053443d133119;
reg [MAX_SUM_WDTH_LONG-1:0]                  I59f419b3bc183a5fe743be3878fac587;
reg [MAX_SUM_WDTH_LONG-1:0]                  I983a5656d68192a7a3d5a78f17f12ff0;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib0804d8bdda49ecd0024300eed52be53;
reg [MAX_SUM_WDTH_LONG-1:0]                  I315445ad2d762b66f94a75d76fbfb839;
reg [MAX_SUM_WDTH_LONG-1:0]                  I37b0efdee34647a5111d698a5a80f367;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7a97a8fe65e56b0a80c242e13e70db09;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id382a04e94d0749d0858041bdc5861be;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2243095f420e4d996f1c69c965932778;
reg [MAX_SUM_WDTH_LONG-1:0]                  I368be992a21201268c41506396dcdcf6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0154a19f9adb43089080304978256c09;
reg [MAX_SUM_WDTH_LONG-1:0]                  I603a008893b5196d9f273b47a9d63144;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib8bdc3b41b3cc7132c43833802115880;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie70d3a768bc09ddff6ac68aaba7d9f2c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I167586906b601ffc473a5b856b213f2b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifb8bd837ada3d8ed5116db29da82d2a9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I094a6ac91aacfdd2f8de8a0d776f732b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I978b93d46e20cb3eda70e5a976d62348;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9d4437c250c28653bbccdea6af8b6280;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib404040d4fb58f47f245184c3be01789;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4afab82ea1a6ad0a36fea0692de1d106;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9c664265c53ebffaad097b70ff3cbbce;
reg [MAX_SUM_WDTH_LONG-1:0]                  I864d41b77a51fda97ea7017ed18b5fea;
reg [MAX_SUM_WDTH_LONG-1:0]                  I781306c6b1ce0741d9c2fa06865f7a19;
reg [MAX_SUM_WDTH_LONG-1:0]                  I758ee12b430cda151b452699eb2039dc;
reg [MAX_SUM_WDTH_LONG-1:0]                  I16fa2e3dc0b3eddbc72811b51d6ac8ed;
reg [MAX_SUM_WDTH_LONG-1:0]                  I134cd61326b70030c027a3821d98a994;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia6f232495726806d01b702b0e248b2f2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I99951d295b9065614c103b3e43fa255c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I66b3734060600caa45d699508c5083d2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I31a4e4f3eac271c84b36c84d7de338fd;
reg [MAX_SUM_WDTH_LONG-1:0]                  I85fae6b23d086235a94a0162e2fb5310;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id36c36d2b2dd9a79f9887c9950b385c3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8d6443d1be42203cb834345ae7e5aff5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I59455b0e53bac4fe6b1cbf609cb03da5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I717332b7f76e9caf9351f1aa69b72a12;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifd633f2ea91cb88aaa2a0bf5579ed1e0;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ieebd34db071409288f489129b70ab599;
reg [MAX_SUM_WDTH_LONG-1:0]                  I87218b174c1db735ac153604b5ff3e15;
reg [MAX_SUM_WDTH_LONG-1:0]                  I917c874137d64a9a495335c8f8ef5374;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4608c92d52306432c114f31b9ba6dd69;
reg [MAX_SUM_WDTH_LONG-1:0]                  I15fb4fb838d4a614c468f7d49261bda3;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iba3f6cde40827d82bc32078344b9bd81;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2eb093d2a38ba8cf4be47d1d7f54ecc4;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib987bde3ee5a0256d0b8b3aa7357cdb2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8f9affdc5cda0fecc35dd15fc5aeb244;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3c33a2bfaa82172457b15f4f621eefee;
reg [MAX_SUM_WDTH_LONG-1:0]                  I615a443d49d1479338d033d2a2cab51f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7ce33eb337b6cacaea13f748061e338a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0635a3270a9653ca0f23c116fd5b2f97;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7a8c5be75d87552ca717a87d1a832d21;
reg [MAX_SUM_WDTH_LONG-1:0]                  I93a7c75ebce8fbf4c613b4d11dc98b72;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id9c9cebf44647040da33567d815c261f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I39334aa9d55bcc001ece37ce2a6c329c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6c522c28a0dc265facb1f21ebe51c564;
reg [MAX_SUM_WDTH_LONG-1:0]                  I07e328d23da9383a296ecb03679ec74b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I86c367b0fd4548d5edfb8863f454653e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8a6e1eace6152af5c98c415804cb60fa;
reg [MAX_SUM_WDTH_LONG-1:0]                  I800271efe85fcbaee8fe733190e90f6d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6ed4d6c350e8691b3a12ab51419cfa65;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia5172996abb4a6bc50046d36ec033c7f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie2b9ed680dac51ac866cb830ca17ef84;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibe20363746d437eef2c85360425739d1;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie439b520bbb0c8b29a5ecea167acb1c9;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iee695b22e8a55479dfcbaa68f5c8b6c9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9f8ef3295578acf5b0a42d074a15a70b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7cdb0bf6c7195df38d701768e655af70;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ief01b06341d489e36ee344fd52084ccf;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1057373671fd4cfba6696f8e88a2d740;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3b72a085b104e17dca3d8b2824f84e97;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7dd9da64c1516e6ae1b703defc4cdc55;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5e1f41e23887493db1d723e1e2cbd996;
reg [MAX_SUM_WDTH_LONG-1:0]                  I58bf5f51208a98b2448e2b4fad3f63ac;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0e6f4c7bdc39bd22833f3d9fcfa55f1d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icb8281c05ea7168d39d6012a1d622e15;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie346802a8898b4b075be289e062b462c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5b16ad2952938bc64f6c9f5ff1ab5a0b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I82ea6f21706a97166ef11af548e80392;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5d5790b480d08bf6c957f26e24467b9a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5f38764f6ecc2dcd1fdd5316102f1f82;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ieb32ca618265eed3419f01907f48527d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id4034bf7a0e92a6c92d0187e00d3df99;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ief90415b272ce5707ba28a8470132f5e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I44692fd63388c57268ea9035a7e4c3ef;
reg [MAX_SUM_WDTH_LONG-1:0]                  I386c79f4301dea9a37c9ce283e8050e4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0c2892a34e5236f1366959eadfd83825;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0d113fab9d7095f8d1693fec58b7c5a6;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iccef2754044e7066e191bc5e1a3805f1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2bbbe9e5d322d9cee76903fa813765ae;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8ace46f1c56cfb3f4773324e0f8cae58;
reg [MAX_SUM_WDTH_LONG-1:0]                  If5317506b6ab92c946af745a65b9e86a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I94ec0139bd827ef5dce2c5ee9eb9aded;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib61ddb3ef6c7239bfc720b1761cc0221;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ied62b116607c549ff5918d5b95e2118f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I70d669976b271b2319d60114c468cae5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9efa5796297bc922bc5fe17f8319a515;
reg [MAX_SUM_WDTH_LONG-1:0]                  I96cb81892e2d1737d6cb25522ea2d9e4;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifa6908d8fda29713d7c1bbaa69b72b53;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6c87926b040d4006c2294c516a3c46fd;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ieb46857229186ce0391cddb2d30f434e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I549670efc854cdc29bad1d9bc03e9f5e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I67fa03f808026b38ca5b4e71e21588bf;
reg [MAX_SUM_WDTH_LONG-1:0]                  If54c0c169048bb3e8a1423a58aed0e70;
reg [MAX_SUM_WDTH_LONG-1:0]                  I70938dfe09b0da9d87dafed6af3fa05c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5c956f39031611db595fbc34e6edad65;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iff30a4e14b6282e9ef92e7f58230b516;
reg [MAX_SUM_WDTH_LONG-1:0]                  I86851725f5d424c4636f9f41e5a7c7e9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I43e0faf8070869ab0528a7a4a5cdc103;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibec300322cef05615c818b163f8a1fef;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib2f0333fac7701ae4a5589d54005b8f3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I09cc443ecf3811a8a672c4aec1f7d6d4;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie4e1491da700923e81b2c1a246e528b1;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iaaf5b9288b4eb557d56908bf072cc642;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie8602467de2ece2013878a6b8d3129a1;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib224ff2bea17f6e694b10bc7cfdb898d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I85c93c62f79b1703cb6928f96737cf27;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ide7d6472bf33f8dcf5c6397c7d7fb733;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3dc816ee6c2a818b32f6d4e1228704bf;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie6193636ea1cba8b71e1d0d5f2e3c1b2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id34d83701e815c01359bc5cd1b9c993c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id631b0a4de889a3c3eff4df79367d3d4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0a20e3e26261ba558d681346649cf0b3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I93d80b8bfb77e7af4d9ac734f26c4e62;
reg [MAX_SUM_WDTH_LONG-1:0]                  I331c6e8dbe2ea1e2232f82766926d0e6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7fba5fee37c5912e7f635feb8c111b3a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie27046fd2751357e4a81dc62086f00be;
reg [MAX_SUM_WDTH_LONG-1:0]                  I22c14ad43399d8a1aee258826a71f50e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0897ceba8201bc14a49ab30318183875;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3bdc4806c5c09de9a7de8d3601c57bfe;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie7b15aa8ce2492bfb433894efeb967f3;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id451569510e0d1bbba9002c2b27bb3d4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I255add08e982f701508a98db221e617d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I16753a377bced0688797a464157d847b;
reg [MAX_SUM_WDTH_LONG-1:0]                  If7ca4919fa1449f38777f742ee1fb875;
reg [MAX_SUM_WDTH_LONG-1:0]                  I76fd17f22401b66bfc0a6239a0518157;
reg [MAX_SUM_WDTH_LONG-1:0]                  I24cafcb5b9825321c54e84827a662fdc;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie56f8b245ab7833b6939cfea43a99874;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3ede71cb7cb39774aedb9889240a2462;
reg [MAX_SUM_WDTH_LONG-1:0]                  I668f8103700f044c7764f2281a5b457e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I24da9598a6840d3ba7b12fe4f638219b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib75c0ca4f8b59afc2fdd7793bff7ad16;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0358ca8833007cec4ce5047db32ab7a3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3d39fa04d24aa69d19a2db8da00eb0d3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I85b5354463c1c15f91ed67292da912c1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I284b4ccbcb23293efe64fa45b2e0ad98;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie93731739ace44811198d0fd95b04a6a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I689ac029a268fe244a8793367c900602;
reg [MAX_SUM_WDTH_LONG-1:0]                  I464926faf4e005ad491b0bf93a365e07;
reg [MAX_SUM_WDTH_LONG-1:0]                  If53dace3e8a7be2524d711de84855015;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icdaaccfead6f2d5ac2ce19caf1104d57;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie3fe635b63e13732c17ae2076b807b4d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I916d6f9429f2b0cc1bd6fb900484cde5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1e196a61113d4db7b51f3d6b18c33da3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0142f9b3d361a0d88522f1c5f54aca84;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic80e494400a5d7dcfdbf96424391e596;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie6871983b4f81b5321519647e628bd0e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I69d20a7aaf2c66ed9b41fdeff0d5c6ec;
reg [MAX_SUM_WDTH_LONG-1:0]                  I17d7be125df22153fc1ed051d4e0770a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I19b667bdb053ebd555aaa540d3a76f95;
reg [MAX_SUM_WDTH_LONG-1:0]                  I50b13959e06243e54fad2088eaf65aa7;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifc3d9cc420aa1274fed24b38c4d9fd8a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7a423d609b492f73d5a322849b4b1cce;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie8a6ed15370edd38bfc92290bf7bb55a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iefec67e214d1868670a34a7297d4a1c8;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ife5a1b49d4b0342f06ef83750ab914d4;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iae7da7fdc002b635ce4285d6916d8156;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9906c49536062867b98ed290e49bbe50;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic561e44b2caeae84df6720f1afa3e8f6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I41be66295070bec696e91d0f9efdc233;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5be062f5b52e104ca67e615ce75a7c80;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4838b956d8a597e78bef9a0fce82542e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iecdde23e34c34ee0055be41f44959a19;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia06cb40e9a3341f34625c5804e02c07f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibe09be9cad0e56d5403868d072d7d628;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4eaad70758412eab097822b2feda7a57;
reg [MAX_SUM_WDTH_LONG-1:0]                  I464e1f3c13acaf466afb354a9b35ba0a;
reg [MAX_SUM_WDTH_LONG-1:0]                  If89e1da3daa6fd3090781723173b140b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I160a465c22073a53510e8a4c489c3321;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9ac67c519fd5a55d0ffb727389781492;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9e86d3e49827861b24f4fbeb308ad3a4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I73799799e5469ae887dec9b46c9c965d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib96b7d796e20967e89a47e01bf424e59;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7ebd7c3f0617cf500deeb8c152c09af2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I565e666f6ba14b4c25e0dd402a3266e1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2ee7d4f522ba17ca941c67079309c398;
reg [MAX_SUM_WDTH_LONG-1:0]                  I97e8bac5becd5128bc70f3bb48f73e6c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I62d13683ba05cfc27d9ae9a82fb04689;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iced39475c6e5e3d8f36d2a5c5a80f146;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic06032eaed49f01d3d5513b2d145eaaf;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idcbd423c2b963c1f693dea2ddf428195;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idba6350812d3c90bee79636db48257e2;
reg [MAX_SUM_WDTH_LONG-1:0]                  If1640e294bdcc51ee12fca5b3a33be6d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6e7ed391604c7e0ff7cca99d5aeddc9f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4754c6c355e632d2ed1336b5a88c3b46;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib78d45cc282f110ed3ddaeb706a0fc12;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1634d703ad5d6e58a97b13ef957bdbec;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0f5d081f9846ad888eac13d4916f5b8c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I804e1e6a01edeb780b0159ecae707b71;
reg [MAX_SUM_WDTH_LONG-1:0]                  I607bdd63c3ee70e2721de3f994d2923e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iea3c0f3c3c3017fe87a3b01647189fe0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5453775d628c6c01c088278b6e090ddf;
reg [MAX_SUM_WDTH_LONG-1:0]                  I756b7d7e6bd3e71afa472e7e4727264a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iff51257cd95c2f3a38c64ae872317410;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifbeae0a2acf80eda6ffd050d3bb07eb3;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie5faf4f522c8d24bc2d3725be57453e3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I990ab4dcb70ee860c2c40f306ef314d3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7952b4b62af35c930dcffe35b1629100;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib131087ea9ccc4bd161c3f9ac2c72303;
reg [MAX_SUM_WDTH_LONG-1:0]                  I47337a0b371f749c3f7f5118362c2301;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9a967ac9d11583faaa783984229aeb2c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I21ea597751b3243936aea7c07cc90f70;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib9921dfcf121e5f4ac4d8be83a868210;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibdce05e98adef0314000dba3c482ace6;
reg [MAX_SUM_WDTH_LONG-1:0]                  If22d8fd45caed08b2c7cee8b7349700f;
reg [MAX_SUM_WDTH_LONG-1:0]                  If0dbc84f59311eeabfb57b5fd0c3b632;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iabf029e67c7f827faf17b6518cd1bfa3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I74f2e7798a8383b78a5e7b816c2370af;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iaeab83001c6285630e3404ae67227f46;
reg [MAX_SUM_WDTH_LONG-1:0]                  I58ee302a3a1faa2b44d9052bffbc2a03;
reg [MAX_SUM_WDTH_LONG-1:0]                  I53ac6d02d2bfc9aca9469148753070a7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I979a71fc0942bf62c06405bb63a717c5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I61992979f60b26d313efd1dc23bb54ab;
reg [MAX_SUM_WDTH_LONG-1:0]                  I30be0ac758b5a0fbacb1c51a36ca8a73;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8b46b3f0835310114208963de7ac8e97;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9c50e0a8a01aaed98ae54530d5c76ba1;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icda26ba6f5c7f77a80776b2c1bbc975d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0daac80ebeec26e428328344a398ce57;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0863565b3ae88137a2384750436f9e19;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6739f13ea431943bb5bacb4a05140063;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id646110f8d09cd47dc7695e05f73efc6;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifa0e560fe6445b006ab74096a807b90f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5999eef2304e579a3d47e4f15ba336e1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9595c0fd77d6a0610eb859dcd2b67d1d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idd302bdc6ff8368a6b73d53bbc8f8425;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6f3e685e70fa700b52bec62d0aed942c;

reg     [22-1:0]          Ib58043c04b5c4c86c1c67e57cc66dcf7;
reg [MAX_SUM_WDTH_LONG-1:0]                Iea07d1adf9016a29cffd61d183e268d0;
reg [MAX_SUM_WDTH_LONG-1:0]                If92db65b39a83e1c699e4cc6d7f9e57b;
reg [MAX_SUM_WDTH_LONG-1:0]                I8f2986bc015fcc64ac5e5395ac6dd851;
reg [MAX_SUM_WDTH_LONG-1:0]                I355725a804e0df68b4acf96ca98f2448;
reg [MAX_SUM_WDTH_LONG-1:0]                I78212ae965ab2dcb2eed0b060d6b253f;
reg [MAX_SUM_WDTH_LONG-1:0]                I0b56aa7a1b7549c91dddd3a06ecbaacf;
reg [MAX_SUM_WDTH_LONG-1:0]                I71412803cc5229025487255aec62ec4f;
reg [MAX_SUM_WDTH_LONG-1:0]                I32fcb28a27356bc6f403528836ea4c1f;
reg [MAX_SUM_WDTH_LONG-1:0]                Iad354d876cb9fc72fc0143e6f7da9357;
reg [MAX_SUM_WDTH_LONG-1:0]                If6e745bb85abba7282dae1f6f701225e;
reg [MAX_SUM_WDTH_LONG-1:0]                I93bb43c1b89d4c70a57bdc019d64fd22;
reg [MAX_SUM_WDTH_LONG-1:0]                I7a2e554d07bbea291f2cfc18694fca3a;
reg [MAX_SUM_WDTH_LONG-1:0]                I3e59b2419c7dd1553b792d536208514e;
reg [MAX_SUM_WDTH_LONG-1:0]                I46894c6526983bf1ce4b503159131b41;
reg [MAX_SUM_WDTH_LONG-1:0]                I6404d0df952b5bf8292c753e4c6f35d8;
reg [MAX_SUM_WDTH_LONG-1:0]                I8522c402e654d007abffcb0e904af5e6;
reg [MAX_SUM_WDTH_LONG-1:0]                I5ed85845c39337c37791f16e718069b4;
reg [MAX_SUM_WDTH_LONG-1:0]                I89013d61c1ea8da8b1c6071cc21c316f;
reg [MAX_SUM_WDTH_LONG-1:0]                I4102100fa5f1dd299af0190862efcc42;
reg [MAX_SUM_WDTH_LONG-1:0]                I4939f69abb1eac56d5021e06406a93b5;
reg [MAX_SUM_WDTH_LONG-1:0]                Iadbd245bf842aebb456417579a3e6296;
reg [MAX_SUM_WDTH_LONG-1:0]                Ifc8ece44a4e68c3117eda9e65f3084d2;
reg     [22-1:0]          Ibc0871b3c992fd278815fdbefcd2bac0;
reg [MAX_SUM_WDTH_LONG-1:0]                I91679dfab57a372eddc7f9b94a231edb;
reg [MAX_SUM_WDTH_LONG-1:0]                I2213c1a2b831f421707a261f5a58b1b1;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic53b875b2ddcba11406eb2ca39354757;
reg [MAX_SUM_WDTH_LONG-1:0]                I634484f00590216c0f74f975c9c83400;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib3b1db2d8b669988c887ed780e439b26;
reg [MAX_SUM_WDTH_LONG-1:0]                I735db8b0ee0ec98e4cce0030b11508da;
reg [MAX_SUM_WDTH_LONG-1:0]                If1607e907e626902ee26d15020a64c21;
reg [MAX_SUM_WDTH_LONG-1:0]                I081b38dbb37d4c14a6a9fd3fefa13daa;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibac5e7b6d4bf5cd6926358318f0c418f;
reg [MAX_SUM_WDTH_LONG-1:0]                Iadfc60386481092ae85cc148a2c40abb;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie0ee5445c56a5f9b41640b57422206de;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie5f8620371236cb11c9e88c16b509ee8;
reg [MAX_SUM_WDTH_LONG-1:0]                I8d7c1fe2e33bbd45379b0325a3c5e989;
reg [MAX_SUM_WDTH_LONG-1:0]                I4fbdc4ee57a3be42b62d9bd43078d6ef;
reg [MAX_SUM_WDTH_LONG-1:0]                I5510b88bfd65811b3200adf4ef975b48;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib57ef2f577cca54713c16717cbbd1ce9;
reg [MAX_SUM_WDTH_LONG-1:0]                I15943aa74e9fbbaebdc0d54eb6a3bffa;
reg [MAX_SUM_WDTH_LONG-1:0]                I6ac24c46319a787daa5c545de8c6eeea;
reg [MAX_SUM_WDTH_LONG-1:0]                I52403a0454e5fa002e79eaab7ea497bd;
reg [MAX_SUM_WDTH_LONG-1:0]                I634f0ce28934600a1a31ab0d8e59b4a9;
reg [MAX_SUM_WDTH_LONG-1:0]                I7103aa739616a39c03e675ea0efb0335;
reg [MAX_SUM_WDTH_LONG-1:0]                I0296d01fd3f9a269a617efd4beea9b8b;
reg     [22-1:0]          I8695e1e94cbfcbe4b9eae315b042529e;
reg [MAX_SUM_WDTH_LONG-1:0]                I065a81ba25962785215583e7ece27661;
reg [MAX_SUM_WDTH_LONG-1:0]                I631a3300cb6685f47da7781940ec5d27;
reg [MAX_SUM_WDTH_LONG-1:0]                I8bbe1a2ace8f51aa22cca5d9fc66f136;
reg [MAX_SUM_WDTH_LONG-1:0]                I38c3e3e136acb79c8a0ff850bcc55f16;
reg [MAX_SUM_WDTH_LONG-1:0]                I35b2c7e9cdc53a98913e1c16a3a47b37;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib1a2b31d49ae476e2f1fb9acba2d5af0;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic72f41f9bbf470aee3c9b9b8787b31c3;
reg [MAX_SUM_WDTH_LONG-1:0]                I3ea4c33a9419820ed54460eb64134dff;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia0d940e16c8cbd4f7544f5a5cd7d83b2;
reg [MAX_SUM_WDTH_LONG-1:0]                I4a8abfa0896ce414d9b98093ef84455f;
reg [MAX_SUM_WDTH_LONG-1:0]                I680be647bf2a62e0ee9b5d379dc87b4f;
reg [MAX_SUM_WDTH_LONG-1:0]                If4d75f83299a21802b6fbe136913489f;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibddfda6413e3dd2f483c3174ea836b6a;
reg [MAX_SUM_WDTH_LONG-1:0]                I33bddb0adcc2af7b12a83bf843036385;
reg [MAX_SUM_WDTH_LONG-1:0]                I529f92b82248efe2cf64f7da0ec8283c;
reg [MAX_SUM_WDTH_LONG-1:0]                I2f34af0036985cd94ade9cc905bec065;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia1a0d8d7dfd6e877f15cce773f85f5b7;
reg [MAX_SUM_WDTH_LONG-1:0]                I5dd29fd1a73df5662d2b636e7285bad9;
reg [MAX_SUM_WDTH_LONG-1:0]                Ide530e6f4622c8a7b101b6dce9650e42;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibaf00a6780325882067a79f0c4d693d2;
reg [MAX_SUM_WDTH_LONG-1:0]                I16e3559c63ebfed83d6698fc9a9cd93a;
reg [MAX_SUM_WDTH_LONG-1:0]                I9747a02384abb1c2dd1f52b3a5a999cc;
reg     [22-1:0]          Ifeb6f8e9d7d86fb01ee8faed3bad6d6e;
reg [MAX_SUM_WDTH_LONG-1:0]                Iceb7a1d4c23806b8f5824016779ad129;
reg [MAX_SUM_WDTH_LONG-1:0]                I40ef50004a60ae58aedc49eb5e6797c9;
reg [MAX_SUM_WDTH_LONG-1:0]                I753f92da60980736440aba814a156f1e;
reg [MAX_SUM_WDTH_LONG-1:0]                I4ac79b67a8904b95f7912d24af420585;
reg [MAX_SUM_WDTH_LONG-1:0]                Iad44c932cfa5c249c5e59f8c706173a8;
reg [MAX_SUM_WDTH_LONG-1:0]                I10f14b6433498e3b9e9bf021b60115e8;
reg [MAX_SUM_WDTH_LONG-1:0]                I96008f47b9f134c9c4274cfcfb28e550;
reg [MAX_SUM_WDTH_LONG-1:0]                Id0344146d1a53d418add6d2b185377dd;
reg [MAX_SUM_WDTH_LONG-1:0]                I1eede74f12d37331b399eb7136bc621f;
reg [MAX_SUM_WDTH_LONG-1:0]                I3e4754acc31d99bc71525789bdee0c1a;
reg [MAX_SUM_WDTH_LONG-1:0]                I11c1fc94a3bd6dffa17e1571cc6ae97c;
reg [MAX_SUM_WDTH_LONG-1:0]                I5395ee57418c31e11cf847f0f514ec19;
reg [MAX_SUM_WDTH_LONG-1:0]                Iff125392fa39afebae1637a19c4e23ec;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia6308e16fae5428f4ab6560f5b21479a;
reg [MAX_SUM_WDTH_LONG-1:0]                I5ea02b5349cd4d99ccbcb6b26f0cfdd7;
reg [MAX_SUM_WDTH_LONG-1:0]                I21de4f6194dec9e3c401934db92c25e7;
reg [MAX_SUM_WDTH_LONG-1:0]                I57d0920119f8901bd4dea2d5f8fb5d90;
reg [MAX_SUM_WDTH_LONG-1:0]                I89537301987d6da0dbe6cff3caab3ff4;
reg [MAX_SUM_WDTH_LONG-1:0]                Iaf0bbbe791bb71d0f557dc71caa5fb87;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic7ff9cde71054c1ee9eef81eabdd7061;
reg [MAX_SUM_WDTH_LONG-1:0]                I88c10c47ae424fbdcb852fbf1e94127c;
reg [MAX_SUM_WDTH_LONG-1:0]                Icd2e75e47cab1d539ba9ff1b6e1d7155;
reg     [23-1:0]          I61f0c04673dfb262ef6912eb2df39120;
reg [MAX_SUM_WDTH_LONG-1:0]                I37e6bc7aff363ed0ed1f84b23c5f3e34;
reg [MAX_SUM_WDTH_LONG-1:0]                I733605337bf6972630c089d32fd7f98f;
reg [MAX_SUM_WDTH_LONG-1:0]                Idcb1d8bbdeaed6768c2a418c3048e6ee;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia89da2f1890524ad3519ab403dd0686c;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie33a780b0221084898c9fc5b237b244a;
reg [MAX_SUM_WDTH_LONG-1:0]                Iabbd1668e0014df518ede5216232834c;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibd89458312687610aa166a9538968851;
reg [MAX_SUM_WDTH_LONG-1:0]                Icbaf92a8e9875bcb19a1d074779a9ea5;
reg [MAX_SUM_WDTH_LONG-1:0]                I80f3c8559da8e97bc5397bb8b621a0bd;
reg [MAX_SUM_WDTH_LONG-1:0]                I7a0eada108891aba06cecab5071232c9;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie21a2c9b22e7bf8425fb5c0f33e5f4f7;
reg [MAX_SUM_WDTH_LONG-1:0]                Iaa5b2807e5cc2403c5787eeb3d10ca6b;
reg [MAX_SUM_WDTH_LONG-1:0]                I6da2b3a481ee71b85f3087b36b399288;
reg [MAX_SUM_WDTH_LONG-1:0]                I11094e852295755925c3c61f1df81643;
reg [MAX_SUM_WDTH_LONG-1:0]                I9c633aa620cca127b0ff8cf882178e76;
reg [MAX_SUM_WDTH_LONG-1:0]                I694d471fd353eb54aae08a2afa7b645a;
reg [MAX_SUM_WDTH_LONG-1:0]                I816704585ad393f685731104ad3ec64f;
reg [MAX_SUM_WDTH_LONG-1:0]                I85d95015a9ce27a18ccbf73bbbcdbd70;
reg [MAX_SUM_WDTH_LONG-1:0]                I992e7c551b4aa818606c3465d33eb798;
reg [MAX_SUM_WDTH_LONG-1:0]                I2ead0e9941e2280309ab53535b1e1ac1;
reg [MAX_SUM_WDTH_LONG-1:0]                I56873feb8418005b5661c7382f2dbeec;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib6ea4a822da2ea32e0abf6cf8a33d295;
reg [MAX_SUM_WDTH_LONG-1:0]                Id1659ccdeaea3e59eb2d3f65a65ebd05;
reg     [23-1:0]          Ibeb5edab51cd6aedad9c2ecedaded6f5;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic2171967791a0329f3e39fc19d0a6bc8;
reg [MAX_SUM_WDTH_LONG-1:0]                I7d5041a6796c00188f74936d283defe6;
reg [MAX_SUM_WDTH_LONG-1:0]                Iba7608ee0a01af103e022bcaf564bf6b;
reg [MAX_SUM_WDTH_LONG-1:0]                Iedbe9d0e48bd36064f59faea51afddb9;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic3871325d57b310c95ca02fcaca529eb;
reg [MAX_SUM_WDTH_LONG-1:0]                I42f9b1f8ef24ad56c10086852678b456;
reg [MAX_SUM_WDTH_LONG-1:0]                I3ed5d0fca86f35b3d4b4a89c6147d0cd;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib0126fb335e32793c400a97c5a4a337c;
reg [MAX_SUM_WDTH_LONG-1:0]                I20590d8fb97ec0b2164ffe17826136a7;
reg [MAX_SUM_WDTH_LONG-1:0]                I3c128efc9f80c9b8334bf7b61de71b43;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic7147944f8835e26b9838fdbdc18ca41;
reg [MAX_SUM_WDTH_LONG-1:0]                I698b1dbc9d8664d1c86c7a763d97b3b7;
reg [MAX_SUM_WDTH_LONG-1:0]                I508bbade361787127e1a2e8687ec884c;
reg [MAX_SUM_WDTH_LONG-1:0]                I2afeb2a7b199c0c6738938f156ae4274;
reg [MAX_SUM_WDTH_LONG-1:0]                I86255756ddd1f88b74e070b19f8c3bfa;
reg [MAX_SUM_WDTH_LONG-1:0]                I7d4924388dc5373ad7936dca76797473;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie317e5ea2ca4ba2060d0f491290af96f;
reg [MAX_SUM_WDTH_LONG-1:0]                I56ea52c50a188ec47e48740839a031c9;
reg [MAX_SUM_WDTH_LONG-1:0]                Id9b9a8fe43992ec0793845715dd2226c;
reg [MAX_SUM_WDTH_LONG-1:0]                I93b69bfb228db4b569a6772179d603be;
reg [MAX_SUM_WDTH_LONG-1:0]                I71afab29cdb962e1f1ca21b61dfb50c6;
reg [MAX_SUM_WDTH_LONG-1:0]                I9905e2686b350e8a6e7f790563a91294;
reg [MAX_SUM_WDTH_LONG-1:0]                I524e78ae6a4204e17ba4532dba047d4b;
reg     [23-1:0]          Iceb64ab2ff8a2e0dfdb74803811d4cfe;
reg [MAX_SUM_WDTH_LONG-1:0]                I71228fe4188ab1d9796081184a422094;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie19b39200436b0bfca13502ad36c21b9;
reg [MAX_SUM_WDTH_LONG-1:0]                If6657f90c84ca5e2ba08ec705f34be03;
reg [MAX_SUM_WDTH_LONG-1:0]                I60ec7459bbe99fce295406bee1f2af46;
reg [MAX_SUM_WDTH_LONG-1:0]                I29ab844f80c105d247c5c15faa35863c;
reg [MAX_SUM_WDTH_LONG-1:0]                I856fa68463aa5ef1ae53442699d38b33;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic3d00a27f15f8983a120395082854d6b;
reg [MAX_SUM_WDTH_LONG-1:0]                I6b1d01c3cb8fb51e43cdb788b89816be;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib74a56900c1f8b159ad381f61acee801;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia5eba52d169755c507b9e0094e467fab;
reg [MAX_SUM_WDTH_LONG-1:0]                I0899e8fec1a7209cd94757c0b2f87c9a;
reg [MAX_SUM_WDTH_LONG-1:0]                I08ece7cd684e593e02321612b7a88cee;
reg [MAX_SUM_WDTH_LONG-1:0]                I691c84d81c60a462e28e2b2bae3ea845;
reg [MAX_SUM_WDTH_LONG-1:0]                I58dc9cce6384160c0a85c6efb3319cdb;
reg [MAX_SUM_WDTH_LONG-1:0]                I56bf74b5890ec67090f499afdc0a9c88;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibaf2f1f8bda2f6b932dc30f8369c0e1f;
reg [MAX_SUM_WDTH_LONG-1:0]                Id9364a29fd79b52d0442e18dc0227854;
reg [MAX_SUM_WDTH_LONG-1:0]                Ica3a41ace27f7d94377981079952f4f7;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib57795a63d642a73456324bab41384b6;
reg [MAX_SUM_WDTH_LONG-1:0]                Iabf572c97b48c6a7dcc19e56676e3a82;
reg [MAX_SUM_WDTH_LONG-1:0]                Iefd370d0df1a93639af482f78a1e8706;
reg [MAX_SUM_WDTH_LONG-1:0]                I995d2809ffaf0ecda6a004d01cb9c8c4;
reg [MAX_SUM_WDTH_LONG-1:0]                I4e8ebc46bc068c3f9889d970db131112;
reg     [23-1:0]          I5b7caaeb34c43e66e8d095a859e708fe;
reg [MAX_SUM_WDTH_LONG-1:0]                I7b561638da1b4a45ff59be81243e4471;
reg [MAX_SUM_WDTH_LONG-1:0]                If0a3b88a66a816b25f17ced5d0e8f775;
reg [MAX_SUM_WDTH_LONG-1:0]                I0374ada4fe50717f2158468b7ad205d4;
reg [MAX_SUM_WDTH_LONG-1:0]                I357137b41bb91e0659b1ac6ead9b5c12;
reg [MAX_SUM_WDTH_LONG-1:0]                I5d70bc64cf7b3d3ef4180e082e533237;
reg [MAX_SUM_WDTH_LONG-1:0]                I7d9ad929660cd212387d893266b681da;
reg [MAX_SUM_WDTH_LONG-1:0]                I34be4b353cf75603301372840c2f91c2;
reg [MAX_SUM_WDTH_LONG-1:0]                I14834fc8e6489775359bcecf5a37ff4d;
reg [MAX_SUM_WDTH_LONG-1:0]                I633a74e4dfa841c9fd13dbb6564c8493;
reg [MAX_SUM_WDTH_LONG-1:0]                I157bd468200e63385583b9045758d81e;
reg [MAX_SUM_WDTH_LONG-1:0]                I918c46173eebc5b2a95e041cfd91d958;
reg [MAX_SUM_WDTH_LONG-1:0]                I4f8792c18bd07b23e82bbc44b4ca947f;
reg [MAX_SUM_WDTH_LONG-1:0]                I8d0a1ae4c47edf1f2b99d1175aaa7197;
reg [MAX_SUM_WDTH_LONG-1:0]                I734e601f5f9d568a44a48834559e04db;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie421da1dc5aaea57c50d0c7d9c5a2717;
reg [MAX_SUM_WDTH_LONG-1:0]                Ief5cbddfbfb98fce4812a676849b9a98;
reg [MAX_SUM_WDTH_LONG-1:0]                Id113cab2dd1949d32e3c1c15273185c8;
reg [MAX_SUM_WDTH_LONG-1:0]                Icfe1a689e33b2b9aa9dba692d6d610b9;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia4b671f3360f3ce55db0dc0e4d78ddbe;
reg [MAX_SUM_WDTH_LONG-1:0]                I60cbd4369e7ba9b6532f279e5c59084c;
reg [MAX_SUM_WDTH_LONG-1:0]                Ifb6c65a00d9a2c31d8b1119b949828d8;
reg [MAX_SUM_WDTH_LONG-1:0]                I4a777f0dd62b19dd340ad31517c4e789;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib75747cb32130d44b338ed8c8af8ca11;
reg     [10-1:0]          Ib0bf69cc797f330fb2546eb46d2d6f76;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic7e35cf8d5cd230b94c40714f16e2418;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic51bb9184dfd103703cd0c6ad6edff4b;
reg [MAX_SUM_WDTH_LONG-1:0]                I103f1449c78c47396d6a54dc1c810934;
reg [MAX_SUM_WDTH_LONG-1:0]                I56b3a97dc3037f0bb2eed93a9482c813;
reg [MAX_SUM_WDTH_LONG-1:0]                I51e98035b35a35fdc52f5bab8f19c152;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia6a7f9beaceb08d81012f0e72171252f;
reg [MAX_SUM_WDTH_LONG-1:0]                I21b062856ced09cb9131c01b5e166f32;
reg [MAX_SUM_WDTH_LONG-1:0]                I4f1221ce7880729fe584b42ef3afe6b2;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie7f3f1d6cee7f02ae1b17740ed54c049;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib196f5bcf9152703dc32c5101076600a;
reg     [10-1:0]          Iec7404bc79c58d4d2538fcdf659e9134;
reg [MAX_SUM_WDTH_LONG-1:0]                Ide9ef5a16d8fe32353c2c2a30e8ee3b0;
reg [MAX_SUM_WDTH_LONG-1:0]                Iee6f2484a381bd42e441ff072ec582e4;
reg [MAX_SUM_WDTH_LONG-1:0]                I53121a39de0bcba91a4d0438be2ae958;
reg [MAX_SUM_WDTH_LONG-1:0]                Iff7950f24f0a6b0073942c37fff49d37;
reg [MAX_SUM_WDTH_LONG-1:0]                Ide86f019e9573706c25bd8b4552396a8;
reg [MAX_SUM_WDTH_LONG-1:0]                I2370042234b0e93bb66e44b97fca3e43;
reg [MAX_SUM_WDTH_LONG-1:0]                If9efe7a1c359ec03014a52870ac13aec;
reg [MAX_SUM_WDTH_LONG-1:0]                I6a6eb62960b616043415406ebfc21346;
reg [MAX_SUM_WDTH_LONG-1:0]                I06c7728ef64be8311f48d10d766d0c44;
reg [MAX_SUM_WDTH_LONG-1:0]                I9fe11f6c8147391aa4a5afd1a4e4f731;
reg     [10-1:0]          Ie1cd04c7668d3f450c387a6c1ad778c7;
reg [MAX_SUM_WDTH_LONG-1:0]                Id50edc56fce48130247fdbc42eeff9ea;
reg [MAX_SUM_WDTH_LONG-1:0]                If3e5161254eb9056914c46263b865c10;
reg [MAX_SUM_WDTH_LONG-1:0]                I58703e8b6d04f8c69ac38f5fcfdc4efc;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie1f41720e296ced1b74cb325b666d88f;
reg [MAX_SUM_WDTH_LONG-1:0]                I5d5701435c96f1078e741921b56e3c65;
reg [MAX_SUM_WDTH_LONG-1:0]                Id96e744d9b10dcddd1ae0115ea57a76a;
reg [MAX_SUM_WDTH_LONG-1:0]                I0c0060fe260afa3cdc72f35ffb6938ff;
reg [MAX_SUM_WDTH_LONG-1:0]                Iaec1f186cb4a65da21d41e637fc628f7;
reg [MAX_SUM_WDTH_LONG-1:0]                I9c15a6a5c0db11ede80ff6d04c9a56d8;
reg [MAX_SUM_WDTH_LONG-1:0]                I8922487573e02d684a3d71448c3828f5;
reg     [10-1:0]          If511a6ea6aa5cda5353658d8e192791f;
reg [MAX_SUM_WDTH_LONG-1:0]                I47f17afcd5871fc3ac378316fd3d7ae9;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia9642d79bb50567348083b4435c7d66d;
reg [MAX_SUM_WDTH_LONG-1:0]                I2b2bd845428c49346ef8e94e95b618f8;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib730fdb59198f23d1e590f6d6039e96a;
reg [MAX_SUM_WDTH_LONG-1:0]                I644e83f0a7d432fba38ffb2d99088eca;
reg [MAX_SUM_WDTH_LONG-1:0]                I97f2b15ce0a74e68d5a4438111adcb0a;
reg [MAX_SUM_WDTH_LONG-1:0]                I84c88b631bed5311cb6e99e58941149e;
reg [MAX_SUM_WDTH_LONG-1:0]                I45c5e6710240685bf54b73b0d7a64271;
reg [MAX_SUM_WDTH_LONG-1:0]                I5827bc87b5db1801b7db16e1e61515db;
reg [MAX_SUM_WDTH_LONG-1:0]                I1c85c8f73ef80a6808c6aec0c8eca8ab;
reg     [5-1:0]          Id88b9265ff08e0730e6a41abe1f80a32;
reg [MAX_SUM_WDTH_LONG-1:0]                Id13c99b7f7500c8195b54627efbc4232;
reg [MAX_SUM_WDTH_LONG-1:0]                I4636821315d702a677dc93113872e647;
reg [MAX_SUM_WDTH_LONG-1:0]                I9c981b0614a29386ca5e8ebc06a17f15;
reg [MAX_SUM_WDTH_LONG-1:0]                I4df3d4dac24877b14e6d361bafc1a800;
reg [MAX_SUM_WDTH_LONG-1:0]                I913d818403024510c55b65b56a38dd89;
reg     [5-1:0]          I6330943c9295298c53e889d47c7904d9;
reg [MAX_SUM_WDTH_LONG-1:0]                I57015930f5b09a6c6b030ed01dad2177;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib54d55a70605119e37e9898b940ff636;
reg [MAX_SUM_WDTH_LONG-1:0]                If7e146da4f3bd255b8457fd6902005f6;
reg [MAX_SUM_WDTH_LONG-1:0]                Ied00d87af99ae55144fdde41ebfc1357;
reg [MAX_SUM_WDTH_LONG-1:0]                I7774313f1ae5a2de98855aad572b3676;
reg     [5-1:0]          I5686b595177e07dd5bf231a35ee41659;
reg [MAX_SUM_WDTH_LONG-1:0]                I679baea452c3c6d04c53baa88edd8eb3;
reg [MAX_SUM_WDTH_LONG-1:0]                If4132b39ddb92aa02d8d0346fb0e6691;
reg [MAX_SUM_WDTH_LONG-1:0]                Iba70e737d52e6812a67c159520e5192f;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib9ceb8315f0cd848f861bab677c2c694;
reg [MAX_SUM_WDTH_LONG-1:0]                I7846bc2cc11e08d05f7c853c4920d555;
reg     [5-1:0]          I9c0b88a0be66d62f8ab061aeaee7e60f;
reg [MAX_SUM_WDTH_LONG-1:0]                I0865623d3350645e63fa6e6c9b78ac57;
reg [MAX_SUM_WDTH_LONG-1:0]                I0262b30a4efa9f1cfb11d1c3940de9e7;
reg [MAX_SUM_WDTH_LONG-1:0]                I7a2e79d42779ad235bca6ce3757cf588;
reg [MAX_SUM_WDTH_LONG-1:0]                I09e9a3cd4c12d204f760758e873a177b;
reg [MAX_SUM_WDTH_LONG-1:0]                I30b0b1d54912c1a41a02a25ab238bb54;
reg     [5-1:0]          I9ef21ef20099af28d9a8c794f70d45a5;
reg [MAX_SUM_WDTH_LONG-1:0]                I49fb0909ddf66fc0073e6400f1a07844;
reg [MAX_SUM_WDTH_LONG-1:0]                I9938397dc94002481984f5b560fadc58;
reg [MAX_SUM_WDTH_LONG-1:0]                I4378d139db4b710e3587aa72df22b70d;
reg [MAX_SUM_WDTH_LONG-1:0]                Ifa43d74fa91b7b9884969f575ef9ca8e;
reg [MAX_SUM_WDTH_LONG-1:0]                I7c19a79f441ecbb73685db5a505e7479;
reg     [5-1:0]          Ic2941d16ae6a5cbce70e8546a18ca4ff;
reg [MAX_SUM_WDTH_LONG-1:0]                If2af8106efc1f7dd02c074af68278b3d;
reg [MAX_SUM_WDTH_LONG-1:0]                I89a3f8d5f760d1a650f85814cbfdc017;
reg [MAX_SUM_WDTH_LONG-1:0]                Ifae345c79662c3df3dff0fe68ad68746;
reg [MAX_SUM_WDTH_LONG-1:0]                I88a61cf72347d695489909d0819332ab;
reg [MAX_SUM_WDTH_LONG-1:0]                I9aaa036a6158d11c235bdc8406d79f4c;
reg     [5-1:0]          I8e29ebe9ee25ea8ef3e52ff56fc29157;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie8df350430970b5f1229cda772440f85;
reg [MAX_SUM_WDTH_LONG-1:0]                I7d77ac9b64b2e8cae21c6e36947e3ca2;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic1faed76fca5a9ceb7db26c2f43623d9;
reg [MAX_SUM_WDTH_LONG-1:0]                I3ca2b9b77ed8d78a10aff42a07a53b07;
reg [MAX_SUM_WDTH_LONG-1:0]                I1f00849ea055a7893df386aed162a7b6;
reg     [5-1:0]          Ic3742290179b27b9865f9d1f88d66266;
reg [MAX_SUM_WDTH_LONG-1:0]                Iaf8a19fde3de660c3fa925593bebbe0c;
reg [MAX_SUM_WDTH_LONG-1:0]                Icd1da43a4d95230e79dbd35a7ae41066;
reg [MAX_SUM_WDTH_LONG-1:0]                Ice9079fb6e08d629f8c0c9ce332c8f11;
reg [MAX_SUM_WDTH_LONG-1:0]                I15fafe2baba4d2f28037023a81ce0a81;
reg [MAX_SUM_WDTH_LONG-1:0]                If4d5b48882e9e628cf51ad2ac2f38c22;
reg     [14-1:0]          I04302edb2671c5bc0ca2673cd53935e1;
reg [MAX_SUM_WDTH_LONG-1:0]                Id0eef1adba01447c14a6f005782dd9a2;
reg [MAX_SUM_WDTH_LONG-1:0]                I1d1a7c5928982c278d068ebd262254da;
reg [MAX_SUM_WDTH_LONG-1:0]                I6354a0e638340378124e4df7f3d145b8;
reg [MAX_SUM_WDTH_LONG-1:0]                I0236c912c6d684bf4862b725be9d5951;
reg [MAX_SUM_WDTH_LONG-1:0]                I6f3be51d69b2b64a04e55b8946d5dd56;
reg [MAX_SUM_WDTH_LONG-1:0]                Icde3e6dbcf985682041f30903ad95572;
reg [MAX_SUM_WDTH_LONG-1:0]                I46ee30b46020d91707689f3468f00e26;
reg [MAX_SUM_WDTH_LONG-1:0]                I2605f078c1a9006c93855a9a2b0cf6b9;
reg [MAX_SUM_WDTH_LONG-1:0]                I4d226dd2f0bfcdbea6a2e6a6613c1b64;
reg [MAX_SUM_WDTH_LONG-1:0]                I5c942076b173cf527e1be2ddb8560e84;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic95191bccb18e26c10e56be395ca6b1a;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia284f974dd8a526f31eb81ed71a06e94;
reg [MAX_SUM_WDTH_LONG-1:0]                Icc93450a007cee4c0a42717ed7600528;
reg [MAX_SUM_WDTH_LONG-1:0]                I9ec9f389d0489908d497487e44c6edcd;
reg     [14-1:0]          I480a0f6d6c3eb936de10a72749f6cd3f;
reg [MAX_SUM_WDTH_LONG-1:0]                If8a527cc7f06a9963a80a880d225d34c;
reg [MAX_SUM_WDTH_LONG-1:0]                I39ff4663007dbc89b403f3b08a69bb6c;
reg [MAX_SUM_WDTH_LONG-1:0]                I9590eb28a81c730b83b92ef7653e71a1;
reg [MAX_SUM_WDTH_LONG-1:0]                I2ba1acca919bddcc22a41a28d43a4e3e;
reg [MAX_SUM_WDTH_LONG-1:0]                I62d8efd4227cb3dc88aa08b6585fafc8;
reg [MAX_SUM_WDTH_LONG-1:0]                I749e987266a20840bb8a4b1a2a2fc5b0;
reg [MAX_SUM_WDTH_LONG-1:0]                I7607af5d98e8070e3d15cee23cdf877e;
reg [MAX_SUM_WDTH_LONG-1:0]                I2e11a697d7f17ac30302eadb500de72d;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia0886ce792e062e22d0c224158cdfb7d;
reg [MAX_SUM_WDTH_LONG-1:0]                I6b3cd79aa87235ff174c0299b855dd3d;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie4ae993ddb776bdffec843db0def2f5c;
reg [MAX_SUM_WDTH_LONG-1:0]                I3ed2da9b53daac0852a06ad1acfad21b;
reg [MAX_SUM_WDTH_LONG-1:0]                Idefa29d4d4e2a6e9147f84893520096f;
reg [MAX_SUM_WDTH_LONG-1:0]                Id1fbbe0594dae272856566522633bb3d;
reg     [14-1:0]          I50976b0051e84b6a42fc1dbabd7d20ae;
reg [MAX_SUM_WDTH_LONG-1:0]                I8070a3b7d8b1a7ae90c1a2d27aed09aa;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie88285ce2b9c71de02ebd62e8f44ca72;
reg [MAX_SUM_WDTH_LONG-1:0]                Ica1997c6c569c1d1f45224fbaa4e6b59;
reg [MAX_SUM_WDTH_LONG-1:0]                Iaf08bcaaeb15bb0c971432f7f8b16d0a;
reg [MAX_SUM_WDTH_LONG-1:0]                Idcb37cfc357cc088c775409fb9225b51;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic419255414995e7168afb97b051fa64f;
reg [MAX_SUM_WDTH_LONG-1:0]                Iee6da3120d73373627b25ab7c0dedd28;
reg [MAX_SUM_WDTH_LONG-1:0]                I56fc99a22960232b305d6e683c66fcc7;
reg [MAX_SUM_WDTH_LONG-1:0]                I0a9a09b0ab43d2a0f1d1d01e13f0333c;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibc73d07e0c97a6fcae791e04106cb082;
reg [MAX_SUM_WDTH_LONG-1:0]                I224bbdf94ac86c5c376d1db4f4d4e060;
reg [MAX_SUM_WDTH_LONG-1:0]                I43f2b69c6b427de3095c44d4166b77cd;
reg [MAX_SUM_WDTH_LONG-1:0]                I1e50c90010a3df1a8ce1cff811cc7a0c;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie1817cbf3a80dae435a5571dfbd2f5ad;
reg     [14-1:0]          I82e0e091fba6f79cef97eacac4b43ecb;
reg [MAX_SUM_WDTH_LONG-1:0]                I0052d562fb3182890c8828e52d437b11;
reg [MAX_SUM_WDTH_LONG-1:0]                I1eedecb1d8ff505c75be7787199afada;
reg [MAX_SUM_WDTH_LONG-1:0]                I7ef544597a185b1de63b4ffc4a1d44c2;
reg [MAX_SUM_WDTH_LONG-1:0]                Iadeedf3870f0b1eae98d0f7dbbeff04a;
reg [MAX_SUM_WDTH_LONG-1:0]                I70ae07db9b44d530be220f06401d3d3d;
reg [MAX_SUM_WDTH_LONG-1:0]                I7992ea31927b4f0e268462a3b0f18c5d;
reg [MAX_SUM_WDTH_LONG-1:0]                Iadf927d18644a232ad1f1eba7db82934;
reg [MAX_SUM_WDTH_LONG-1:0]                I2a9c673cdd7ded79e09ada38c0f47e6f;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia86740e870d8063f0266b68ad6d7481d;
reg [MAX_SUM_WDTH_LONG-1:0]                I6627bcdbaa8afb115123777abd45435b;
reg [MAX_SUM_WDTH_LONG-1:0]                I96fe3eb633eff6958ac575b997460bb9;
reg [MAX_SUM_WDTH_LONG-1:0]                Iefdcb71f2903b11f5cb0b8857f7a1727;
reg [MAX_SUM_WDTH_LONG-1:0]                I2eb90278aaa54b9c8212b3b4af7c3617;
reg [MAX_SUM_WDTH_LONG-1:0]                I43493f70f0336453d77caf7f27503daa;
reg     [7-1:0]          I3d50cfeaa4b69c09bb648b8873a6bc24;
reg [MAX_SUM_WDTH_LONG-1:0]                I26a7fe395eb583258c1ac58aaaa3234a;
reg [MAX_SUM_WDTH_LONG-1:0]                I21668ff77cf75570cae97f575cbcf644;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie48be9e6b6fd63baa104d0a6a4561a1a;
reg [MAX_SUM_WDTH_LONG-1:0]                I05370777439b01811fe7f750d2f724f4;
reg [MAX_SUM_WDTH_LONG-1:0]                Icdcd83341f6b5c404f91ec7e97d0550c;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibba4e82d1510ddc16eb4ef64893cec02;
reg [MAX_SUM_WDTH_LONG-1:0]                Ifb00ae47340bc99669c71da34cccc59e;
reg     [7-1:0]          I33a6ffad80ddf99a4d316a049078244d;
reg [MAX_SUM_WDTH_LONG-1:0]                I75a4cf2948bebc58e12bb039ed273ff2;
reg [MAX_SUM_WDTH_LONG-1:0]                I5a9fdec7d7ff99fe33ad6cd8afd9e059;
reg [MAX_SUM_WDTH_LONG-1:0]                I47b1695a74e4d27389b97543415dcc67;
reg [MAX_SUM_WDTH_LONG-1:0]                Ieb38fa62119a5a77c060d6634e051298;
reg [MAX_SUM_WDTH_LONG-1:0]                I3459d98131faef5a5040a03847890b55;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie9b9221b2122087cd5f309570b6d31ca;
reg [MAX_SUM_WDTH_LONG-1:0]                Id4451722e8e2393d627dcd0175dc9903;
reg     [7-1:0]          I980165c1147ac5ff86619c841c6031dc;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic10356f9069e3651b9c045c906e63512;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic3a431f39c678b7175ed30fde1fa6424;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib01cfd833a63500e03333f263805db3d;
reg [MAX_SUM_WDTH_LONG-1:0]                I0b7b4c0a8503c751229edfe0237cc903;
reg [MAX_SUM_WDTH_LONG-1:0]                Iace01234164c8a9f7c98eeb83268745b;
reg [MAX_SUM_WDTH_LONG-1:0]                Iace8b3b3a4c16763132b5aaa6b24212d;
reg [MAX_SUM_WDTH_LONG-1:0]                I80a89644e278e96b1cd1c4b7f764dc34;
reg     [7-1:0]          I19df055705f322292a3601fa63f0e5f9;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia92d2276a8a23521ad1b88df7c27bc2e;
reg [MAX_SUM_WDTH_LONG-1:0]                I39bbec42c442d1e8c818f46ad9c096a8;
reg [MAX_SUM_WDTH_LONG-1:0]                I88f1b5c12759a5efb2d2ded8483c9ed2;
reg [MAX_SUM_WDTH_LONG-1:0]                Iaf4ae293c576af16f5f43a8b86c1aa3d;
reg [MAX_SUM_WDTH_LONG-1:0]                I68b575fcbc5321d4d26a22bcdbb506f6;
reg [MAX_SUM_WDTH_LONG-1:0]                Idf600b93ee1018ecf969ed7944b6bc7b;
reg [MAX_SUM_WDTH_LONG-1:0]                I1cd93172cf5996bc870063aa642188a2;
reg     [13-1:0]          I0e0b15868b02ca52b260f17f150d237e;
reg [MAX_SUM_WDTH_LONG-1:0]                I4af080cb4e5cc525db95e5f401019e8c;
reg [MAX_SUM_WDTH_LONG-1:0]                I6fc8044eb226a14ff1a786ddc96d2414;
reg [MAX_SUM_WDTH_LONG-1:0]                I27fd0073dbcdee599fbe85cf48806efc;
reg [MAX_SUM_WDTH_LONG-1:0]                Iaee6d725a8b2653eeac6d5acb91f8f36;
reg [MAX_SUM_WDTH_LONG-1:0]                I4afdeba4fc2a12a6cbe3567a519367fc;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib42816335dd8475dcc78662c4c0786c1;
reg [MAX_SUM_WDTH_LONG-1:0]                I343c9efe71164c01e9c7d599e032864a;
reg [MAX_SUM_WDTH_LONG-1:0]                I108c269ceec4adcff9afeda01101b838;
reg [MAX_SUM_WDTH_LONG-1:0]                I761983331fb6e3c6c437b3f1660f0b6b;
reg [MAX_SUM_WDTH_LONG-1:0]                I70d32affde22f9dcb2d77430fca39069;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic08e85346f61da036a15345a13ac12f0;
reg [MAX_SUM_WDTH_LONG-1:0]                If5dfdadb3868ed5a495007362f7db648;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia1ee5579358b564de06c08ca418a9bf4;
reg     [13-1:0]          I3c0b6f53f0a5cda5b6758b2ee2c83b92;
reg [MAX_SUM_WDTH_LONG-1:0]                I9bb81dda8102b829441be46460eb8900;
reg [MAX_SUM_WDTH_LONG-1:0]                I8eef6ca0a61a21882ea28b3d63735228;
reg [MAX_SUM_WDTH_LONG-1:0]                I438522d92cce6f7010246424746ca255;
reg [MAX_SUM_WDTH_LONG-1:0]                I92496f68b44a94565af28a2c28d6fbae;
reg [MAX_SUM_WDTH_LONG-1:0]                I66528f43f614f0edb715564eba3c77c1;
reg [MAX_SUM_WDTH_LONG-1:0]                I8cab9fba615b94fd4bb6934325be8ab8;
reg [MAX_SUM_WDTH_LONG-1:0]                I92d9fec22d36b1baac8bd78abfc1bbd5;
reg [MAX_SUM_WDTH_LONG-1:0]                I4eadce87f47df6d8f0e4acd057de5a09;
reg [MAX_SUM_WDTH_LONG-1:0]                I73203143fe37933c16fff873c1abf512;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibed2a63af723a7abf96dacf1951e5266;
reg [MAX_SUM_WDTH_LONG-1:0]                Id667c80003b5541de9f84d3b8709c828;
reg [MAX_SUM_WDTH_LONG-1:0]                I02cbb4255db2b21ea32140f9e9ddb36b;
reg [MAX_SUM_WDTH_LONG-1:0]                I65354f2069de0c25bbe7cd50fbe892aa;
reg     [13-1:0]          I8e591d83170c8ba46d31c61935311b22;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic279867ebf3055980f3d813d5dc8dec6;
reg [MAX_SUM_WDTH_LONG-1:0]                I5c05da8a222ad5effb9815cbf3ec25f3;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib8bf21f32c0e8b9cfa42a53807bfe3a3;
reg [MAX_SUM_WDTH_LONG-1:0]                I7208256bb198bfce1be71390b01bc028;
reg [MAX_SUM_WDTH_LONG-1:0]                I49f2a06ceb3a59773c65b19f54ff362b;
reg [MAX_SUM_WDTH_LONG-1:0]                I86e495dc894d2aace15c1aff89798bf7;
reg [MAX_SUM_WDTH_LONG-1:0]                I0d53bb5344cabe5fa5ce3ecf7122a260;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib2f5f5fc77ea8b529f2471c54388f2d1;
reg [MAX_SUM_WDTH_LONG-1:0]                Idcada1bfb3c0d1f2a09aab58a2071a57;
reg [MAX_SUM_WDTH_LONG-1:0]                I814b62120953991f9da055f118967e05;
reg [MAX_SUM_WDTH_LONG-1:0]                I123a212546a8ac394051425db4924812;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie95f1a7e0effcec0aa423dc803056a13;
reg [MAX_SUM_WDTH_LONG-1:0]                I106deaff50b8480eac31ddbae2ec7c61;
reg     [13-1:0]          I02b62fafd371de339f299f8aefec6c43;
reg [MAX_SUM_WDTH_LONG-1:0]                I68528be9951f5b8805411711cd11ea59;
reg [MAX_SUM_WDTH_LONG-1:0]                I0f034a8f077b0ab231727b6298e366d8;
reg [MAX_SUM_WDTH_LONG-1:0]                If9c12f8662333fb54a45cfa1bc5da487;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie1681d905517daafcc7584725cd6014c;
reg [MAX_SUM_WDTH_LONG-1:0]                I2ff3edcdb6158f1e3c9a555aeefc0850;
reg [MAX_SUM_WDTH_LONG-1:0]                I43b380be6df7df0d354223d0a0d6d6b6;
reg [MAX_SUM_WDTH_LONG-1:0]                I23eb1dc4d1c992f804dd04a2d823c778;
reg [MAX_SUM_WDTH_LONG-1:0]                I7f90f96c0260560ad5e6dc7448b2670a;
reg [MAX_SUM_WDTH_LONG-1:0]                I07b417cdcc99eaea3413f563e26ddc73;
reg [MAX_SUM_WDTH_LONG-1:0]                I2f3ab9654e515a54e22e73d6c130ccc3;
reg [MAX_SUM_WDTH_LONG-1:0]                Iebdc41368d57498a04fa73e30b10a966;
reg [MAX_SUM_WDTH_LONG-1:0]                I5b4305bef5b4350c1d7ae143667afddd;
reg [MAX_SUM_WDTH_LONG-1:0]                I2795d21d343b83a69146314a2407cfa2;
reg     [6-1:0]          I6ebab438dc55ccf6c1600313891d9c38;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic6386d7d8813731d612e24b715740275;
reg [MAX_SUM_WDTH_LONG-1:0]                I4c366a57920ff090a98a2cb8b9caa00b;
reg [MAX_SUM_WDTH_LONG-1:0]                I14cf5d43fc9864820a8a25efcc5c6d86;
reg [MAX_SUM_WDTH_LONG-1:0]                I33b99994abbb5ecf8eed4de39033e4f8;
reg [MAX_SUM_WDTH_LONG-1:0]                I7c3291f0250d13ca94802b0b071a95c6;
reg [MAX_SUM_WDTH_LONG-1:0]                I2c926fd9d306e9ae13364e07c4b0395b;
reg     [6-1:0]          I2fbf89398a148c47810456812dbee5a6;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib23edc35fa5bbfe0415fcf0861a22d9b;
reg [MAX_SUM_WDTH_LONG-1:0]                I3e0e682047f7cc36142e668828cbff1e;
reg [MAX_SUM_WDTH_LONG-1:0]                I99fb9030e8361e57818c07511479a9b8;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic87c3d7762a18772972552162e1d1a8c;
reg [MAX_SUM_WDTH_LONG-1:0]                I7e393e6c1d1bc44daaab120d55f5dd59;
reg [MAX_SUM_WDTH_LONG-1:0]                I448f126fd3932d5065abbe7bb2d92c56;
reg     [6-1:0]          Icac5a9001ee113e612e3457b4b49ee68;
reg [MAX_SUM_WDTH_LONG-1:0]                Ifc8c6df8904b97674f2970ebc95b523c;
reg [MAX_SUM_WDTH_LONG-1:0]                Icd0622a90782b9c451950e7ab0399567;
reg [MAX_SUM_WDTH_LONG-1:0]                I6493b3c087d4685a6b3f98c73dc2ff49;
reg [MAX_SUM_WDTH_LONG-1:0]                I20c2057240417146df144b518b43d052;
reg [MAX_SUM_WDTH_LONG-1:0]                Ied029d0bdea3bf134744c99426fa72dc;
reg [MAX_SUM_WDTH_LONG-1:0]                Icb82c9ff4cb58159a1c3115c6fdd5f8c;
reg     [6-1:0]          I9461e92a5880cb9e04fcece2ef4674f0;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia3450e134e4086c35acbdee1e6042396;
reg [MAX_SUM_WDTH_LONG-1:0]                I5a0f27df5158309f32f0df31e8ae3ae3;
reg [MAX_SUM_WDTH_LONG-1:0]                I17d9e19854cef197fd3267618617efc3;
reg [MAX_SUM_WDTH_LONG-1:0]                I2993acb61f1abe529f8a60c94a438550;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic8be2c94235fb40f78da33179ce4873a;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib3367565e4456da15e7c2315dccdb5e4;
reg     [8-1:0]          I07930a807994815de45864af579902c4;
reg [MAX_SUM_WDTH_LONG-1:0]                I15a1671def323cd294591564ae6ef8b1;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic512effb493a06ece58a2af155135004;
reg [MAX_SUM_WDTH_LONG-1:0]                I2c72248cbe49ec0a0febac2437b8a6dc;
reg [MAX_SUM_WDTH_LONG-1:0]                I964e17c41a134c080e9c43412a514f3f;
reg [MAX_SUM_WDTH_LONG-1:0]                I94f1724740defe5bb7e40041d0e266a0;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic19486b6ab0373b9c0ad8f7597782d8f;
reg [MAX_SUM_WDTH_LONG-1:0]                I31243de90dc2a1656ca9d5e03bdd78da;
reg [MAX_SUM_WDTH_LONG-1:0]                I242a30bdc8699d8ff550b25dd53d6c59;
reg     [8-1:0]          I72a2f42b727a0503d43332c0f22d5ae3;
reg [MAX_SUM_WDTH_LONG-1:0]                I9d15f76bb68b214057566cba4b511214;
reg [MAX_SUM_WDTH_LONG-1:0]                I9cc16a00912e7dfc05fb505a9db23cd8;
reg [MAX_SUM_WDTH_LONG-1:0]                Iacf9640cbf486411d6ceb8fe1a2fd5c9;
reg [MAX_SUM_WDTH_LONG-1:0]                I9015033ab0caf3fa41dae4de43f24a82;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia630e59cbce82a570ae3890a6c0221e5;
reg [MAX_SUM_WDTH_LONG-1:0]                I4904ab14b19fa1b6befc218bc7be3842;
reg [MAX_SUM_WDTH_LONG-1:0]                I282d2eb4e74e034694e33273b9cb19d5;
reg [MAX_SUM_WDTH_LONG-1:0]                I3f33901c407a87e10d86c13c83dd52eb;
reg     [8-1:0]          I8b8b9c4777e6df3eb2b9313e69ef2c8c;
reg [MAX_SUM_WDTH_LONG-1:0]                I43f41bf07836cee48069e9890c1de2a0;
reg [MAX_SUM_WDTH_LONG-1:0]                Id88480a0a350bb5fcf01ed5fff0bbd4c;
reg [MAX_SUM_WDTH_LONG-1:0]                I1d9b9ff357667a362f0442f19986f451;
reg [MAX_SUM_WDTH_LONG-1:0]                Ice73589836da9028def6efb24a04dbbd;
reg [MAX_SUM_WDTH_LONG-1:0]                Idb72c046c5996fbbd80b706666ffbd92;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie5757e7b1647ab7d43cdbcf98cbb77fc;
reg [MAX_SUM_WDTH_LONG-1:0]                I6072331f838d82329a07a4ffa340c7b6;
reg [MAX_SUM_WDTH_LONG-1:0]                Idf6875955525d80dc660ce956f4a84e7;
reg     [8-1:0]          I4a16e8e7946d9a8220304fc1be3fb362;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia96955d9c0a8a587e0afab37c8415d8c;
reg [MAX_SUM_WDTH_LONG-1:0]                Ifec374bce7f5507438f550df22d61a01;
reg [MAX_SUM_WDTH_LONG-1:0]                Ief67e897e57b96e2ec200e82bbc7caeb;
reg [MAX_SUM_WDTH_LONG-1:0]                Ide604e9bbe35cb55892a4602e18b2527;
reg [MAX_SUM_WDTH_LONG-1:0]                I262f2390e77ec486ccd3a6ed05816e2d;
reg [MAX_SUM_WDTH_LONG-1:0]                I280e20c20c0b4f26278b3de9b2ff84e4;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib3a0307176d424a4733720416d71069d;
reg [MAX_SUM_WDTH_LONG-1:0]                I76060709de3ea188748849f043c59ac0;
reg     [9-1:0]          Ic2580cbeec8c11a19bd1e2ebc29d255e;
reg [MAX_SUM_WDTH_LONG-1:0]                I8be20605d26d218911e80a883a90d085;
reg [MAX_SUM_WDTH_LONG-1:0]                Ieafa9d74d4a61d28ac4a913db460bf33;
reg [MAX_SUM_WDTH_LONG-1:0]                I6fd1b4395af175eff85b3bfeef4c329b;
reg [MAX_SUM_WDTH_LONG-1:0]                I39e6d3fb468aa40ea73535e81556ea65;
reg [MAX_SUM_WDTH_LONG-1:0]                Iae449b74e50e0907feae9e60f2329426;
reg [MAX_SUM_WDTH_LONG-1:0]                Iebf769a6bdaf214c1006c55c608d4eda;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia030c08757123aae947f86ab8bfb6d94;
reg [MAX_SUM_WDTH_LONG-1:0]                I8c35c5b343b552c22000e194c517ca12;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibf80bb564263ea85bd886a8617f09bb2;
reg     [9-1:0]          If79ed5ee2b8710da0608c1e245d07d55;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib8dfd9b8badef282ca00a4f793c3c868;
reg [MAX_SUM_WDTH_LONG-1:0]                I596ad7e132f272cb196b74faa8c75aa4;
reg [MAX_SUM_WDTH_LONG-1:0]                Idc629414f6d0236ce0714cfaae23f065;
reg [MAX_SUM_WDTH_LONG-1:0]                I157fdf8775206858c08682db3039b084;
reg [MAX_SUM_WDTH_LONG-1:0]                Iacbb4daf5ce5c7eb1a2afe30d0cb5382;
reg [MAX_SUM_WDTH_LONG-1:0]                I4e08021c0235fafb60200aab97827a8f;
reg [MAX_SUM_WDTH_LONG-1:0]                I730634ea15ac94d241f3ad2d6393a227;
reg [MAX_SUM_WDTH_LONG-1:0]                Iee367c535d9c39f872d2ec043e7e7b33;
reg [MAX_SUM_WDTH_LONG-1:0]                I68bb1f26f878862f288c1f57049cf58b;
reg     [9-1:0]          I9497bbb4f746969a95cff948a3ee9ade;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia9b5d9ede006c56a6d83905529c77b7b;
reg [MAX_SUM_WDTH_LONG-1:0]                I1487170cb1f3370ad45efc801cefc8ab;
reg [MAX_SUM_WDTH_LONG-1:0]                Id88568dd34fbee42c9cb8cc15ac5c31d;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia30539545e66c4cfc16828140149180a;
reg [MAX_SUM_WDTH_LONG-1:0]                Icbfbb37bad6344005dd233b3605a784f;
reg [MAX_SUM_WDTH_LONG-1:0]                I91a6408a11fab36a8ba3dbd3f895a803;
reg [MAX_SUM_WDTH_LONG-1:0]                I47b878f27c30f79a37e97e022307e9e9;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie76b0739aec66f8860870e66e87a6445;
reg [MAX_SUM_WDTH_LONG-1:0]                I50383e3d7c172eedfa00aa50a9faac4c;
reg     [9-1:0]          I651d700a00d7004d8728bc7356f30926;
reg [MAX_SUM_WDTH_LONG-1:0]                Ifeaa99e03bda8ded058f98387de3d49d;
reg [MAX_SUM_WDTH_LONG-1:0]                I4255ac1af4367c321567c4e46b06ab25;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia445bdc7def7d8c1eec31ab892c25c41;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic3b4752136ac08e343933ccc3a4ec47c;
reg [MAX_SUM_WDTH_LONG-1:0]                Ica6707efd6d44ba6bbb87c0593a3d828;
reg [MAX_SUM_WDTH_LONG-1:0]                I739267bcc50c54b8a685cb3c6afc5cc1;
reg [MAX_SUM_WDTH_LONG-1:0]                I9160d11439c5140c0109b5190eb82e6b;
reg [MAX_SUM_WDTH_LONG-1:0]                I6ff7b86cd7f63f9243646f1be10b2577;
reg [MAX_SUM_WDTH_LONG-1:0]                I165653ab165cfafe2b74cd441331f9e1;
reg     [16-1:0]          I6f5c991e5fdcf56d582c6f80eb6731df;
reg [MAX_SUM_WDTH_LONG-1:0]                I08a8cd6965c23af6650568b654831b20;
reg [MAX_SUM_WDTH_LONG-1:0]                I9b6a674dbcbfcf65f1ae0deb8fc3566d;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie3a336de822ac7baf8486b1618ef1126;
reg [MAX_SUM_WDTH_LONG-1:0]                I5fc3c26d6c5aa893dfd5caa0f677233a;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie22b94121b58f17af14c75bfb27f96dd;
reg [MAX_SUM_WDTH_LONG-1:0]                I0d9f8c99194d9d6e187b4ad02fcce8b4;
reg [MAX_SUM_WDTH_LONG-1:0]                I71e101962e766a4d1484b3235359a4b5;
reg [MAX_SUM_WDTH_LONG-1:0]                If2539da6722562bbf31786fd0036666a;
reg [MAX_SUM_WDTH_LONG-1:0]                I22c8ccd4a9018ad1c129aa058bf579d8;
reg [MAX_SUM_WDTH_LONG-1:0]                I83330fef69470d2f5def8e6d7d9c50d2;
reg [MAX_SUM_WDTH_LONG-1:0]                I0539d598bbe3d50940329a282c801328;
reg [MAX_SUM_WDTH_LONG-1:0]                I202f88fdc946494d55fc8831c2e8a34c;
reg [MAX_SUM_WDTH_LONG-1:0]                I3ee10f6a7785a236db317515fdd23a2d;
reg [MAX_SUM_WDTH_LONG-1:0]                I453fdf4fbb5af5bd28a20d7643da9eb2;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic4a6c02880a9aead7353332708e3f388;
reg [MAX_SUM_WDTH_LONG-1:0]                I7fb3b66cb48521f8715f66bf5642cdb2;
reg     [16-1:0]          Ia5cc3055ba3365e64cf59c4d4fd3f093;
reg [MAX_SUM_WDTH_LONG-1:0]                I2fd872df07f50688486c0d602cfc5549;
reg [MAX_SUM_WDTH_LONG-1:0]                Iccefa45795486757515d95e5908b306a;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib1357cb20f471f1670ac2448f964f8eb;
reg [MAX_SUM_WDTH_LONG-1:0]                Iab953a8974a1eb619dc0f074c003b5f9;
reg [MAX_SUM_WDTH_LONG-1:0]                I6e37582849c2c98fd15ad92d22c222da;
reg [MAX_SUM_WDTH_LONG-1:0]                If004de0cac6e5f7701a1fce48c6936d5;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic1efa395cc1fd2c5a1d1559fb169a5a0;
reg [MAX_SUM_WDTH_LONG-1:0]                I8e96c69e7d872be23229353808c34953;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib6aded6c73a8cc3cb964b0ae895b859e;
reg [MAX_SUM_WDTH_LONG-1:0]                I939368b76d98b43826c68c7f468a5632;
reg [MAX_SUM_WDTH_LONG-1:0]                I544f6263f16cd5e0b7cf28c511a8f6e3;
reg [MAX_SUM_WDTH_LONG-1:0]                I484545c4d2c869d79eb17f51e11070a3;
reg [MAX_SUM_WDTH_LONG-1:0]                I39289e6385a9bc378a9b8dd440249a7f;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie9cce5746a83479a567bbaeac6dbf497;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic044d7419cc43736d278c2df33b4a3cc;
reg [MAX_SUM_WDTH_LONG-1:0]                I6714551e8885ef5e4490673fe1b2dad1;
reg     [16-1:0]          Iea7da1f43ba202d753b0edb0be8b3fcf;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie9ab3c88ac62369e3d92d110165a94a8;
reg [MAX_SUM_WDTH_LONG-1:0]                If38feb4f76f761dce6145731ad235d7f;
reg [MAX_SUM_WDTH_LONG-1:0]                I6359856a1843d8c8b65dc478bccb3acd;
reg [MAX_SUM_WDTH_LONG-1:0]                If6f3d91c3c7a43622b9a522492cd83d3;
reg [MAX_SUM_WDTH_LONG-1:0]                Id023a6298e65da1f4da3831f5136afc2;
reg [MAX_SUM_WDTH_LONG-1:0]                I6b24690f394792edb0d82b3b9e110851;
reg [MAX_SUM_WDTH_LONG-1:0]                I5b55c285f7e3e78447fee68532ab9f7f;
reg [MAX_SUM_WDTH_LONG-1:0]                I32701d9e4b96853c53f0ab651a6a4ba2;
reg [MAX_SUM_WDTH_LONG-1:0]                I82f266e5792cdb6e7ebd264e246161f5;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibfacfe5b83819afe7fbd4bffa2d6d4e2;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib8e68a77ad8b9e7cf415bee17645c3f9;
reg [MAX_SUM_WDTH_LONG-1:0]                I644ee0055a55f54ab3544bb532e39c61;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic5467e42aa377c6ffd8f70673808774f;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic57eb4a034247a4c952d8224ea9f2bac;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia642db613c0ec1ca4e69afde7a14a839;
reg [MAX_SUM_WDTH_LONG-1:0]                I432aa7cb844286c442356954f8814260;
reg     [16-1:0]          I872f61d20baf011e867b44dc5539fc37;
reg [MAX_SUM_WDTH_LONG-1:0]                If520c1cd27f9d4bc52d0d029f693b660;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie87075ac979410cc11099a356966b8a2;
reg [MAX_SUM_WDTH_LONG-1:0]                I6fab46b1766878b26b53f352fee98223;
reg [MAX_SUM_WDTH_LONG-1:0]                Ieaf14683f40374c4531326d228cb43c3;
reg [MAX_SUM_WDTH_LONG-1:0]                I5149125aaaad943d891df6a3c2be93a0;
reg [MAX_SUM_WDTH_LONG-1:0]                I770dff588ee1f52f58bea1921cb23383;
reg [MAX_SUM_WDTH_LONG-1:0]                I8f0a90e761111a613d2488285534a500;
reg [MAX_SUM_WDTH_LONG-1:0]                I765a8825e42180a6c63f7b33703bb483;
reg [MAX_SUM_WDTH_LONG-1:0]                I512cc8f6519aa08aee18225b56d47c9f;
reg [MAX_SUM_WDTH_LONG-1:0]                If08370fd0e8af818c6db20f43e74034d;
reg [MAX_SUM_WDTH_LONG-1:0]                I0ff382edfc8051459657ffa3899f5f73;
reg [MAX_SUM_WDTH_LONG-1:0]                I9d2864024148337277523ef7fa2e1600;
reg [MAX_SUM_WDTH_LONG-1:0]                I1c85a2d1df6749a194072eb731506bfe;
reg [MAX_SUM_WDTH_LONG-1:0]                I3e3ce8b4ead150a6eae2e5c701c7b598;
reg [MAX_SUM_WDTH_LONG-1:0]                I45bc13ae0e0554a79c62cd9c6aa8f2a5;
reg [MAX_SUM_WDTH_LONG-1:0]                I92678f5b52c9c55556ff7f17f0f607b7;
reg     [9-1:0]          Ieb244944e7ee8236a207924f56fbc689;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib4bdc9069d0c08655f5e87f705943eda;
reg [MAX_SUM_WDTH_LONG-1:0]                Idbf9094c94c931f16fba468b9dd59a25;
reg [MAX_SUM_WDTH_LONG-1:0]                I1c3c4ce44610e04c5eef2fcbc2ea5114;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie84be0ae8311d906eff08f7f5b214943;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic90b98708faa8c8b75d4bd9a52c292f7;
reg [MAX_SUM_WDTH_LONG-1:0]                I8eba6f14f42701d22859fbea94bd1871;
reg [MAX_SUM_WDTH_LONG-1:0]                I6d83efa9f988328f487e9232bf2633a2;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic23e01562c8a753fd70c343297be288a;
reg [MAX_SUM_WDTH_LONG-1:0]                I5669856f88f5e2c98f64df696db76414;
reg     [9-1:0]          Ie9b2be4c32334220e134e041ca8dfc06;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic3a608b850709286ea0ad2f67425d9ac;
reg [MAX_SUM_WDTH_LONG-1:0]                I5267fa34449e6eebe891017fc32d0749;
reg [MAX_SUM_WDTH_LONG-1:0]                I599d01cfe6e54d8e45d64446c446818d;
reg [MAX_SUM_WDTH_LONG-1:0]                I8f94dbafaac589ac9f14b56d4556ff96;
reg [MAX_SUM_WDTH_LONG-1:0]                I754563caea429d3d0e22df5d193b84eb;
reg [MAX_SUM_WDTH_LONG-1:0]                If7f373506cac70f8ba1222db135c27e8;
reg [MAX_SUM_WDTH_LONG-1:0]                I69f563e7b7ad483893ac9c4684349769;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia0a02781c674fe5d769206448d475245;
reg [MAX_SUM_WDTH_LONG-1:0]                I1b7a401bc11741e6f011fb9895b5c797;
reg     [9-1:0]          Id6f07dee3e47f39e3b43329c26f690f7;
reg [MAX_SUM_WDTH_LONG-1:0]                Ieb528d666fdb708279184bb59eac25d9;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic3ff7ce12c836bf0693252b9a7a7cfe8;
reg [MAX_SUM_WDTH_LONG-1:0]                I19bba6a58ad3ef959b33701f82761984;
reg [MAX_SUM_WDTH_LONG-1:0]                I8acc93b34974c1e708b0e1591f7b2d3d;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib60d4ac0fcadcdfce5a14fb92f58423f;
reg [MAX_SUM_WDTH_LONG-1:0]                I039f05d5be891a37e04556f1eae674d2;
reg [MAX_SUM_WDTH_LONG-1:0]                Id0f75e19b94541ed5c5c352d13390d2d;
reg [MAX_SUM_WDTH_LONG-1:0]                Ife1190f76c2e251704c2960c23330a48;
reg [MAX_SUM_WDTH_LONG-1:0]                Id3e0c98bff2636e216b4d3a0ffd51054;
reg     [9-1:0]          Ic7f04c065f8ff82c2288f1de77d37189;
reg [MAX_SUM_WDTH_LONG-1:0]                If4d3b31b87c0f723241d35ce7e854eba;
reg [MAX_SUM_WDTH_LONG-1:0]                I72369dedfe36cb22269033cc305b730c;
reg [MAX_SUM_WDTH_LONG-1:0]                Iec71fe7fcebccf1ae0d10a5d187fcc44;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie11da10808c4ca84f399535df6261307;
reg [MAX_SUM_WDTH_LONG-1:0]                I280fa9d114e227cd649bf0e55e845651;
reg [MAX_SUM_WDTH_LONG-1:0]                I94c4e11670b4233fa072517a8f19c901;
reg [MAX_SUM_WDTH_LONG-1:0]                I4dca2dd40a7127ce44f83b430a34c738;
reg [MAX_SUM_WDTH_LONG-1:0]                I1a24e98165afa62bd14986911a36fb6e;
reg [MAX_SUM_WDTH_LONG-1:0]                Ife1164cad7cda4aa9a08d94dfe86add6;
reg     [12-1:0]          I4267622319ca65909a3b40484dc74d3a;
reg [MAX_SUM_WDTH_LONG-1:0]                I8d8d95ff26f33f69a182b32ccde23905;
reg [MAX_SUM_WDTH_LONG-1:0]                I2508854bcbab37bd09c9465c377c06aa;
reg [MAX_SUM_WDTH_LONG-1:0]                I140078292f7209eccacd53a8bab18016;
reg [MAX_SUM_WDTH_LONG-1:0]                I141fb1cbe09f9abe282cffd4de815d25;
reg [MAX_SUM_WDTH_LONG-1:0]                If79d1d378f7c6fd29fc3335ec5f5c51d;
reg [MAX_SUM_WDTH_LONG-1:0]                I4a41999cea9357a85c73a0af509eeac9;
reg [MAX_SUM_WDTH_LONG-1:0]                I8e517c401d62dbb10dcc96ab536f6afb;
reg [MAX_SUM_WDTH_LONG-1:0]                I8ad3627f171eadcc960a688ac0afcbc0;
reg [MAX_SUM_WDTH_LONG-1:0]                I85c4d3d6c8408c6f38741257ed177ca6;
reg [MAX_SUM_WDTH_LONG-1:0]                Id66c47fd69c175a4393e975a269cf053;
reg [MAX_SUM_WDTH_LONG-1:0]                I37dca40506d61bdeab1255ed4892ca20;
reg [MAX_SUM_WDTH_LONG-1:0]                I340c98b886123c541a1b8d9fc8a6d48c;
reg     [12-1:0]          Iedd7d4ea8d082b40244c04946dfb14a0;
reg [MAX_SUM_WDTH_LONG-1:0]                I2dc64c3b06588542b027f997437bee63;
reg [MAX_SUM_WDTH_LONG-1:0]                Id92a37c091100e9df08e24498ecb4022;
reg [MAX_SUM_WDTH_LONG-1:0]                I74a4b9365391fd20c34588002ad40547;
reg [MAX_SUM_WDTH_LONG-1:0]                I461195b7ae78743e09ee50486ad6ebe5;
reg [MAX_SUM_WDTH_LONG-1:0]                I356d747600182675699a2d2634d4c5ce;
reg [MAX_SUM_WDTH_LONG-1:0]                I87d6a5d30c3e4202cf51f33c7a770c51;
reg [MAX_SUM_WDTH_LONG-1:0]                I960768a84aec9d5b8bc7c1c523024a25;
reg [MAX_SUM_WDTH_LONG-1:0]                I09b5273bb15d48a7fd78559930fa6d1c;
reg [MAX_SUM_WDTH_LONG-1:0]                I5814a85c45fd0f7be21ed325235fe4b7;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib06b60cf9933dd8952206c5f3ccced8e;
reg [MAX_SUM_WDTH_LONG-1:0]                I67347c413b5efd8ff9e0d5bc7ab2a047;
reg [MAX_SUM_WDTH_LONG-1:0]                I72b1bb104bf2843f161448baf7aab44b;
reg     [12-1:0]          I56e1fe0c7a62589c123876f2b4e57a26;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib23d889edb5a6d9f27de977d3b1a2616;
reg [MAX_SUM_WDTH_LONG-1:0]                Ifaff9dd032cf96487be819c59b03000a;
reg [MAX_SUM_WDTH_LONG-1:0]                I028ce03be0618b816e0ecdf43d4cd6e6;
reg [MAX_SUM_WDTH_LONG-1:0]                I6ae2523095237282533e0b5f1c26b488;
reg [MAX_SUM_WDTH_LONG-1:0]                I5aba6218461e8d571be03a3ef041ebaa;
reg [MAX_SUM_WDTH_LONG-1:0]                I6ca8a1fa2c72b1c61d11dc7d1ba5f37b;
reg [MAX_SUM_WDTH_LONG-1:0]                I3ec5819176ad4b0895a9118d90ab22b5;
reg [MAX_SUM_WDTH_LONG-1:0]                I49b64469d298012dbb131d879bff38d6;
reg [MAX_SUM_WDTH_LONG-1:0]                I95361d5f524ccb9feb42811af5c482e2;
reg [MAX_SUM_WDTH_LONG-1:0]                I9c4b34b5fb1d59c132bcaeb6258675df;
reg [MAX_SUM_WDTH_LONG-1:0]                I613d4b1e3b9e812b785c9cf14fefdfe6;
reg [MAX_SUM_WDTH_LONG-1:0]                I848ed394bd4f0b199d11c0ff458394a7;
reg     [12-1:0]          Ia8a468877c9f96713c8141df9205f92a;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie65a0634454381e24bb3223a333e3ad0;
reg [MAX_SUM_WDTH_LONG-1:0]                Iad166146f7df5e8068fc6efe4d3e4141;
reg [MAX_SUM_WDTH_LONG-1:0]                I63e45abd4d27219bddcef06108b72021;
reg [MAX_SUM_WDTH_LONG-1:0]                Id1bacd13718f7c29c26b63c239d04dd8;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia3104c69fb4f7abfb5efa3874169a7ad;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie1b7257c99831ec5864f65958ecf14fb;
reg [MAX_SUM_WDTH_LONG-1:0]                I4accbad1b451ed2b622e15ef9ae16d13;
reg [MAX_SUM_WDTH_LONG-1:0]                I5ce8b2f633011e89356243a1a71edeb6;
reg [MAX_SUM_WDTH_LONG-1:0]                I3e5139f24e3d082eb31b0e61ea9fa1aa;
reg [MAX_SUM_WDTH_LONG-1:0]                I61cc8a0f49e393721a62a776e4793deb;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie631e40caade823a196370fc3358f042;
reg [MAX_SUM_WDTH_LONG-1:0]                I4c971e714427664c59c6371e14781bae;
reg     [1-1:0]          Ida6059c6e0890f730536f97dfb83770b;
reg [MAX_SUM_WDTH_LONG-1:0]                I36ca732e811d67cd742d24fd4cae887b;
reg     [1-1:0]          I1993c1ed200d7cdf838d23c72a0c1c0b;
reg [MAX_SUM_WDTH_LONG-1:0]                I354fdd241d5d07f0d8380fe8924e0a8c;
reg     [1-1:0]          I07e04e352df9aa1988ccf05d9cb2d1d7;
reg [MAX_SUM_WDTH_LONG-1:0]                Id38b705f5d2863a020a475ffffc8afd6;
reg     [1-1:0]          Ic4c0ebcc3711c9844a3aa3875483d2f7;
reg [MAX_SUM_WDTH_LONG-1:0]                Id6e5d67e7bb7c4b999459374ea80459a;
reg     [1-1:0]          I28e344560ba76bb3b76d01d8c53693a9;
reg [MAX_SUM_WDTH_LONG-1:0]                I05341013abd4206eb66fcddfd63bfe26;
reg     [1-1:0]          I0600def6e6caada88ba6dedbb0d322ac;
reg [MAX_SUM_WDTH_LONG-1:0]                I15da71a21f5842cb65b543d9bc3e267b;
reg     [1-1:0]          Iddbf50612c89b5b95a5c9efb5575cae3;
reg [MAX_SUM_WDTH_LONG-1:0]                Iccf255fb3422c558465e45226068a16d;
reg     [1-1:0]          Iadc8f7f87b50bfff53d2d12d82489829;
reg [MAX_SUM_WDTH_LONG-1:0]                I1c2674b2e6b269ed539827412c5199a5;
reg     [1-1:0]          I53a658b443200b9f11f1830547b5f42d;
reg [MAX_SUM_WDTH_LONG-1:0]                I6a3f405bb4a0c4448d9b9d3dd95d036c;
reg     [1-1:0]          I170f424df45651abe215ec74d649a9eb;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib528bb7a64cce4f694081d151fa6fa86;
reg     [1-1:0]          I3c897bfed190017a876c44fd73a7ecea;
reg [MAX_SUM_WDTH_LONG-1:0]                Iaa40bd3abf668a21e0f87c7bda7b3f69;
reg     [1-1:0]          Iaecbbae967be2c62cacf2fa7f9801899;
reg [MAX_SUM_WDTH_LONG-1:0]                I919d36a7f6ad42c4bbc23222beb73106;
reg     [1-1:0]          I52f867f1009f2e8d18b50a777942bde3;
reg [MAX_SUM_WDTH_LONG-1:0]                I648d2a279dd1f587b1e45eeb35f2fa90;
reg     [1-1:0]          I56a39a0c67b1de0a3cab6c61af3eebcf;
reg [MAX_SUM_WDTH_LONG-1:0]                I194a64bef92ecf6714141eaa5d41c9d4;
reg     [1-1:0]          I490a65b3f7b30540906262ec5e12717b;
reg [MAX_SUM_WDTH_LONG-1:0]                Id332e7f482524adeac7f7cdafcf5ca46;
reg     [1-1:0]          Ib3c52fef8251d95e9abc8df0aad45d4e;
reg [MAX_SUM_WDTH_LONG-1:0]                I226383d68f89db716cfd8d08b837865a;
reg     [1-1:0]          If75725e534dcb00364d73a42769539fb;
reg [MAX_SUM_WDTH_LONG-1:0]                I2bdf5d319ba9089a4da34b108f5c5ae5;
reg     [1-1:0]          I9ddc427eef437ecc3ac4a2cf52aad4c3;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia91800792941ec7cc60415c3f844e4ed;
reg     [1-1:0]          I8999ca1f2fe9d4a30bd38fcb0daad2a4;
reg [MAX_SUM_WDTH_LONG-1:0]                Id7c507d96098ee7a955af8a48ee5d72a;
reg     [1-1:0]          Ie11cf6677812bb739255b053a9c9cd56;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie15e4c1bcdb0e18085d4b320ac6a925c;
reg     [1-1:0]          Iacc1d5a5c7811f0c9326ef80d1154fbb;
reg [MAX_SUM_WDTH_LONG-1:0]                I5485d9edcafc6202f6e5f0969979802f;
reg     [1-1:0]          I0efdadfd49c035a49d92243391395bca;
reg [MAX_SUM_WDTH_LONG-1:0]                I7fe364f9f537cbef782e7007848a1c10;
reg     [1-1:0]          Ie34d59bc77e06807937fe6f6860527e9;
reg [MAX_SUM_WDTH_LONG-1:0]                I52dcf5bace9cadcf8a895aaa6a8c1da8;
reg     [1-1:0]          I9661cb126908d8550b585e2bad383bd6;
reg [MAX_SUM_WDTH_LONG-1:0]                I13a9eec6175e695ab8bc4516cf57d6ec;
reg     [1-1:0]          Ic0b832fbcbdb57745fefcc1ac1438808;
reg [MAX_SUM_WDTH_LONG-1:0]                Iee73a7c685a4cee03f33d3ef379b1c8a;
reg     [1-1:0]          I2afd96714b26f30483c3935c2a68e64f;
reg [MAX_SUM_WDTH_LONG-1:0]                I740dc91716e3906ad078e2c7cc3c925a;
reg     [1-1:0]          Id6d4165b752630a1ce7ceb77fdcee477;
reg [MAX_SUM_WDTH_LONG-1:0]                I514d2dc697e9b39ba027c418a6df6cb9;
reg     [1-1:0]          I59baaf1ad22721cde9064b8aad65ac76;
reg [MAX_SUM_WDTH_LONG-1:0]                I782726e317a2aada9e755bcbc4b0d3fa;
reg     [1-1:0]          I9094f4e9c5b60add3acee212118a1dfa;
reg [MAX_SUM_WDTH_LONG-1:0]                I11eb26cf0f0b3a334e8f7317bf8d9eb0;
reg     [1-1:0]          I13168bab2231ed22a3509142f990e408;
reg [MAX_SUM_WDTH_LONG-1:0]                I26cb63ba20245b2c332b09e25c4409aa;
reg     [1-1:0]          I280145f996e5e249788cacca7caf0095;
reg [MAX_SUM_WDTH_LONG-1:0]                Idd7691d31f8d0c09ee988116d574ec59;
reg     [1-1:0]          Ia9db6d176e9b9579a1aa5f257cd1a9f6;
reg [MAX_SUM_WDTH_LONG-1:0]                Iecc02842a2d2b9b9e8187f2d39e62e05;
reg     [1-1:0]          I0ed43cf9eec83545457c57cfb6181d3c;
reg [MAX_SUM_WDTH_LONG-1:0]                I5551342f1751fc64f32744a46b9649be;
reg     [1-1:0]          I5b74f5fc705a0406ff2376cb8ac11db4;
reg [MAX_SUM_WDTH_LONG-1:0]                Iff7c29299f005c1cd5a16b64601e727e;
reg     [1-1:0]          I14f0d3ad4fec9ca492d6b36eb29a5dea;
reg [MAX_SUM_WDTH_LONG-1:0]                I17a5446e942bcc1dc2c96930e0a87a70;
reg     [1-1:0]          I3a25c80d9bf7655f4ce70cf29843db43;
reg [MAX_SUM_WDTH_LONG-1:0]                I719b67f84e07e90dfd29a8cd5d94cf39;
reg     [1-1:0]          I260dc9154b3a9fe38b0948e807bdb42d;
reg [MAX_SUM_WDTH_LONG-1:0]                I2c835dfb3596b8bf057a7cc21122c81f;
reg     [1-1:0]          Ic49b2c150e2face8c362e33f2d87f9c4;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib71b3d357c98dcdfae5c777ca3082275;
reg     [1-1:0]          I714350b3b56a3249aad06d5f59fbb291;
reg [MAX_SUM_WDTH_LONG-1:0]                I086bf19f620c8a8f6888e775cb1ed7f4;
reg     [1-1:0]          Ia318eb500b8bd71048bde375c1db65a6;
reg [MAX_SUM_WDTH_LONG-1:0]                I802c554d5b04af6b949677819a4966ed;
reg     [1-1:0]          Ia2c4192b1e4f180402550aebcf1dcd1f;
reg [MAX_SUM_WDTH_LONG-1:0]                Iceefb06cb3715e1b41e6f7d89420e5ba;
reg     [1-1:0]          I1686a95674ecad0c4e234b8aa6e22dd9;
reg [MAX_SUM_WDTH_LONG-1:0]                I56948bc48c0220893d68004615a6ebaa;
reg     [1-1:0]          I5ee21680396395f8338477fa2bb314ec;
reg [MAX_SUM_WDTH_LONG-1:0]                Iec1368f034655d61354ab5b5e94d7d89;
reg     [1-1:0]          I005e89f0a9a9a52aec92752813a70f81;
reg [MAX_SUM_WDTH_LONG-1:0]                I1e43c0aeeb8a2461d208eba24967af30;
reg     [1-1:0]          I0daca3ad02a67285295cd9fc330d8027;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia6eb85b127cf9c1a437611556296b967;
reg     [1-1:0]          I0d2ddde9edfef483482e6c177a084f6e;
reg [MAX_SUM_WDTH_LONG-1:0]                Ieba89aa901e61218074af53a2484a74b;
reg     [1-1:0]          I932ad562b582e2c9795f241c82901188;
reg [MAX_SUM_WDTH_LONG-1:0]                I8b3b875c6c07bd97ba598a5139156fa4;
reg     [1-1:0]          Ifee4aa12e36833c935c54ef27b1917da;
reg [MAX_SUM_WDTH_LONG-1:0]                I7b33ddad346077928620344542b9481e;
reg     [1-1:0]          I51e5b79f738795719ac21c6a88711a01;
reg [MAX_SUM_WDTH_LONG-1:0]                I11d967a5c5d14c88b5587d4cfed1d05f;
reg     [1-1:0]          I4e41e628a8af629421544cb4c6f45265;
reg [MAX_SUM_WDTH_LONG-1:0]                I27458d76b3ac6520fb379405c6b2956f;
reg     [1-1:0]          I9b2ec7db66661f7c9d85cfb1bc41893b;
reg [MAX_SUM_WDTH_LONG-1:0]                I2525111a2fb5f10d64bbd16e148653b8;
reg     [1-1:0]          I0a594a36728c7ac6244c504b8ea9c9af;
reg [MAX_SUM_WDTH_LONG-1:0]                I7b7cbcd1c6d2a2eeaaff474536a69eed;
reg     [1-1:0]          Ibd943ebf64fe56a1818d2bb8b9f9f8bd;
reg [MAX_SUM_WDTH_LONG-1:0]                Id2a7f0781d18dccc7c4e0b383b7cddfa;
reg     [1-1:0]          I8c3ba90c84f9375001e727b711dead8d;
reg [MAX_SUM_WDTH_LONG-1:0]                If8bc141d98ebe1be7fa81cde5c65868e;
reg     [1-1:0]          I387ca23d0e2183522ab041ec48bffef4;
reg [MAX_SUM_WDTH_LONG-1:0]                I8645e1326c66f5efef4b9c923599d1a3;
reg     [1-1:0]          Ib933575f5224d414f87bc71fa7498534;
reg [MAX_SUM_WDTH_LONG-1:0]                I0426ef66185128dd1ef4dbb68dcda585;
reg     [1-1:0]          Ibfe1bddf32fa63ea87c68de7a3af1815;
reg [MAX_SUM_WDTH_LONG-1:0]                Iddd954df5bae9b4240e0512f746669a9;
reg     [1-1:0]          I719c50f9bbc66decebe794fe6ea017dd;
reg [MAX_SUM_WDTH_LONG-1:0]                I29e940970d87e8e09b26ab1b0b8f2286;
reg     [1-1:0]          I833b0433a33dac70cb215bc8cc9f4863;
reg [MAX_SUM_WDTH_LONG-1:0]                I488f6d9676aa85a55d030bf12e8997a7;
reg     [1-1:0]          I9769761eb863e3273f9253ace4c69585;
reg [MAX_SUM_WDTH_LONG-1:0]                I99d761b75ade1fb2e8afbb1a77752609;
reg     [1-1:0]          I1fc63f388d047207a9375842c85e87f7;
reg [MAX_SUM_WDTH_LONG-1:0]                Iac4e3d20178049f9c59abf374752dccc;
reg     [1-1:0]          I414c4d389ecc00197f2138eff0b6454e;
reg [MAX_SUM_WDTH_LONG-1:0]                I618d33f26badabfa578908903a613bce;
reg     [1-1:0]          Ibe387e8fe6f35588e028ba29cda5b912;
reg [MAX_SUM_WDTH_LONG-1:0]                I822d7973afe090b2764335f1b72dfd0e;
reg     [1-1:0]          I98191a7e6c56aae1b56e3d623004ed75;
reg [MAX_SUM_WDTH_LONG-1:0]                I12c1035353e553b3b6a13bb174ce6020;
reg     [1-1:0]          Icd0f5c370462670cd18d30dfc0c81c02;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia6d61947d36fc128c689808c82db80f6;
reg     [1-1:0]          I15c59dc8eba10ff8eadfa6078678773b;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie9b042f686381739b9ff219041f1e0ce;
reg     [1-1:0]          I3870d672343c002ad9c83c816fd40567;
reg [MAX_SUM_WDTH_LONG-1:0]                I0c4268c01aed70ce4fc71531bf4bb862;
reg     [1-1:0]          Ic341b9d947f2d3ac57aa41f408214434;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia34e42f8de91fa4861b0c6cac5dcfc29;
reg     [1-1:0]          Ied40f6b7847158bd08cbd932254dd6ba;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib7c5850b4f7cc77be2048d114a2128d9;
reg     [1-1:0]          I6ab04d323306b7290cc89ed66dbd93bf;
reg [MAX_SUM_WDTH_LONG-1:0]                I32bb50faa2b246b2d3b462a79be597c5;
reg     [1-1:0]          Iac4a5fdede87b021e6a8150d3bf34b66;
reg [MAX_SUM_WDTH_LONG-1:0]                Idc6d40a49f05c5422758cee50f787eb1;
reg     [1-1:0]          Id92b1676e19c5818fa813d06dc9a01f3;
reg [MAX_SUM_WDTH_LONG-1:0]                Ide1d7dc22a4b271ef764df14ac22366a;
reg     [1-1:0]          I93da1192f27c33e21e03b9a2748774ea;
reg [MAX_SUM_WDTH_LONG-1:0]                I7ace6778ac86b3e05939a3fcc716136f;
reg     [1-1:0]          I69a0c79d41af6b6340430b8b337fb0ca;
reg [MAX_SUM_WDTH_LONG-1:0]                I044e01e8d2df46e03f00a0af2beb0bf5;
reg     [1-1:0]          Ibd47f48d306ec44d94865a0a81e4f9dc;
reg [MAX_SUM_WDTH_LONG-1:0]                I45a7ddcda2662e36b7617dfe64514346;
reg     [1-1:0]          Ia5707d1275138a5145b2a42190d95183;
reg [MAX_SUM_WDTH_LONG-1:0]                Idada779a1ac7b844867571d77054b657;
reg     [1-1:0]          I33bc2f42d997a2963b063326eb210d1c;
reg [MAX_SUM_WDTH_LONG-1:0]                Ieeba01b18a244ab8c0ac263c138fabcc;
reg     [1-1:0]          Ib22e39b701614cd9986061c32adfbc66;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie4c9797a955778694dd8615219cb51e7;
reg     [1-1:0]          I9b08176fde1cd08c9d7686a659213580;
reg [MAX_SUM_WDTH_LONG-1:0]                I28a5ed4c239e64c76bb6e566b50cfd23;
reg     [1-1:0]          I1b4e65357a818998d08b83d21584e18c;
reg [MAX_SUM_WDTH_LONG-1:0]                I79a705ee1e414fe4a5fb14e9b3ce9597;
reg     [1-1:0]          Ibb865ea5891db706b7b54e5c6fa383d0;
reg [MAX_SUM_WDTH_LONG-1:0]                I04f90a907f10a7fa1ae3591b48094d5c;
reg     [1-1:0]          I32d42cfd2d516af2e68fc2db4d5dce03;
reg [MAX_SUM_WDTH_LONG-1:0]                I31d25b1b49e65216e90b39aa27acd6be;
reg     [1-1:0]          I4d0e8d475a5d2a7da24daca60f23f3d6;
reg [MAX_SUM_WDTH_LONG-1:0]                I1f6540c5f037d861dee2c0091cba01ec;
reg     [1-1:0]          Ie3850345b207e59aaaa5c944dab40b90;
reg [MAX_SUM_WDTH_LONG-1:0]                I9632bb500b7faaaaeb649d74c21cbe8c;
reg     [1-1:0]          I4a9a1c932db30dcf04cb105a8d7384f9;
reg [MAX_SUM_WDTH_LONG-1:0]                Idd0217a35c3adc8abc7bb581a5df7a2d;
reg     [1-1:0]          I0ef689822226332f5feaf79fcf8f6674;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic05b46168884322644db4e331d37d759;
reg     [1-1:0]          Ib5744c2130bb5a9d0ccdd975fdf2ff9c;
reg [MAX_SUM_WDTH_LONG-1:0]                I53c88dc237bb2cd02d50fd7f0a168a48;
reg     [1-1:0]          I039a7ddcb25972501d80c45c938cf683;
reg [MAX_SUM_WDTH_LONG-1:0]                I7450d4ab3ef0227e93a02bfd620d047b;
reg     [1-1:0]          Ic5f36c15ebad061dfbd5301e02ce2ffe;
reg [MAX_SUM_WDTH_LONG-1:0]                I2b16e5b4e279bb29c3c675b72083e5fe;
reg     [1-1:0]          Idf0d9dac06522293f8d7e00a93b6bbb5;
reg [MAX_SUM_WDTH_LONG-1:0]                I70c92e8ada46476d15ef4b3c620d2601;
reg     [1-1:0]          Id557db735a70dbb14504bc3088e8798e;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib193b07804d6d5f111b06bda487bfa5f;
reg     [1-1:0]          I150d31ef31093fdfc5f145d84bb35156;
reg [MAX_SUM_WDTH_LONG-1:0]                I885433b0ab16c6d87abe45af13c9e529;
reg     [1-1:0]          I7e40e6f9d82d9b9fc546672e8e8621bb;
reg [MAX_SUM_WDTH_LONG-1:0]                I198c055930cb89d0390c336eda8fed4f;
reg     [1-1:0]          I14133cbbfa6521c5b81477fa1c229cbf;
reg [MAX_SUM_WDTH_LONG-1:0]                I688a2c72e69b217d2673e8da75146a83;
reg     [1-1:0]          I3728e31a7cf48639ce873d9135dc87fb;
reg [MAX_SUM_WDTH_LONG-1:0]                I3b6fde4ed14cd68af1468ae1d4cc1a22;
reg     [1-1:0]          Ic6be12e390bd3c25c66d9b9e7c0532b8;
reg [MAX_SUM_WDTH_LONG-1:0]                I5d3df1e7563630311f56143ee6d97a8e;
reg     [1-1:0]          Icc50e1923274729fe472ca578b68c0f5;
reg [MAX_SUM_WDTH_LONG-1:0]                I90a7ea789d3bf7f9126c786474a56da0;
reg     [1-1:0]          I4d98064f544a41b977ba945d2eecdf21;
reg [MAX_SUM_WDTH_LONG-1:0]                I5029424c9d9fe923eeb858b1e62cd758;
reg     [1-1:0]          I12f2a9f1e3e715d7e684ff39dd7942f0;
reg [MAX_SUM_WDTH_LONG-1:0]                I1e805c70d50c2765b4a03ad2982dc421;
reg     [1-1:0]          Iaa4e3c53a0d55e8f42f60ff40893427e;
reg [MAX_SUM_WDTH_LONG-1:0]                Iba58175a7fd5c5da650222193caff0b3;
reg     [1-1:0]          I26aae317b0b320df86ca4004f64aab88;
reg [MAX_SUM_WDTH_LONG-1:0]                I7401a0501ba69c5559fbf00c77e58dc5;
reg     [1-1:0]          I9344825cc2e5864f691043a1f94f86a4;
reg [MAX_SUM_WDTH_LONG-1:0]                Idd9f7ea657ea9cdcb45a7e4b573b9d50;
reg     [1-1:0]          I82988c3879c1de76fe2140c469f6a4c1;
reg [MAX_SUM_WDTH_LONG-1:0]                I53f275395dd6be17961a5edc3e8da7f2;
reg     [1-1:0]          I6bdd8334512c7c6a3226ebb4e928a270;
reg [MAX_SUM_WDTH_LONG-1:0]                Icab010d78cd66b02e089c74f04bf4e75;
reg     [1-1:0]          I0debec6ace7160558cce7f111dd1bea6;
reg [MAX_SUM_WDTH_LONG-1:0]                I376a48b7e0195a5aacc76a0ad8bd14b2;
reg     [1-1:0]          I8ee02e65ce9183683f0f3168bfd755c5;
reg [MAX_SUM_WDTH_LONG-1:0]                I241622b0367dde514f96ece55c8c3964;
reg     [1-1:0]          I80e6d2c9c5f7b6bc6bffa063c4959115;
reg [MAX_SUM_WDTH_LONG-1:0]                If94a1abfb972f63629d07e64dc23863c;
reg     [1-1:0]          I0f21fb041239a7a8895c9506f2754595;
reg [MAX_SUM_WDTH_LONG-1:0]                I07b9b1f4fa01b16cc69356057d3b6154;
reg     [1-1:0]          I8ce37a8e81b54043276835c11e394df5;
reg [MAX_SUM_WDTH_LONG-1:0]                I2288a6ad3b748b716249f4adc42d52c4;
reg     [1-1:0]          Idf7d1f78735ce1e9695d99a532a7726e;
reg [MAX_SUM_WDTH_LONG-1:0]                I022df337bcc05ac5648b8ae2e42f3a76;
reg     [1-1:0]          I96a552ed2d18c0ba3fc6cb6d6b6a0f44;
reg [MAX_SUM_WDTH_LONG-1:0]                I60d9a7f95fb8623753002ecaf9a4efcc;
reg     [1-1:0]          I3c76936e8e3467378210a13645a401d4;
reg [MAX_SUM_WDTH_LONG-1:0]                I23a74ea5e7174d95e6d16a5e85ac236b;
reg     [1-1:0]          Ic9a1d599fcfd5dd51265e5d0989719b6;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie697d28d757df82b3901564bda43251c;
reg     [1-1:0]          I60156470e631268c392040d3c5582eca;
reg [MAX_SUM_WDTH_LONG-1:0]                I8572aedc94f7243ce5eacb332c81eae2;
reg     [1-1:0]          I821126d1516ad7e8191a7b2a3b5e4b47;
reg [MAX_SUM_WDTH_LONG-1:0]                I6734123aaf6320da75638b212812732f;
reg     [1-1:0]          Ibe72e9f6d2c3cbbcf98f6b5aa6a4f93b;
reg [MAX_SUM_WDTH_LONG-1:0]                I7f6dc6f0f403c58f9aaaa70c2383a666;
reg     [1-1:0]          I1e8b6306d2dfde4a36ee9b9c2caf1c85;
reg [MAX_SUM_WDTH_LONG-1:0]                I66391978843c39b6acbdb4847a01050a;
reg     [1-1:0]          I48ed92480f457fc3cc2ff0dd7d177a10;
reg [MAX_SUM_WDTH_LONG-1:0]                I4f756e4125c8af5c412944b273e01cb0;
reg     [1-1:0]          Iaed28d88a651f0151501ec4ea6ee3346;
reg [MAX_SUM_WDTH_LONG-1:0]                Id2c9f7ac95de07148c54803f69347f56;
reg     [1-1:0]          I9d94d9b5414662de841443d7866e66b1;
reg [MAX_SUM_WDTH_LONG-1:0]                I5061e13a179d27e1ba5f89ce8ee0fd4a;
reg     [1-1:0]          I870b8a3b11be215a8704ba05568f05e2;
reg [MAX_SUM_WDTH_LONG-1:0]                I0f7c32fc1548fb49b8041f55c157498a;
reg     [1-1:0]          Ia8bbf21e040b326058a9acb7d198a835;
reg [MAX_SUM_WDTH_LONG-1:0]                I89ffab735ee30423c82e079ed98216c5;
reg     [1-1:0]          Ie852f207c8f537621b080ffa0a89bfdc;
reg [MAX_SUM_WDTH_LONG-1:0]                I9494921d8487ee0b314f75cf0380fd2f;
reg     [1-1:0]          If53029b05bea46d656a6ef72fb6d6642;
reg [MAX_SUM_WDTH_LONG-1:0]                If2b3e7d1541cbd8ffc2b4cfc3ad13a57;
reg     [1-1:0]          I8e8a740d09e000444ba1f4931b5cccf4;
reg [MAX_SUM_WDTH_LONG-1:0]                Idf3d79da44f2d686f5bd43c3c1427430;
reg     [1-1:0]          I46605d823e06af5485e50b256b5c3f22;
reg [MAX_SUM_WDTH_LONG-1:0]                If8125ad3c9e7f0a2b84106064d320996;
reg     [1-1:0]          I38344d68127f5c035193bb9030ce4d4d;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic9018b88fa91fb638bbab0613795ae13;
reg     [1-1:0]          Iba9f33c08db89a7f120cc1e3eaf05dec;
reg [MAX_SUM_WDTH_LONG-1:0]                Iad4ea0196eb32f9a152c9e6fe5059e46;
reg     [1-1:0]          Ibde51eb91b3ca50a8a0513c94bd7be15;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia8ff29ed728e7f2ae4213f00328b495d;
reg     [1-1:0]          Ifb94196d1653a0166567e170f06ec0db;
reg [MAX_SUM_WDTH_LONG-1:0]                I70717726200ec02929f679ef05496455;
reg     [1-1:0]          I9cf7557e2cac4532a77fcb212712db0f;
reg [MAX_SUM_WDTH_LONG-1:0]                Iaf1e4c7dae6ad89567836877c08f57d2;
reg     [1-1:0]          I3159d7faeee1a904c409bde1967d2c21;
reg [MAX_SUM_WDTH_LONG-1:0]                Icd09aa81e9b43528af73e23b2f0f80cb;
reg     [1-1:0]          I35dfb5ece5e04504d6e74739ae99c9cc;
reg [MAX_SUM_WDTH_LONG-1:0]                I6ebb2b94f0f80425f8401ae823d92a1d;
reg     [1-1:0]          Iabff939ae4acf7d7b038e028c29b6166;
reg [MAX_SUM_WDTH_LONG-1:0]                I4a2c3204a6a9936d4a215b46c0ffd045;
reg     [1-1:0]          Ia14159444578c6dc88f2d5ea0317774b;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib02c0694762c4815448b2c8d3df767c2;
reg     [1-1:0]          Ie2306a5c441d621388b73195027fc118;
reg [MAX_SUM_WDTH_LONG-1:0]                I98cee6efbbe565d3a4de16703189782f;
reg     [1-1:0]          I700a0fbf81e57d4970ce07090ec4f2e2;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibf981c01a9d44cbea3c6d8ead92bc2ab;
reg     [1-1:0]          I6007914b3fb3011c3ab2f9a9d7794ab2;
reg [MAX_SUM_WDTH_LONG-1:0]                I864c33e8ea204d20a9baef4584f22d4e;
reg     [1-1:0]          I2096f40fe62e9d6f1ff96f258ffdbe33;
reg [MAX_SUM_WDTH_LONG-1:0]                I6ad3228e0e2e1f19648d73e83ba5a229;
reg     [1-1:0]          I93d8b7a24702bacbfc528242991516a9;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie099210a99a4899c53baf39559592690;
reg     [1-1:0]          If0863fae91b2ec980ebdb26cfc90ae2e;
reg [MAX_SUM_WDTH_LONG-1:0]                Ieeec71d9df4613555fade2ced7b3baf1;
reg     [1-1:0]          I9ec29a319384efd562c2337e1857cb4e;
reg [MAX_SUM_WDTH_LONG-1:0]                I4931884e3544af182bcda9061091a42d;
reg     [1-1:0]          Ia56ecc024eae608d7de1509d75139dc2;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib3fb10da528d450251764a9b9ede0dba;
reg     [1-1:0]          Iebcd65ea41cd38bfe3c8577277809acd;
reg [MAX_SUM_WDTH_LONG-1:0]                Icdc9e676957b2223d60c413331fa982f;
reg     [1-1:0]          I75be12b14694ebcb5aff6e5d3e576315;
reg [MAX_SUM_WDTH_LONG-1:0]                I381f6051282c062ccf53866830344cd4;
reg     [1-1:0]          I8e06fe414cd04103baf3882771a63e2c;
reg [MAX_SUM_WDTH_LONG-1:0]                Icfc21935c007fbbceb2a67ebe1a68a0b;
reg     [1-1:0]          I0fe8574049166c363c7cc816b1435009;
reg [MAX_SUM_WDTH_LONG-1:0]                I120d597a80158374726e064fb0f099fb;
reg     [1-1:0]          Id5f435c07240d5fe4a0e48c8f25ad0b7;
reg [MAX_SUM_WDTH_LONG-1:0]                I2520aa556aadf851f58f0b1820498730;
reg     [1-1:0]          I1ae21e0db88f955c4f08f6d52f58974d;
reg [MAX_SUM_WDTH_LONG-1:0]                I6203f49a08107f7185ebadeecf2c16b0;
reg     [1-1:0]          I92efddd59e1ea92902a295c0b8385c68;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia706fb593b63cebbee0321c154cb859b;
reg     [1-1:0]          I56948ad2b2cc245bb1003fd71ae5f899;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia4b5f2b07556629673fc6576bc49a5dc;
reg     [1-1:0]          I5fb5081b7a2da89115c0080b0967974d;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic532c6b85b156f821e0742f47239a65c;

/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [22-1:0] [MAX_SUM_WDTH_LONG-1:0]      I583b1bfc712ec29d08acc68c27675882;
reg  [22-1:0] [MAX_SUM_WDTH_LONG-1:0]      I95878a848ec38c4f334bc1915576e6d6;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [22-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ifba287889bea3585954fef5efdf5bb24;
reg  [22-1:0] [MAX_SUM_WDTH_LONG-1:0]      I3eb1902edf9266038f39c281d134c26c;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [22-1:0] [MAX_SUM_WDTH_LONG-1:0]      I8e5ae9e6fa38cea8e5d320fe582c0729;
reg  [22-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ie791b43e8d5c9d1669743ea4d6e3139c;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [22-1:0] [MAX_SUM_WDTH_LONG-1:0]      I67315420a608e257df8cfb520ef9f0a1;
reg  [22-1:0] [MAX_SUM_WDTH_LONG-1:0]      I5b892f00b2642ca102f7755ab512d067;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [23-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ic80a23c7b47f2236087fd7818d8d7c7f;
reg  [23-1:0] [MAX_SUM_WDTH_LONG-1:0]      I8f906015dba99b4a73dcf767cbd948ee;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [23-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ie53d62e3ef9caf35092d7a63be1f565f;
reg  [23-1:0] [MAX_SUM_WDTH_LONG-1:0]      I9ab4bbe4191d0f284defcdce6b885054;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [23-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ia73bc9712b861f909d0e3683ec91ea1c;
reg  [23-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ic8a3b3e2aacd0eb24cbc429e9bb734ee;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [23-1:0] [MAX_SUM_WDTH_LONG-1:0]      I97d2ee9c3120e78ebcda2f0dbb888b49;
reg  [23-1:0] [MAX_SUM_WDTH_LONG-1:0]      I6ff6fafd1a3364131b269724ad273ba5;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [10-1:0] [MAX_SUM_WDTH_LONG-1:0]      I07b2a00225c337eed1e5a350f3361240;
reg  [10-1:0] [MAX_SUM_WDTH_LONG-1:0]      I154fcd3171f1231e825ee603d53ecfe8;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [10-1:0] [MAX_SUM_WDTH_LONG-1:0]      I64c650bb94f04521a5a33efa937d9cfc;
reg  [10-1:0] [MAX_SUM_WDTH_LONG-1:0]      I489e70342dbba4a551097e3064dc9835;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [10-1:0] [MAX_SUM_WDTH_LONG-1:0]      I34152d4ef2dadfcc943a004e81d175f1;
reg  [10-1:0] [MAX_SUM_WDTH_LONG-1:0]      I0b0a1f577a212bd9024c8b9a44c92e00;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [10-1:0] [MAX_SUM_WDTH_LONG-1:0]      I745f84653760acc2d83607dcbe1eec73;
reg  [10-1:0] [MAX_SUM_WDTH_LONG-1:0]      I40d311bab75b73e3788c50115a205270;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [5-1:0] [MAX_SUM_WDTH_LONG-1:0]      I9efcf5ce8571b24b590d2d4c8161d49d;
reg  [5-1:0] [MAX_SUM_WDTH_LONG-1:0]      I5fa015a360308bffc46921d119b60c1b;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [5-1:0] [MAX_SUM_WDTH_LONG-1:0]      I60a6ef79e3a8244ad32b9833a6ec196b;
reg  [5-1:0] [MAX_SUM_WDTH_LONG-1:0]      I9e42bc767599ce3cc4e2d886e5ef2e62;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [5-1:0] [MAX_SUM_WDTH_LONG-1:0]      I849584bb1c2436f764968afcbb14a61b;
reg  [5-1:0] [MAX_SUM_WDTH_LONG-1:0]      Iea43b150eabf3c7781275821eee3e0c1;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [5-1:0] [MAX_SUM_WDTH_LONG-1:0]      I3ed70f2b460f9278ddeebaf6919b77e8;
reg  [5-1:0] [MAX_SUM_WDTH_LONG-1:0]      I8012eea3d53fa4e000eb28b121e02ada;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [5-1:0] [MAX_SUM_WDTH_LONG-1:0]      I37b4978577c93e476e4a0bc15b9008c9;
reg  [5-1:0] [MAX_SUM_WDTH_LONG-1:0]      I49804415d20c0c087f802b25dd609887;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [5-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ieeaf46eef680115f0d2d108b84b5d3da;
reg  [5-1:0] [MAX_SUM_WDTH_LONG-1:0]      Id270f05bf5c3fc0bb211d1665d149044;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [5-1:0] [MAX_SUM_WDTH_LONG-1:0]      I8b4ff33c17efa28c7eff64664384cffe;
reg  [5-1:0] [MAX_SUM_WDTH_LONG-1:0]      If091fe044c792be711325c103b84cf1d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [5-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ia453e66ce9c1335efac95deebe00c249;
reg  [5-1:0] [MAX_SUM_WDTH_LONG-1:0]      I1550db301291ab131a5536147fb938f6;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [14-1:0] [MAX_SUM_WDTH_LONG-1:0]      I9c5decf5be3d3e4222559a9c244afc6b;
reg  [14-1:0] [MAX_SUM_WDTH_LONG-1:0]      I74d1345ee56f5688f875823a5d7c1f4f;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [14-1:0] [MAX_SUM_WDTH_LONG-1:0]      I56c4270727a90e00c295c578183a4dce;
reg  [14-1:0] [MAX_SUM_WDTH_LONG-1:0]      I187371a49a27a988920854b2bb61bea5;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [14-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ib3e1c6976da60eb724a8d00f19368423;
reg  [14-1:0] [MAX_SUM_WDTH_LONG-1:0]      I48c4c6e7414394e3aeff9d17ec25d020;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [14-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ib53ea6bc0e3ac45d5a8eecd5dce775d8;
reg  [14-1:0] [MAX_SUM_WDTH_LONG-1:0]      I3cba0f4c2ca8c7c200df8e1071ab429d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [7-1:0] [MAX_SUM_WDTH_LONG-1:0]      I922408509703b8175883356d89806972;
reg  [7-1:0] [MAX_SUM_WDTH_LONG-1:0]      I35688678e1a83ec39d737d9cdfd44ba3;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [7-1:0] [MAX_SUM_WDTH_LONG-1:0]      I6cabc68155bc4aef952a07f101ea2802;
reg  [7-1:0] [MAX_SUM_WDTH_LONG-1:0]      I94b86d31e8226723950096e91855b6d3;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [7-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ia894c8a3585def468e93aa51039d405c;
reg  [7-1:0] [MAX_SUM_WDTH_LONG-1:0]      I0ea7c4721ee0c13ad15a9b0fa7b15ad3;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [7-1:0] [MAX_SUM_WDTH_LONG-1:0]      Iaf1c895fc85487f017d3c084e125551c;
reg  [7-1:0] [MAX_SUM_WDTH_LONG-1:0]      I29dd5fb1c2673cd4daa9cafaf24d8e7c;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [13-1:0] [MAX_SUM_WDTH_LONG-1:0]      I63d67a9bf5a46800216b38df1eb185eb;
reg  [13-1:0] [MAX_SUM_WDTH_LONG-1:0]      Iead4c81d836e3befae55049797c30d6b;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [13-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ic087eef7b3d2a51f34f317a6b9e49144;
reg  [13-1:0] [MAX_SUM_WDTH_LONG-1:0]      I23e22f44791c167acaba27c91ef3b497;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [13-1:0] [MAX_SUM_WDTH_LONG-1:0]      I6d360540762be9eab571c0bfe0500f67;
reg  [13-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ic91f087829e0b9e0c964229a2dc567bc;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [13-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ieb702849c7e744c5d04be8f86a00a4fa;
reg  [13-1:0] [MAX_SUM_WDTH_LONG-1:0]      I0fd9bcdcf8faaaabf94649881419c66f;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [6-1:0] [MAX_SUM_WDTH_LONG-1:0]      I8519162455bacafeb7f45c170c0b5e7e;
reg  [6-1:0] [MAX_SUM_WDTH_LONG-1:0]      I7cbcdd5018de9ceb49554b140e5665e8;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [6-1:0] [MAX_SUM_WDTH_LONG-1:0]      I0d7c184fb7627c9c50a0026ac5052448;
reg  [6-1:0] [MAX_SUM_WDTH_LONG-1:0]      I5a79c19fd2093d974b574e85245b5617;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [6-1:0] [MAX_SUM_WDTH_LONG-1:0]      If5cd4834f1cb99b40cd4084fea388070;
reg  [6-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ica937143b618734fa099683949153130;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [6-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ia3aa64fb9d2eb1168da1f7e178c05c4e;
reg  [6-1:0] [MAX_SUM_WDTH_LONG-1:0]      I2d4d5d2694718b39e80b89b422d690cc;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [8-1:0] [MAX_SUM_WDTH_LONG-1:0]      I58c319fa3e05e8f7ca440775482ba8fe;
reg  [8-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ic2faea3d4bb97dda16ecc29c27939ca6;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [8-1:0] [MAX_SUM_WDTH_LONG-1:0]      I23f3a4487998f2384d9323f9103f7aca;
reg  [8-1:0] [MAX_SUM_WDTH_LONG-1:0]      I503e83a1146c42d5c1ef011ecb280807;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [8-1:0] [MAX_SUM_WDTH_LONG-1:0]      I081087845b5c62dc79fd5b9882339572;
reg  [8-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ib9886c1fcd27ceb24afb2d0d7da85c26;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [8-1:0] [MAX_SUM_WDTH_LONG-1:0]      I8aa441e2ed6f41bca12ddbeaac9f5c3d;
reg  [8-1:0] [MAX_SUM_WDTH_LONG-1:0]      Icd90612c09423a2817a72f750e585309;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [9-1:0] [MAX_SUM_WDTH_LONG-1:0]      I4bc30140a67bbc7b19449fcf946a17aa;
reg  [9-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ib7b7884d2653893806af34579f7c0760;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [9-1:0] [MAX_SUM_WDTH_LONG-1:0]      I943f523a14e49f42d9c6ceb3ad1dd841;
reg  [9-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ic3f0ad21d8a446c31afec49309a18133;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [9-1:0] [MAX_SUM_WDTH_LONG-1:0]      I10ab80965b99680e93ea304f6e261094;
reg  [9-1:0] [MAX_SUM_WDTH_LONG-1:0]      I2dd65bec7d2bc4778b7fc48a413d2ba7;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [9-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ibfef15cf57c5850241c05384f18da5ea;
reg  [9-1:0] [MAX_SUM_WDTH_LONG-1:0]      I36b5867a3da6f2ed529e791166640d3f;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [16-1:0] [MAX_SUM_WDTH_LONG-1:0]      I0aa8bcd235f4c4f32c3075d5f39bc20f;
reg  [16-1:0] [MAX_SUM_WDTH_LONG-1:0]      Iedc20522d3322bbe3f55e2aa611d76df;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [16-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ic5e951c3193081b1880ccf868e740e92;
reg  [16-1:0] [MAX_SUM_WDTH_LONG-1:0]      I6821e897aea31f7c237ca1a553bf0cd1;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [16-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ie8edae9436451bc0a4dbdbf531401682;
reg  [16-1:0] [MAX_SUM_WDTH_LONG-1:0]      I290499340d94dd8e234f53f9962a182b;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [16-1:0] [MAX_SUM_WDTH_LONG-1:0]      I84a56b9dce9dfafc97fbdc2ad3b2ae68;
reg  [16-1:0] [MAX_SUM_WDTH_LONG-1:0]      I5ce387684404cf922955e4af33ed2367;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [9-1:0] [MAX_SUM_WDTH_LONG-1:0]      I8afac763670df6f56525d3192e04e784;
reg  [9-1:0] [MAX_SUM_WDTH_LONG-1:0]      I1ae87f851f8bd64e6e1428a143e82151;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [9-1:0] [MAX_SUM_WDTH_LONG-1:0]      I8cd574c061a4f1bb0da529d2a892324b;
reg  [9-1:0] [MAX_SUM_WDTH_LONG-1:0]      I646767a2d4b3029ed7acb73a15af1682;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [9-1:0] [MAX_SUM_WDTH_LONG-1:0]      I919a7f8471a46de33447530b4f3b591d;
reg  [9-1:0] [MAX_SUM_WDTH_LONG-1:0]      I48001f5c6554999a2178308ae271b70e;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [9-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ib1f53b5c820345ccdba27ab5be3fa49f;
reg  [9-1:0] [MAX_SUM_WDTH_LONG-1:0]      I7fe6d853fc1c11142b64ff8f40783246;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [12-1:0] [MAX_SUM_WDTH_LONG-1:0]      I384c493c3195d97eea0a9faaec860f78;
reg  [12-1:0] [MAX_SUM_WDTH_LONG-1:0]      Iadc98deb917f599574e99a90e3230e88;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [12-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ida1ee79b7a153e40e91549c2180d8425;
reg  [12-1:0] [MAX_SUM_WDTH_LONG-1:0]      I3d79461a85cd6a58bf9f96f6e0d704ac;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [12-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ib6bfc051a54fef77204b41e38cdfc6a8;
reg  [12-1:0] [MAX_SUM_WDTH_LONG-1:0]      I2fcbccd884710be9c6a34f78d2ae6a18;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [12-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ie6d740bc0451311c5f93f4954812613d;
reg  [12-1:0] [MAX_SUM_WDTH_LONG-1:0]      I3d3df5d4d89adf508497bac8d75ef0c6;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ia6ac09257dfd071a132e96619a662f57;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Iadecdac113e45cd08e095317d07766e5;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Id2e5704c73c707a217875dbf2743e6f3;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I2e4a339cb29f80caa8cbd630a0372ae8;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      If152a76f9c612e979151b8f51262efc1;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I423e8e9a9f19cf712372622e5c80c732;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ifdb6febe29caf3ce300d9cea4954927a;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I5434db7480d96327d98156af57961745;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Icfb2b3a2e096f55ba29dd2f9b5761852;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I20ebcbecf2c13a53be05ff26552b4e72;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I06c6597547e69bb46e1bede7b7b7f24a;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I7ba72e4bac9bd64d046733ce50f43769;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I325f629c52919e62b3c0075481267744;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I6614526a756edaabd6a25e858b472d14;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I56dc657b33a933d2e5d3ac517a9d1fef;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I47b2e8ee0c69e5301365a25d512b1ece;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ie17d5d171cb71e3748dd0b6c800263ca;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ibb72eb38996b41ce253875df0f620eb7;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I9cabb772f5988b877afae0c3b65f340a;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I66944cd8c5bc22cd92a5cfcd68cee426;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ie29294b754845c1c5602dade95c9e762;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I8f2ff78b78e43fe7f6780f19d92ff7b8;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ibfc5db8e8f393324f06568278da33b4e;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ieea0e49da41cdf0d062217a6e6591728;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I44aace203d154a4d0fc8f10f2cdc5626;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I699c35d4b3c36c35ecaadb87c8b35d9a;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I75526eea62d190615e13ac2731e07074;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ie6c95c6ddde379ca7437e78c42a8245e;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I67bc090d5c81788569b837217febf22d;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I85e05de515eb28d7172a95ba55da82a2;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I28d725840d5db12ad4940ef965775cc4;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I7ed14b994ecbeae0536a721e16c88489;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ia9e617fb96d7ae3706736fafa5dce67c;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Iad29b892bf50a3e83e4eb9b7c271292a;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ie033e6fdf59cdfd67ff238b68924dfb5;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I35d2bc3f0efd23ded421f195b62a6a33;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I6190c7e2fd99fcb3394fc330e0b08678;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I4aaa94237ac5b28ce1d0db0d4e15ff81;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I91f50b160f3a0bc73c84123d977fa4ab;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I137145b608dfe5138d4bdbea237743bd;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ic05ea9ae53b9396b54c4484a56c7ec79;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I68a784efb51b172af79e3dec88d529e1;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Icf4d6deb47e202e607a07639d064ca55;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ic3036adab4495c6a59055dd34a28b2e5;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I85ee05cc8e67b77acbd3ddc7fdfd6bca;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I84a699063d2a7944f4a1b72b67ab5b4f;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I803822a38e626e789a50bade0961edab;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I63acf3ed504ad084a12a219790842b4a;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      If93330fbf9bc863d2837ffc2a0466e70;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I23a2a7fb24650eec8812d8671d92bf2b;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I8ac880ea1c849c493c66a82534400d8c;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I6f9156b7b5e13529ec0c34da34cb2b04;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I7cf96d4e28b02fd623d8c76161410eb6;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I09a4c92baceef72d764c6880fb62c1f7;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I637636f1d78f96c75bf5c3841419e9fe;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I13a44a5dfbb198be64c99845122a6e97;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Icc7d8812ba512a84d2905f1182e69d0a;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I2b57472e34677b9aafb852a3e421270d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Iba60ce25380dc39b44ba505a04453614;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ic96e056f2208c211122e5008d5fd8ced;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I9a6a2b184e5122aaa964c2bc818c255d;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ie6b1ee6dfca427a82e4d1016585682d9;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I4dea7825b6a0eab3aebeb7c4889cdae9;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ieb0276790e2d912809acc7f3a409ac37;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I4809ebf07d855a2e48f92df77ac08b89;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I9883bdcc250c2eb1f8e691d0f18b3cbc;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ie0a958d83a20d204b3e7a9b4235c4b19;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I28f58fec52ea2df3fa3d8e4a2722468b;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I8280db7b6ab8c525afd18dc79c0715fb;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ibf1bb88a30c8519cf22f684a9bc552e9;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ifd4e06675d2b57e0064369490c20b8ba;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I9d2131bc965972708385d8d79c5b1687;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I887915cd3be831277d41e47417ae42e7;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I65dc268c49445ceeef922f9c273df755;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ic3af54bfe225c905cd146c6ccd3e34e6;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I7c0af5fba885dca550df150029e9ee36;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ida4ab0033193d0b40f4ab5d8b74d7625;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      If26299fbf3d11a469aa2bc573760fed0;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ic0c2d77062c77982f91941bd99eea68a;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I2ba80daf0c2b625370644ab47cef63e9;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I783f9d09de5fce4d69c179fb398a58ae;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I0911e01c831a9e46568122fa6dab2357;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I0af2bc8f858473a4b6f9467d5635f2ed;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ic8f0aa27dadc689b1bfb5b284fc13562;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Id882b47b85085b9603449499ecfcdb49;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I5ad4c6aba210a8b2d343ab17b49c38a3;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I5b2752f489336c41887046ed4673a717;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I34947a54412d287f3ff730332211dc5a;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I75b2328b94afd38404e28c46d7358b22;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ia6ac380b9be591fb53c0f36f4d417a7e;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I7a642ae71b9f5454a31702d6c3197c79;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ia5d5342af30d46f66f0e4f41e5170b87;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I0f8357de84a9c9e19d35ddd0715b7be4;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ica011579f46e949eda7f8eed2e4d3ada;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I76599476765ec5b54c1ed75efddc909d;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I88b214aeebaffa768ccf7c70423fb0c3;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I9e277097d3f55ad75b5b0e819d6d3651;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      If46340645f788fdde3bb8f4d176aae52;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ibade670ce04ec07f3b5174fcfc67fabb;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ib59f285283d8c3013c20aad73ed9d148;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I19a9636de4b8153208ebef0cfbf811ea;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I3229ea9a0c348b17fcaedf6565d6d7cc;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ieb302f84fbd92b0fa4a5747cb1764926;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I3ba17818aa7ea9bbfcebb2a5f405fec1;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      If88f7bba0fc9ca004e41cf047f6e6410;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I2ad1769ceb4cf0013f7b032c6e583745;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I5989aa844d0d73de1a11b8902002efee;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ib35d4bfa08a9364f7f6c8be7feaf15ba;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ia683e321a3334e9668b39f5fea591cd4;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I216edc2024d31f612d05617f6696c6c5;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ic16cfcc11cd03b06afab4b96ab13a350;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I2be51c29373fe2ddfe456265a54bcc08;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Icb19ea7dbeb8d826bf85e1e8518e7558;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ib3561cb8090e7787ad8c324db3a5456a;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ie1c0888b2c811ca399501f4669dd8267;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I5d701e34c6fea83dccbac286a36fcbbc;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I65008ba6af7af0ee93fd085692ff4705;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ie479179aee4de4208dda8af63ed9fb66;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I0818a864ca9a381fd4b8492410037437;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I0acbd9a7ed1409c7958d6c630a7f96d7;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I11e799346dda7e851c5d48f116216d5a;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I390dbe9907497b62162445c90f2f27fc;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I1bea6ddcb374caef97e35af1eb33d878;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I01d386885d97d770ff2ab01da72631a0;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Iae87b81938ba6be7fcfb902e35b55ff2;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Iedbfdad739e796202d764f909e6ac6b2;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I2cf76e56c5212c0921ac6725ca41be3c;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I41ded014d071bd714d053a8aed21cf5a;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I21cf97f59f8387bdd451934e800a501d;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I1f14df209c8c73fe390873ae05063afe;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I9c91a8ca3a41b5df249ad6e0cd9b6601;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I510a362375a9b9c75436ad01388de6db;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I02e4ad55fc6e12cd60370ae782bbd36b;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ic2f0b44a83961b8b49f4637ec6750f27;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I5192b23d7d4742e17ffcf58679d96734;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Id5cbccb1a2ccacf28b64ece8eec0099e;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I0aaea02d5fbc4cfe6478060df6a92441;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I9686b2d0e5248bfb6d3ef9b7c687ed05;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I64476c4b13b6612ab90845870c8fcec6;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ibe5129eb30f626925a3ab5ed5e239bb3;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I46cb13c147e8087f9f93618f946d0f75;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I2a656dad40cec86a53e732e78f00c269;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ida1dc39acb508dea4487357625f65a62;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      If06132c6a0060efdbd695b31c338faf6;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ief0a83a4d2ab6337a9a842850ed9c8d2;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I02fd20ab9e4fa12009b63fbe41d647fb;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Iabc0481ca8b87650597db2ab82d9526a;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ibb97d541a2ed2b0cbad273a09fef5594;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I273daf63e8da53e5e9b99de802715b44;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I0905c7e3678f66095194058bb72d22fe;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I9bec797aec01899ccab507296d7f4d53;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I81433ae67b7cb4dee0b2091f3819ea88;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Id769ce05d2596a106b4e750d272b6d86;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ia6249382442d1dd3062acc63f891465b;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ifcd0ef96ba3a7a7ef8ab4f64c5671f80;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ie4bd4c14051455f00efdb023c3b58173;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I2789f24264b92b82f7e9f34a5ccaa489;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ie64e67a2316af18c5835c3a32ae9290f;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ic9f02e5a9bad9928c784d38980f709ff;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Icaf94b3fea3e29ff77d4793b389c9d14;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I5729f3c3121489f404f8964abb3e842a;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I334991f6bfe06389e35b7a580982de1f;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      If076d265cc6b8f7baf4059ea5fa7525d;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I6390495458553670944cdbf57bd6ce7b;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I7acc5316ae2768ce90598a82ad196eca;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ibafc73f0a3486943914e197a7af4505c;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Idc81e8df0b1b36ee2885c180c992a8db;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I2ec83b82756dda6035ddff10dd41fed5;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I2f587d7d70873b05956908ded54c36f9;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I5f6abb1000e5416dd4d43fcd052321fb;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I7f013f76d9fcc1b14984188e7af2ec0d;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Icc865d7264dd89944317be21610dcf9d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ica4903599938b7e1996702a51a7e9ec8;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I6a301412ef9235f3a609baf10a4200dd;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I53484a61ff8b4273d872779c33b292d5;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I9840f42586460341bb39256726d39ca1;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Iae00c13f4457b91d9a252b5b2aa67780;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I0837554bfb175a9ac8a4cb17e091fa9e;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I208b29bdae3040b547e8e40ffdc96d34;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Iacd698956b9ea6f1649063ee612c7e76;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ic6378ae3bd73ac1ddfb25e7d7882c671;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I68928b2759202e358f75b08e162e6a68;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I81f95de60a5dd186e51f9f4bf0b624da;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I609f881624ec9034823c9f54f4fb9b6d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ic05bdf0bf00ca3ba90c6ee7728b2d49b;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I075a0a1afc1463e92edb5f7658395424;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ic74ef5ce41d9db0920015b60cd80dada;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Idf1030f0e2aa5e2605bcea5fbe0428f8;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      If54ee451267f16296945fca60801b6da;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I1b82e98260c3bdeb5183a3af470e2d4a;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I22af03550c9ffd5ee75db6b34f444612;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I75338af3ebc7b7061a499e98a5be1674;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I76d5529e20b89a706595f65abe004da2;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I9f863d33f3c727e13eb52e7563ef9d1e;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Iebca060c7873173db59d0e1a244a5f62;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I56b8e0a7e6d2229baa9908843c0208ce;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I39ebf0c6f66596aeb1c56eaf50bc6b55;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I3d04bcd17aa2b98b69dcd671b9666c50;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I685db637ba885fcd9a37a9457b56c827;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Id254880ed38db79c53facbdc0c4a6d1a;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      If659617a922c1800e53f789111d7f946;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I988a7c2c284c38fcd6682236dc2d6151;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I3cde77dbb4b236619f7d00d6212d8f46;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ida4c48caeba43eccdddd1748824ec551;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ic1f7f01098e573cdab8482bd3f0dfe0c;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      If9936b476bb351a9ecbb97e2088cdd6f;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ic229657d83879de9bd470c1739254faa;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I6cbccfdeeb675a8a99d4c394bc8e71cd;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I3e69a3b20cf7ac74e77887b37fc3a5d7;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I79a4a9dfcecca4073c101bdd9b738c7c;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ief74f9042bd0058f17af181156b58456;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ice57a50f53d13e7eaf25af23547b5fb0;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ide1209ba9c80b0f69b0f17a1320b7a33;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I8ff8106a70daac7c8932e88aeb6d198b;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ib8c08ba5cf3c7bd8233532cc8ecb4825;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I8f9d1ec03357f7f045196050511341a2;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I812e31439ca7c94df3d6bf578b60beaf;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ic423bfa7639075130324da59f2cca2fc;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ie93978ee93511b6ed29aad9aed8ee903;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I4eed402353a7fa22fcb11f2adbf6be03;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      If0c12a1750d279b90738aacac5b35e04;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ieb579bed6711928456b296873c5da9cd;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I0501ec6e9230839738818ae2b19a5b65;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ifdf316d14ef99080247091609b2c2a8f;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I9e9c3529814bb741e0e425dba9ba0abf;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I2a1afeffe5592e35349bfd4384de834e;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I3898f311fc81d9bbcda50e18e7f978e1;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I93f88eac6c04d26228b5d7a3b1d00a42;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I4bf59374718f169f17fea6adb9d9c7e1;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I8c32ed7572af2a6a41a415ff6c580f3d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ide127cda229e55eca7ef703c0d794e6e;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I9cc4cd2860ebe1e5d43eb6024ea32dcf;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I482955b75319360d2646b1f712acdbde;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I35b73e275ce37c06d10c227595c7c3f6;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I158984c3dfe52e5107e4aa64548c1ab5;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Iac4ee00e62d47494b2bfe3aff55506ea;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ibdfb487053f2567b45db76d12e9eb75a;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I6023ec90efcd1ac53ea71eeee1c996e2;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I1fc2b706279a62a29d90f261f211c3a9;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I6f2b0c5e254aeb7e967f86e914876171;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I988227c12ad87b2ced8fd8fd89eb138d;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ie9353d9dd97f3536dfa6bcc2c662bf40;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Id537c7ec3b2e195d892f7fb1a63dcf46;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I09fd28ae4656b1282feb899a40b9b233;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I92a93c16158990f624973e9cc487fc00;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Iabbb1734d7e19cd9c7329b30cb26cd3b;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Iab0879a7d17f0fbf2c2ed147e41d3f32;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Iacc03e49c3cd6749e4c49e13c8c8593e;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I762ebc964e606e803121e347086668e4;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I7913101e04088970adf3f1e7429cd06a;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I032010a0a18eaf23274cdff5c99442bc;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ibddcea3450984eb0b3cc3ca6961fa646;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I24956c032de466de716b6ab57dd8a265;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I0a863fcba425a8683ebbb35195ea70a4;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      If816e24bfd42448c3c0fb03b6e9e9404;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I8138f45ab1b8a10869a2a6078b6c214c;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I0903046199323180f148f13aedaa0ab3;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ie4c27f8574c8bad0b923796d2544f858;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I25ec8dfa866fe300e67a01944f893bf6;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ibea29d15c71d594e4e9cbe6a58ebc550;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I77ac8c7c5ea03d948931590d57c8d649;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I0b249349485591abcc09c4587efca78d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ief5d16bc74276d3aec10a56fe8234b8a;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I6bbe05bfdabac8f312c7800eca53be62;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I6bec62410ca887855fafaa4be4c09d72;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ie28e38c9881297e7ffae5c3aed4dfdd3;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I290223476b30aa41df98af3016119109;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I1358b8ab0933bd596c33b622d2f9523f;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I07e3ae59ec05fa46d6ca3398a42e287c;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I46ce01ea907e88cafb7d96d22b5fffd6;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I7b019b5e5991ad8497a048367d83341f;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I64c0e39b2f3c34d724ecf0f511a413c9;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I80f8ed713e4b0281f94804a0b66fadcf;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I6ffbd03867a92aea248506af197c2e86;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I8cd2472defb068d6e3af7070c97c25ef;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ie0a0c3e63be2145dc838faf227a84044;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I3689f559a9636f9dd4558e99424d6c80;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I58265e8a07eede7063d5a80db2412214;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I77c454b260ff3c291b59ac8679966ab1;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I6734d5f87b795f4a05510778c22b555c;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Iddb9b8c346479631362bfc4aa039b746;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I314ced88cfc50d8b2edf129a6a3bf1a6;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I3db9cdf51e4437b6e979f8c1a0be96df;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I8cc6f1dc58a26262f18f334b751385ea;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I2a2352cab4f2edc64f156ef7b5e5595b;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I18d34c481f17aae6b16b6d0a5aa85357;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Iee3314c9bfca7066dcbb138d5f46d1f8;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ib54b35abe1088393d275f4f45f7ed966;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I4883185d078ac45e5eb2d6dbcd2c875b;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ie339493197828e5bd69bc49ca91aeb1d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ie6242ba25d061a37a41d7ca41370e919;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ic5084e34e9626f2e423283a87ea0d91d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I99d9fb1f21a8aba32da690b3bbb786df;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I3fee16f7ef907bcf1e2f5b2e7ec77866;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I1328d62797b528de9c98372d828d4af0;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Iee529a0d30e79cdc9b33dd3d876a0f23;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Id71c488586e019260c79018420d61673;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I6c7373fafcfbb14c527e38e0f4440404;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I6f2d4122c89e56e6640df3cec76c3c48;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Ided1b79349f8806da8f5c6898cea94bc;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I37d02ddb7b52ae3495a3a182a3d4708a;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      Id77e3ee5aded95fe141c26ad08639538;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I30b006cb2cf34c967066041123ac3698;
reg  [1-1:0] [MAX_SUM_WDTH_LONG-1:0]      I3c286283659a38021c27b5e5346b59b0;


reg [MAX_SUM_WDTH_LONG-1: 0]                I748f85f6680918a2e992df339b4b6558;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ib0f57837099e3fdf1b908d78bcda4a43;
reg [MAX_SUM_WDTH_LONG-1: 0]                If75e99660e3997f53f7b903bc366f47f;
reg [MAX_SUM_WDTH_LONG-1: 0]                I3253481bee7dbfc0f3eac94c3252ee4e;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ia80693da8182ee2c3708b6ec21d397d2;
reg [MAX_SUM_WDTH_LONG-1: 0]                I7fa3f2648baacebf9e4b59c179601fa6;
reg [MAX_SUM_WDTH_LONG-1: 0]                Id7699f8f89380c315303644fdebacb32;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ibf3e1ead3776901898d4b154aeb61267;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ie486617fc1d6354c7f347692cdbd894d;
reg [MAX_SUM_WDTH_LONG-1: 0]                I7ba403c6745e7d026282ad704e065702;
reg [MAX_SUM_WDTH_LONG-1: 0]                I93cb3974b8594665b2e7ce5593fde69b;
reg [MAX_SUM_WDTH_LONG-1: 0]                Id6a9ab06d58c3a01e1fe04fcf61406fd;
reg [MAX_SUM_WDTH_LONG-1: 0]                I261bd53528b82128acabd405389c8d60;
reg [MAX_SUM_WDTH_LONG-1: 0]                If7fa833bf1b1438e7a5bc783ee745252;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ibb103853fc21f8f3d466ca16557ccd3e;
reg [MAX_SUM_WDTH_LONG-1: 0]                I37446eb66ccfd268cb418655b8160fe1;
reg [MAX_SUM_WDTH_LONG-1: 0]                Id17f6250f8c7f1d7f75fd27f92698da3;
reg [MAX_SUM_WDTH_LONG-1: 0]                I9957b02e8d0d888e6950eb553d9084d7;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ic71258b745437bc8463fb4f847c55e27;
reg [MAX_SUM_WDTH_LONG-1: 0]                I24bb5c315eacf0f4e8c86f6582389e39;
reg [MAX_SUM_WDTH_LONG-1: 0]                I607f203694ff76930cfee4103cb73c30;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ica8e4c56ebb37e189ca8e6b3daafdb80;
reg [MAX_SUM_WDTH_LONG-1: 0]                I7089386c94261e0febf3b4f7dc1aec30;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ia1e4f20f32f7371cb0078d6e80fe8b7e;
reg [MAX_SUM_WDTH_LONG-1: 0]                I790cbca796af58b1726d0a4680cc164f;
reg [MAX_SUM_WDTH_LONG-1: 0]                I0a93f095f9efb1542116a295c0db9c8b;
reg [MAX_SUM_WDTH_LONG-1: 0]                I989ba39f188a44475a83e65a4960d2af;
reg [MAX_SUM_WDTH_LONG-1: 0]                I9bcc1d9b3dd258fa7b6042f0185d48cb;
reg [MAX_SUM_WDTH_LONG-1: 0]                I9ba14715d9f33ef45681ad52f5be9593;
reg [MAX_SUM_WDTH_LONG-1: 0]                I396a897f79b519f4fa02af39d0274f64;
reg [MAX_SUM_WDTH_LONG-1: 0]                I197c0cd576e16ee2197a28c86397f801;
reg [MAX_SUM_WDTH_LONG-1: 0]                I094a178e55425f27ac1ff6195217396b;
reg [MAX_SUM_WDTH_LONG-1: 0]                I3177408f7d08b431be99297fb10586e6;
reg [MAX_SUM_WDTH_LONG-1: 0]                Id4948c876d48bdbf317d32f135e645b4;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ice5ff01d4fb4583898498651a0ac0171;
reg [MAX_SUM_WDTH_LONG-1: 0]                I0fb33a5ced3d15622c9aefa188052e24;
reg [MAX_SUM_WDTH_LONG-1: 0]                I0074e1c3ca0ff903a9201ac5fe7ca841;
reg [MAX_SUM_WDTH_LONG-1: 0]                If65f587e987a51c093e8dd4df532e26c;
reg [MAX_SUM_WDTH_LONG-1: 0]                I33d7e77d08590f0dfb1867e741dd8b6b;
reg [MAX_SUM_WDTH_LONG-1: 0]                I678c22563e0273403b046df4261f21cf;
reg [MAX_SUM_WDTH_LONG-1: 0]                Icca700c12ae2e8155ca6b41e692e8a8c;
reg [MAX_SUM_WDTH_LONG-1: 0]                I5ed74e81d2497681af5a0ca13fe23088;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ic7fa6b8cdfcf7d83d4e101d9c8b7b34f;
reg [MAX_SUM_WDTH_LONG-1: 0]                I26010e26e22d8a2ea831e86fae34a24e;
reg [MAX_SUM_WDTH_LONG-1: 0]                I578efe5c2c504f12c8f2466a7f734215;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ida86d05f907d23ff9fed06927c2ec9d9;
reg [MAX_SUM_WDTH_LONG-1: 0]                I9d9f8c7a23d9750ec44e706bf763df76;
reg [MAX_SUM_WDTH_LONG-1: 0]                I0b41b002a32b8e9e2fe68e819f228fb7;
reg [MAX_SUM_WDTH_LONG-1: 0]                I0e872d4c07169cac84549178fa144274;
reg [MAX_SUM_WDTH_LONG-1: 0]                I6f4ef0f404ae046519b8436171d51e09;
reg [MAX_SUM_WDTH_LONG-1: 0]                I4d04e66ad9103a685fbe088b74517452;
reg [MAX_SUM_WDTH_LONG-1: 0]                I988e525020c1e43d238fad41dab4e6ea;
reg [MAX_SUM_WDTH_LONG-1: 0]                I90d92887cb2526a2956d5e8c9fad760c;
reg [MAX_SUM_WDTH_LONG-1: 0]                I00fe3792cde1eeab36e576fd6634c4fa;
reg [MAX_SUM_WDTH_LONG-1: 0]                I6e586c5ac59a28b30c377e51287bf04d;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ib5dc74106d8841d25a793010fdac599a;
reg [MAX_SUM_WDTH_LONG-1: 0]                I3eaf142d2734d2d0decef084dc037b50;
reg [MAX_SUM_WDTH_LONG-1: 0]                I2d171ad83e27a3745d204849a6f46954;
reg [MAX_SUM_WDTH_LONG-1: 0]                I977f1083f5e4f6f8ac38e2c5aecf1b79;
reg [MAX_SUM_WDTH_LONG-1: 0]                I9bcd673a4293e14fd20b48fa20492df7;
reg [MAX_SUM_WDTH_LONG-1: 0]                Icb7422ea46b22b9330c123b40fe343fe;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ic414cdba230d7ea73972b0eda1ec6b1b;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ie4e1e00503dba189b0f871c3c0810d76;
reg [MAX_SUM_WDTH_LONG-1: 0]                I721c43ab62b42a18c3f5228fc0a73262;
reg [MAX_SUM_WDTH_LONG-1: 0]                I1f7cb03cf806b247be1cace4d75de942;
reg [MAX_SUM_WDTH_LONG-1: 0]                I775cc766b069022bc00220050feee4e4;
reg [MAX_SUM_WDTH_LONG-1: 0]                I08b78f774ed494fa7f119977bd92679e;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ic7dc7f94af108ca7c8003a2d07e1e168;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ibe1327961152cc2d26b3f19476a6e2c9;
reg [MAX_SUM_WDTH_LONG-1: 0]                I5ba97de444af4e8c9744c3b707502edc;
reg [MAX_SUM_WDTH_LONG-1: 0]                I3e4f1314042010b5d7384693b580da7b;
reg [MAX_SUM_WDTH_LONG-1: 0]                I4a47ce6e21c1a274578397e480c184c9;
reg [MAX_SUM_WDTH_LONG-1: 0]                Id184731beb200ad6a53ce273b963bb3e;
reg [MAX_SUM_WDTH_LONG-1: 0]                I3317f2f6eef9a8ef1fe1ff68b47c5d03;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ia6b9fa10c79e6f3847f89b35afb4cc59;
reg [MAX_SUM_WDTH_LONG-1: 0]                I91e98b804ef82eea53c5e8eccfec827f;
reg [MAX_SUM_WDTH_LONG-1: 0]                I5f1e0d0c6b50f70a6f5584124e095501;
reg [MAX_SUM_WDTH_LONG-1: 0]                Id61fcc605b4b581f5d42024c2610c8b7;
reg [MAX_SUM_WDTH_LONG-1: 0]                Id64738b7668931553151dbadd5605b71;
reg [MAX_SUM_WDTH_LONG-1: 0]                I3bdfb451eb96d256da542864d39024df;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ia740d8ccd8230b28d078b2ea3e58d6ba;
reg [MAX_SUM_WDTH_LONG-1: 0]                I574050722f82569d34bc2cfae1eedaa9;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ic8f7ec6ee09fb9ee2467e3cea30a44a3;
reg [MAX_SUM_WDTH_LONG-1: 0]                I2b77d922a74fdcef0d57debc789bd539;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ia1d8127af4944b23475bd7deac91d60e;
reg [MAX_SUM_WDTH_LONG-1: 0]                I247abcede9914633c0a33fc402bf58ae;
reg [MAX_SUM_WDTH_LONG-1: 0]                I1f413d3e081c6aea012b122fc94f73d5;
reg [MAX_SUM_WDTH_LONG-1: 0]                I1b812fb764d3b48511c0d15a7efaea29;
reg [MAX_SUM_WDTH_LONG-1: 0]                I88882bd8a9f8718411564221ad85b223;
reg [MAX_SUM_WDTH_LONG-1: 0]                I232f24e2798488ee66003f3b8cc294c0;
reg [MAX_SUM_WDTH_LONG-1: 0]                I856284e951773518eb6c4232ea7f3d40;
reg [MAX_SUM_WDTH_LONG-1: 0]                I82cbeaf5b3e4796b2aaf33dcbd119f4f;
reg [MAX_SUM_WDTH_LONG-1: 0]                Iaa7791bbc193412e5fe25000ceec23d6;
reg [MAX_SUM_WDTH_LONG-1: 0]                I44bdc0baed3d51ef54ce2728618ad339;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ib6bc7e75ce750a26113cbb8895c2f024;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ib4188380f7e96d5afb99f5045674193d;
reg [MAX_SUM_WDTH_LONG-1: 0]                I5bba219c5024301e420e9a5acbdc5845;
reg [MAX_SUM_WDTH_LONG-1: 0]                I1bb52988c9ba03e16b1b69335d3d7e7c;
reg [MAX_SUM_WDTH_LONG-1: 0]                I1b9990aaeae716f66b0f89fb02be0a74;
reg [MAX_SUM_WDTH_LONG-1: 0]                Iceec2cf6aba9138648a3340390f39fe9;
reg [MAX_SUM_WDTH_LONG-1: 0]                Iad7842f3d4672f42c1064c28d4c8ec4e;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ie5a53cf9343fdcdb5788667c45fadc83;
reg [MAX_SUM_WDTH_LONG-1: 0]                I30e06d190906bc9eb6f1c3156c47f9f1;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ieaaaced47e22029ad2945eac9cc45e6c;
reg [MAX_SUM_WDTH_LONG-1: 0]                I08dc6f8e837b1f6b80bd3fc742290dab;
reg [MAX_SUM_WDTH_LONG-1: 0]                I8eb6a9c907c5909dad6cda98022d70b8;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ia5067b1b458af82c3c2cd50653099854;
reg [MAX_SUM_WDTH_LONG-1: 0]                I198c6753cf12d423c709d1512e66fa9b;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ib600dd8a39fda48d28e1289d44d49a84;
reg [MAX_SUM_WDTH_LONG-1: 0]                Iabf09191227584c76d7fbc634b706d12;
reg [MAX_SUM_WDTH_LONG-1: 0]                I4869ba08cab90a6dcbc454b0001a7a20;
reg [MAX_SUM_WDTH_LONG-1: 0]                If97974406672507f8c9a1c507c4b6951;
reg [MAX_SUM_WDTH_LONG-1: 0]                I4210341f99ac7cb08245137999739114;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ic24f4dbd99c8f4d88c8450d4fef762b8;
reg [MAX_SUM_WDTH_LONG-1: 0]                I68dffa1a13eb6ab54615347729c1d6af;
reg [MAX_SUM_WDTH_LONG-1: 0]                I10153d5548b184b9ac2cecdba4ec4b1a;
reg [MAX_SUM_WDTH_LONG-1: 0]                I104b7f0512440cffc0fcce25e477f537;
reg [MAX_SUM_WDTH_LONG-1: 0]                I18b6758319272eebbe76e1eee5ae55b2;
reg [MAX_SUM_WDTH_LONG-1: 0]                I780263b10b98f9bb0eaf66c045d8d37c;
reg [MAX_SUM_WDTH_LONG-1: 0]                I37b772442e55cbcd44ba892a0608d662;
reg [MAX_SUM_WDTH_LONG-1: 0]                I0ac256a6659ff5c6673fd110a8bf578f;
reg [MAX_SUM_WDTH_LONG-1: 0]                If134e1d27e736005e5a390e7a2ea1f4b;
reg [MAX_SUM_WDTH_LONG-1: 0]                I7b37b8f908cd82683832536e02faab0d;
reg [MAX_SUM_WDTH_LONG-1: 0]                I08b4bf60c9c7e7229bd1952cc88bc7b3;
reg [MAX_SUM_WDTH_LONG-1: 0]                I267d637eb63fef9f4723f7978fad88f0;
reg [MAX_SUM_WDTH_LONG-1: 0]                I4fb56a70e5ffa71f58f715da36368e04;
reg [MAX_SUM_WDTH_LONG-1: 0]                I5e9e2acb258baf96ac4b525bba54a462;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ic40f61443a4d8f87769067fc39381cb3;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ieb36710c9a3726f33407436d62639c8d;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ic804af393da2e4b9c8ef25d4a3b4e8d5;
reg [MAX_SUM_WDTH_LONG-1: 0]                I52e4c446693c29a42bb3b665f72d382d;
reg [MAX_SUM_WDTH_LONG-1: 0]                Idbf02cf10add496d30fa44bbb18458c6;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ida095585ad26e215f1c1bf989912da89;
reg [MAX_SUM_WDTH_LONG-1: 0]                I19f1ffa05c7c9a0df5e7014044024c7b;
reg [MAX_SUM_WDTH_LONG-1: 0]                I4d68a2fe778fa93faac38b138138291f;
reg [MAX_SUM_WDTH_LONG-1: 0]                I54393ada6f76ac82c31f2668e228e29d;
reg [MAX_SUM_WDTH_LONG-1: 0]                If5b9ef84f09680f3593250b13a852c1c;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ibb759bc4179e5b7aa759d850c7cfa467;
reg [MAX_SUM_WDTH_LONG-1: 0]                I05e8b5f8b83f07b609b5ebf272bb2229;
reg [MAX_SUM_WDTH_LONG-1: 0]                If6ac15373ec1146d38e7aeb71c3ece64;
reg [MAX_SUM_WDTH_LONG-1: 0]                I2ab3675e1eede757af80716ba980a4e6;
reg [MAX_SUM_WDTH_LONG-1: 0]                I388c271687ab31b57421ad57192273ed;
reg [MAX_SUM_WDTH_LONG-1: 0]                I6121679cec8caa51dc5ff0d1a61f9821;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ia0649b990bf5716cfab230127cd5d47f;
reg [MAX_SUM_WDTH_LONG-1: 0]                I867a0626ca22108b16267d95c0aadf4f;
reg [MAX_SUM_WDTH_LONG-1: 0]                I1af54bcb73d7c6b93e55450871207976;
reg [MAX_SUM_WDTH_LONG-1: 0]                I91883553543d0425e9c6dd726dce3d27;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ie95405659701278e3f87bf1f823a037b;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ia42392e2104b50c0908aad82738a5ee7;
reg [MAX_SUM_WDTH_LONG-1: 0]                I68ad63230a51b9b9e3daffb307ea970d;
reg [MAX_SUM_WDTH_LONG-1: 0]                I7a052d63944ccf42e598efe3a95b88f8;
reg [MAX_SUM_WDTH_LONG-1: 0]                I2b3c6d69f79c8d51e4d1614c62c44fcc;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ifcef0e92f50e3920bf1208af5d64c632;
reg [MAX_SUM_WDTH_LONG-1: 0]                I111340a19625901a3c1b95fd0bd1570e;
reg [MAX_SUM_WDTH_LONG-1: 0]                I11aec4fa85c30f6fe1fd9fa72542ef6c;
reg [MAX_SUM_WDTH_LONG-1: 0]                I80cc333c181c16a96b7bd6501c27c2b3;
reg [MAX_SUM_WDTH_LONG-1: 0]                Idc6354325a6280ae9890da33c06c33ec;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ibb04cf82acc4ac16599ad3ddb0c2ada2;
reg [MAX_SUM_WDTH_LONG-1: 0]                I3ed096dfd8a14f4acb4d53a70cf8aceb;
reg [MAX_SUM_WDTH_LONG-1: 0]                I0fa07f95e96326cb0599c0c3f76e2b48;
reg [MAX_SUM_WDTH_LONG-1: 0]                I87d98fbc97d9a78c2e7d6a6280e7a49a;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ib7ddc4dca877f7cf5697a02c3d1915ba;
reg [MAX_SUM_WDTH_LONG-1: 0]                I3612ef280891f6017fad205d0484bde7;
reg [MAX_SUM_WDTH_LONG-1: 0]                I561547649aeb5b4c3f10d9506db1f3cf;
reg [MAX_SUM_WDTH_LONG-1: 0]                I84cc76c0079b86da7b994844c3ccb875;
reg [MAX_SUM_WDTH_LONG-1: 0]                Iec013c508d0c6401d7eb856e7eb60446;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ifd8979aac6b6b24aa560b46b18240e92;
reg [MAX_SUM_WDTH_LONG-1: 0]                If12394e78dc913b01890b56650856a44;
reg [MAX_SUM_WDTH_LONG-1: 0]                I94d18aa10695f3f22b23246884b72822;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ic90b38835dd7e760dd54067b196f8470;
reg [MAX_SUM_WDTH_LONG-1: 0]                If3691ea51f6efe9b165a31964854d2fe;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ic2ce582555add38a14f5006d3c87eb15;
reg [MAX_SUM_WDTH_LONG-1: 0]                I58cc950ee2cbe56b7c5a619be3792511;
reg [MAX_SUM_WDTH_LONG-1: 0]                I0d8e329ec5873db96df1ec309445a096;
reg [MAX_SUM_WDTH_LONG-1: 0]                I106325488e2ecfdba1cf9e5201e6bc8c;
reg [MAX_SUM_WDTH_LONG-1: 0]                Iff73a0085541a511d3912b64686a82c5;
reg [MAX_SUM_WDTH_LONG-1: 0]                Icdab59de68f2870504598c9ea18f1d2c;
reg [MAX_SUM_WDTH_LONG-1: 0]                I75604d727e82c977741f90113719183a;
reg [MAX_SUM_WDTH_LONG-1: 0]                I6f50c4d0d2639857b2dcca300c2d7b04;
reg [MAX_SUM_WDTH_LONG-1: 0]                I5cd013a2be2e761c10c6a957632517de;
reg [MAX_SUM_WDTH_LONG-1: 0]                Iafeedddd02428bd2610c576e68d4ae25;
reg [MAX_SUM_WDTH_LONG-1: 0]                I912d6325e34180e0f668f0f024e63581;
reg [MAX_SUM_WDTH_LONG-1: 0]                Id1e05294dfd02df499ad0c08bb5c191b;
reg [MAX_SUM_WDTH_LONG-1: 0]                Id3bb9b100ee4302473b49ac14615e9b0;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ief32db1cfc443119b6202b0cc7bf70a2;
reg [MAX_SUM_WDTH_LONG-1: 0]                Iad7dbe9909b5eed3261adf92d3813acc;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ie7daf0789c35caaadbba06cafabd2b70;
reg [MAX_SUM_WDTH_LONG-1: 0]                I2bd1f9b75d9ab94af9ddceb7528935e8;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ic3d9f5c6677758810e4865779ec303e3;
reg [MAX_SUM_WDTH_LONG-1: 0]                I00af04882a25e2832d913a67d4d86d7b;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ic9db631df0a1a9108c10c3e0eca7bf15;
reg [MAX_SUM_WDTH_LONG-1: 0]                I749f9ed1fb2dddd40ebc28f638e02935;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ia45b2a24df24bd5e3c95885c8928686c;
reg [MAX_SUM_WDTH_LONG-1: 0]                I7427464fde340780aba7f9847b4ad564;
reg [MAX_SUM_WDTH_LONG-1: 0]                I33fd1ae225e2b881b2b41e0358675e22;
reg [MAX_SUM_WDTH_LONG-1: 0]                I2e21a35d1cf560936fd19b944a208b6b;
reg [MAX_SUM_WDTH_LONG-1: 0]                I249522a3d42cc75d7a6b9ede1222ee76;
reg [MAX_SUM_WDTH_LONG-1: 0]                I68b4c43d9f40ae4bfd70d2983594392c;
reg [MAX_SUM_WDTH_LONG-1: 0]                I63145e0fec15c7e7c0de105f348bfd31;
reg [MAX_SUM_WDTH_LONG-1: 0]                I8af625de86c04016c3424d116fddab5b;
reg [MAX_SUM_WDTH_LONG-1: 0]                I54c9c10527f83b4ee4e1e22f1e4044ed;
reg [MAX_SUM_WDTH_LONG-1: 0]                I972559e47c7f83bd9000ca1cfc14d8e0;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ib97a7f941eb7ce2a867503a04ff86a67;
reg [MAX_SUM_WDTH_LONG-1: 0]                I5979b55f607c71017537f2b48b40cbea;
reg [MAX_SUM_WDTH_LONG-1: 0]                I6a56760b621f238843b091279c69897f;
reg [MAX_SUM_WDTH_LONG-1: 0]                Icec45bf76c241d37c9a50a5cd092da9d;
reg [MAX_SUM_WDTH_LONG-1: 0]                I2f6d3f61f2890e584d3063a09587e99b;
reg [MAX_SUM_WDTH_LONG-1: 0]                I7c396ea2e959d84fd9a6964617cb29c6;

reg         [ 0:0]                   Ib0973b6e90e7678addcb064fded7ce0f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5033323484d90d6bfbe03749019fc6dd;
reg         [MAX_SUM_WDTH_LONG-1:0]         I97afe24956b7f87cd431f048202bab67;
reg         [MAX_SUM_WDTH_LONG-1:0]         I117235e3ac8e68e4c1ab34db1612aba0;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifd700cc9d18f99b63f1947f3ae631976;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifffbe3d1007fb07a20d3b37902b3ec95;
reg         [MAX_SUM_WDTH_LONG-1:0]         If5443777169422ea6e1e3f709b970e05;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifaf9fc93e4609d818aa46751754c17f1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I419caf964986c655df84d043badc37c9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3095214ac0e6c1323e75ee4ec85e6821;
reg         [ 0:0]                   Iee06707670e19a82d911c1750bcfc811;
reg         [MAX_SUM_WDTH_LONG-1:0]         If5dad13ac41b3034bdb034bc86c9b348;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ided9739bf63937933250a6d0c37535f9;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id0f139b9f3848b45554ac8429230eea2;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id9feed58cf9565255abfd0bf7e3ec068;
reg         [MAX_SUM_WDTH_LONG-1:0]         I30a3be3b5f6ad1880a917eb35659a1bf;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie8148d9aa962a733eb65877b902a187d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I69e98cf3e679183aef6005bb582b18dc;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7f42a504fc61c9548acebdd8b1858eaa;
reg         [MAX_SUM_WDTH_LONG-1:0]         I08b1b4639b5a9ca509b943b977f6d4bb;
reg         [ 0:0]                   Id8d5df9e869aaeb107a41a6bca3b89bd;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iac428f9f798618e1ef495c626c41892b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8d7296627d886566783e79c01b9fa423;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4fc4c97229a8b1f631a3b505941159e4;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib9b16bf51891c328dba2699eb9bcef95;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6c30501ec81fce286817788d614a7824;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia4d4f37baec48121a88808075dd655ef;
reg         [MAX_SUM_WDTH_LONG-1:0]         I385495ea2bf6442a95ab7561456254ac;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5128e03d383c226befa6f7422f3a6f04;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib208908bab4c20713cd17e20139c8db3;
reg         [ 0:0]                   I507f8602a99a1096e4c293ba3c235bbb;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5a6427c8f18b36d2ea18fe60a0831ef1;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id939992b99a11c09f4688c10ca1a34d1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I823453ccb90d5b2b2d9dfc6e8358224d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I279c5c00b92eb1b872b5afa168b0306e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I66f25b1c3c0eb226295179adcca2c3d2;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3068627e91b667d14cd3e55a9371931a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I44c4e0a2d8a7289f8660b81a9ecfa19b;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibe868e258dc87f0dd1460ba6b8354671;
reg         [MAX_SUM_WDTH_LONG-1:0]         Idc3083c3021200345e3edd35a9d4725a;
reg         [ 0:0]                   Ibdf2178bd18783c4797c21e642388d16;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icc29441eac6ca7a138d45743d37505e3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I320d4f19a5b18c23ff407508d47caa77;
reg         [MAX_SUM_WDTH_LONG-1:0]         I16becf3c92615d98d5ec51ee9641cc0a;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifbfacc3b3a0128119943bcbf80176612;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6b4f670c9e8e25984e8891f2440322ab;
reg         [MAX_SUM_WDTH_LONG-1:0]         I19bf0990a30c72421f231772b8627e8e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3ec3eb096ebe3ee8a47e1cba6487b997;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7379ef16405c461ac44b66c4315df831;
reg         [MAX_SUM_WDTH_LONG-1:0]         I79db45b23d21d533a1f9a6e8f94d403d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0979534730cc2b53547d413dbb6b75f4;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5aa2f9c0667d1a6e871efbd4d2bad3a8;
reg         [ 0:0]                   I2c690809d9b9e3482fe5a133b5c00afa;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0e7754dcbc04a4850e052ae4a2fbe328;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iadb28dc990ccf2dd3099544de16b8f16;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1f71aebf698788d6ada66891e9ea756f;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib234e9cf7e7616a1ebc6ab99df2a7ccb;
reg         [MAX_SUM_WDTH_LONG-1:0]         I297d1edcc583ea4d69da780150f0620c;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib0a717cbb4fe38a3fc85520ca0826fd9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I037ecd5945b1f1280b4469d73fe1c7ff;
reg         [MAX_SUM_WDTH_LONG-1:0]         I367ff6b11b884e02a3065fc7fe811e15;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6fab19692b512166fe9c74b5e987788d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I04dd73af505f618ccdb209b3cf97ceec;
reg         [MAX_SUM_WDTH_LONG-1:0]         If8c559905d4120488d431719c4e8ce24;
reg         [ 0:0]                   I369ffa98995ba0834f8029ecce705c56;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia30c019ed8ce395556494a92e7b42a92;
reg         [MAX_SUM_WDTH_LONG-1:0]         I20ed4f6f14e20ce3f0e106d1b7782fcd;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib10626ffa126188c5bf1fc8399107b26;
reg         [MAX_SUM_WDTH_LONG-1:0]         I29007c52357ac7afbda39d72a5bb60af;
reg         [MAX_SUM_WDTH_LONG-1:0]         I66d367c046611f145e607a90911cf499;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9c4c2556f6170a8df61d909855a846ed;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6fadc3e8d995bb4317bf7b4377c3c2c5;
reg         [MAX_SUM_WDTH_LONG-1:0]         I99b20e911c189e0616f02376ab736e91;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5793c12f5dbdd8245dbb202d550ca960;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id0660e9637cad1ce1a73d37188060154;
reg         [MAX_SUM_WDTH_LONG-1:0]         If5a7af7ca023e1393526e888f4220a44;
reg         [ 0:0]                   I9ccef4c47ae7cfab43584de0f2e193d3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9799695ea8244992a6694eaf5c8ae64d;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id043eb50634e803e53adc1168379a5d0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1f866dd0b129267550aea1a267d9c91e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8c4da05c08210fe33139c3d3e5d75d58;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib41f7b823681fdd084b6d8436a407aa8;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic5b50a785b7acac7e3be4095aa92e50a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3ffbe03796b66d00d47fd918be60ab89;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifc92a916da938ef6164db250be635f88;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8ccd42508ce7d5bd897c2cf0c54caeb3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4920e7e82749cc036b58a7cd0a03e327;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie1040b2aa91f272e4449c4b5f9f8f575;
reg         [ 0:0]                   Ief31fe169c1b360d5933558208dbb602;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4524cd664b4cb41f642c675fa484c84b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I65968fb0f63d52ad96cd8fa270126a1b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I839ac8ee59f51d4c3de92ba5cb26e788;
reg         [MAX_SUM_WDTH_LONG-1:0]         I33cd95f1919318a0f3df5df7310d64c6;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4933e8d16fba26cd797b25a9ac2a2de8;
reg         [MAX_SUM_WDTH_LONG-1:0]         I218f7578eb748e31d0002052f30c5842;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2a808d1c42ad758ae3baaaee8129dfb2;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4e851fd3c114af87f5e8c68c02594e3a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0da40f88adc46e90f616acdcdb8e0e2c;
reg         [ 0:0]                   Ib8c0317dafcfb91b3da5eb5afae1f2e2;
reg         [MAX_SUM_WDTH_LONG-1:0]         I64e959d80af111ed2fcd54a5407d21bf;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0dee7767e472a5fd71250ae6c57cc8b5;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9f40be7552b3dd625e5bce0befc5a548;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8fdf98ffd757c8845ed6ffa4ddd1a16b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8103b777314a4fa471e0898fde9cde08;
reg         [MAX_SUM_WDTH_LONG-1:0]         If6c3ee8e0d7dea58043d5be0f4630873;
reg         [MAX_SUM_WDTH_LONG-1:0]         I711a5171f591f472cdbfc9a0f5e1aa17;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic30bc38184dfbbd694af52640692709d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I422f6fd1d273a3834d04b04ab8e2812d;
reg         [ 0:0]                   I54e3f08f6f4cf784da57ac39f246b8fd;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3e0da4bcbab4804b5397fb3aa2c94f51;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia0fdc60b90ad18b6585ec1ad4e89e80b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7809fe7a30d041a7e569ffe890242df8;
reg         [MAX_SUM_WDTH_LONG-1:0]         I672b14ec1b3c4797545f266727505a85;
reg         [MAX_SUM_WDTH_LONG-1:0]         If9620d20ebaae6245a2c386d9bf5fdb1;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic74e22bffd88f32eefe499cde0fafa8a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I76d38ce67387bd76ab45c9cba7d18b31;
reg         [MAX_SUM_WDTH_LONG-1:0]         I44413c6f6f6493f8a86abf6eb32604f6;
reg         [MAX_SUM_WDTH_LONG-1:0]         I67f632fca617fe06565ddcaaee8fa8b8;
reg         [ 0:0]                   I16c7f1b874b0d05c6d120bbede254416;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3740b30d31f3c61d93a14a46e3199c4d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3fd38a71ce6aa3db1d7a5a9f8a991e12;
reg         [MAX_SUM_WDTH_LONG-1:0]         I63e5718bf7d8771ef90b91be73d73264;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie385e1aeb2b0dcf6d2454be3d7708b27;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib2d1b7e105b25b492b45da72536d7578;
reg         [MAX_SUM_WDTH_LONG-1:0]         I588abf5ef4c583f0fec422736a0ce6a0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I58bb95c56c7be17c263a2161210d7d8d;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifaf0e1f21b3bd7393c475b5126540a72;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7027db9e0450724a6d417d708f1043f2;
reg         [ 0:0]                   I0c3cb2de514ecab0dd311e86a4dc3cdb;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibf0a30abfec9031737eada436ac1a0d4;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iebcb7206d8860b5094459c5d10b4efed;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6bbf2b47a7dc50e66a3d8d258d6e31fb;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8459abaa907f5afcd11884b1ec8c06c5;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia16ae2f6ef5000d47b6b84ed058252aa;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ica32690dbc9ea110fefdce92260b125c;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic431d9383cce30b1889c92e2be4cb9d0;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib9cca4c0e58373c26d5fd9f51f793898;
reg         [MAX_SUM_WDTH_LONG-1:0]         I99bf0bc8ac20832b3724b2753f6ca449;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie701008f3c60c51ed72c5f964a8fc36e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3e2d78f8307a1787f8b2eccba94c7557;
reg         [ 0:0]                   Icc5ba4554d7a44bc3b43377efbe3b5f8;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id36e8953a02400a5ab1f4dfdb0422e6d;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic1b4444ab0df9745d29bf893d9b83168;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5f52dbf600656a8f5dc6b6b8a45ccebe;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7f307af79f45ad4b9511e3961c917078;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie17a5be2a16d2efb98c976d7ee882535;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5f19d2adff2f34a4bebe03f929a09c49;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3cd69aeed9e869a2096d6dced5c209a0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I359b6a22c9568a13b81670c741281393;
reg         [MAX_SUM_WDTH_LONG-1:0]         I24ba99614df383c38bbac50ae8b4487e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7498bee46de6b1c946ce95fdcc89f6e5;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0f644f42cabf871b71e5a82871bc7b5d;
reg         [ 0:0]                   I5e51f49adb6dce65a9f19ff736526c4b;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ica71108a53bfcfd1892b4d03ef68110c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I71f9e059726a6cac8bdf0efcc0eadd2b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0c9b2c1da30bfab514bbb556ae7bd4c4;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7918b2e37e96aee94fbccca7e0f75fc4;
reg         [MAX_SUM_WDTH_LONG-1:0]         I76eebd77eb77e0abcbc727d2c511370a;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibb2288e62110bae5b2d3fe901974e5c7;
reg         [MAX_SUM_WDTH_LONG-1:0]         I080f931dfef9d8adfb1dc1ee073eb64c;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ide1106431e3565158bd81ccd6b18f3a1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I63df19931e8d28666cccd79922cbd418;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9a7e4a59447048de90446f877eb06627;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0917e92ed84363ca92fd2074acd74eba;
reg         [ 0:0]                   Id57092394c7cda397f42374df4aa3fec;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7c97629ec6e594f9b2160815ddd133cc;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie3eefdf7b5561a90a6ddd9e6aa432509;
reg         [MAX_SUM_WDTH_LONG-1:0]         I56eeb10d11e886cff629457a640a1c76;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7a9eea89c4e76d856df44b6bdc332840;
reg         [MAX_SUM_WDTH_LONG-1:0]         If8d8f4333e893788fcb9ec54256e5b7a;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie4af0e7e04778d85f5dee73da33376a8;
reg         [MAX_SUM_WDTH_LONG-1:0]         I019a4e997adf54f5f5ca651f80b7901b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I10294667f09abbfd4e2f757c414072fc;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id4e8ab8f15b36bd27d1e4ebc5cbe1495;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6c93588ca9e7c623d75314da39e89a91;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1020412efc78d12a9ebcbaeb83e5dcea;
reg         [ 0:0]                   Idd6a4f8ae94c431f2fa3312b4fd287ba;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4823c8239ace86dc399e906c1b5a0d74;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id0b574f35a83dcfd4481a10043cd1884;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifc577e5c2c7288373a8c5e3969ac1589;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id18a1a17c1cf6e8a2492aa73b62898f2;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id8ce8f636723b9f119bb86c25017e6b3;
reg         [ 0:0]                   I9f1f8590dcf596097bc81001d51684b9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I10ad572ca72c2ea991487c39f7eabd7b;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic29a18d8d504a2d5280c1d7771346518;
reg         [MAX_SUM_WDTH_LONG-1:0]         I96a79193aa2956b8f901d5fcc9cf65cf;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8c97a246c749fbef029f8b1671c772bd;
reg         [MAX_SUM_WDTH_LONG-1:0]         If9ba9d221909ce7499725f6fd7d519f8;
reg         [ 0:0]                   Icecd765baa87877675b0f3972d78c02f;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie9f3fd3a6d16316e55addbe0e336519f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I53a7878f44253f0f1a82d9d27b1a44c3;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie0e928125f9d3d17d123d97e00f1fc34;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2bd0f77efeca09eebe82ea234e9fe638;
reg         [MAX_SUM_WDTH_LONG-1:0]         I94f2e7ef9b3463bd598dc9049f6fb0ef;
reg         [ 0:0]                   I401a38ea1d71dcc71d17a4694ceb0988;
reg         [MAX_SUM_WDTH_LONG-1:0]         I07965bca84276dd56da1af98e64b0adc;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6dc16510af6b61b79b339d0fce77ac24;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic655e213ab81f5d61a018d3ed7016b12;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2ffc4a604025a2f5c4e273c1d070a725;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1c76818a9a3b688ca897aa479f7d807f;
reg         [ 0:0]                   I3db9b61e28a51e974e2d5e323ad53c1e;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic2ade31b8bcf68c4dcc1a371ff14074b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3bfee9d3d88f0569010a4e0101200c19;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5d4738755a26beb6d0f61dd3dec0f804;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2f3c800091275bcb72d1a2a38fba53f3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I378e67cca7c4ff6325683f8346963210;
reg         [MAX_SUM_WDTH_LONG-1:0]         I04c8915a7f4bbde003f7facc84435c1a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3f50b10072f38b6addee6845e6df9118;
reg         [ 0:0]                   I96d0a4387f9b959bc779ac13351182cc;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic0edcf240048fbfde4e938c3e4c5e281;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icc60eb18ba740036d2a17f98f15cfb98;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1677daa18aa8b226753b1a887b9420d1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I36bc2d4c9a4480daa9b0944c08b50738;
reg         [MAX_SUM_WDTH_LONG-1:0]         I38419a6905f50135a6783aacca0384dd;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib48892dcb0715987289662a14672611e;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icd9c94f929dbc71c9b836fda3019630b;
reg         [ 0:0]                   I64082bc75fdbeb69a52a4361ed2d5883;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8b42e89ff5f780d4ef8cd1cd5c99ef61;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5d0249d9a772805b3fba3f3c7f5d35bd;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie97341deb6fb24d49eb8b96bd0fd3f35;
reg         [MAX_SUM_WDTH_LONG-1:0]         I17dd788f9d8e91307b6b1ab7488f9ce2;
reg         [MAX_SUM_WDTH_LONG-1:0]         I92ae370022ed107b152b10fd0aa3d2b7;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iebb39f0d19ec1208bbfba6cf67a3bfc7;
reg         [MAX_SUM_WDTH_LONG-1:0]         I81861f6bb8bbbab6e93407cfb4a852b8;
reg         [ 0:0]                   I62929057b7c214bd38fd532e20ba5623;
reg         [MAX_SUM_WDTH_LONG-1:0]         I70b1b8521b36920707e95fc9418eb8a9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I217b2e3ca0a534fc5b1910adf3c1b57d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8429b08891dc56af24c72ce1b7725457;
reg         [MAX_SUM_WDTH_LONG-1:0]         If96747262303f6c5c6b129e39224bd23;
reg         [MAX_SUM_WDTH_LONG-1:0]         If7012457af15c405baeaa1710319b541;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia0a0229ef71b85195352bb664ea4e4e3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I42aeb7c23accc2ca874c7f8221c3af93;
reg         [ 0:0]                   I641179f37fef63e7deec603b3291381c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4fb1c32a62cbbaeb585c6564a3c938f9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7df6a95bf51f40693c439c6df36510d4;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8fe65f9c344d7ec8657f192abefc3fb6;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4d75c95d34d8d8aeeb528456bbe136e1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I43746054a38c9521f8da9db9d0e91f99;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0430ac2a4b2b2e2fc7f8154bf946553c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I25dc807fd55b81c9f24fd0d1edcaa758;
reg         [ 0:0]                   Iff04b7ec87148f5bd408b4ec4b0590a5;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iefc37daeec14e14ef2fe0716f73109dc;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7881184f1779b9fd4fdf329c5f7664da;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8e6de2d692a307ee8a5a4b2a9265a633;
reg         [MAX_SUM_WDTH_LONG-1:0]         I54b2b18ab051b468808a3d0fc4bc893f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I37ee86e2ca32832862cb57efe76bbedf;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic95f2fc697574803c0f7fa35c2609f0c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I933a30c52c9bec5172530b2d739a3b63;
reg         [ 0:0]                   I198bfb18d6f91c8f62777e6f592a88fa;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibd15f164f6d2ac9e5721a21464bc2c5c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7bbd7df18f85197c22fe8cfe37312af6;
reg         [MAX_SUM_WDTH_LONG-1:0]         I50d5ada7c91c7af16492c6b41151b68f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I32c8e7996b3473d4906c40018799a16b;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic0eacd5a4812ad7ae3fa251ab2db4694;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ideecf8ab87d28a840cd93851169ab05b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1ac6775eb38457b7962241d2e7336b0d;
reg         [ 0:0]                   Ia1562c88b4f56d8935c3a5d6ead0f816;
reg         [MAX_SUM_WDTH_LONG-1:0]         I951dfff9507bb70214d48e03a0ebb3a7;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2ecaa89698604fddd863d7e28d643a57;
reg         [MAX_SUM_WDTH_LONG-1:0]         I273e0fe9c51c8549c8dfff393ca2e4e1;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifb1fc76002f6920a1f44c7b1bbcd0020;
reg         [MAX_SUM_WDTH_LONG-1:0]         Idf6d4e3aa753aa396a9bffb27732f851;
reg         [MAX_SUM_WDTH_LONG-1:0]         If14ca1f5d1c2977f9da79eaebaad1bf9;
reg         [MAX_SUM_WDTH_LONG-1:0]         If8f1505d9f10e30bd3320f500d34932f;
reg         [ 0:0]                   Iaccba3030d9d9f8a56f86d6e34ed6325;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie78e30b2a2eda75d0df7d10fd67b5e36;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id32aa77c6406b35a00168bb5452b12fb;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9a73686acefeb361337511f6943b036b;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib6eb7ce5a070f3a87bcf0e18be8c855d;
reg         [MAX_SUM_WDTH_LONG-1:0]         If69b0b717c35d33fc8c0e59b07eb9edc;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibb0d73078b779585e6b0e228391ecb96;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2894546e399fe3e33d7579772a1310df;
reg         [ 0:0]                   I953dfeeacee8c44c08d0a425fa549e49;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia0b83a372dd4115dc4d61eb8ff0811b9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I97f99a266267859aed199b278a430417;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie18cc792329941a3654322376a937d8d;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie914a99f08d60b74c3c36a632a4ca9b0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I82916e9dc3894ad88e12de01a68d6aa5;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6cbf576b3d652e34c0221f8316b5a392;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9141b2516d7f855cd186472780af7b67;
reg         [ 0:0]                   I214a50bf9f879fe747904f4679fdd1f6;
reg         [MAX_SUM_WDTH_LONG-1:0]         If5c5bcbbea01aa22f242b913f0d01929;
reg         [MAX_SUM_WDTH_LONG-1:0]         I07bf32ed72de9c02abf700c64853af61;
reg         [MAX_SUM_WDTH_LONG-1:0]         I52663a2999fb9571834d517538691b6f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8dcb88c94506367aabe8d7ed62cc56c2;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie676a4bee61154145391d9cc473fe91d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9502c8fbf6b48749bf9f84a89a937dfe;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0c91e540e7106f32ae59491d8ed1853e;
reg         [ 0:0]                   Ic88f2c344a8ad254fc7d7034cb594f6d;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iccba58cd3519fb4cc75a61b50da1d562;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iddfb8a8e261389eb4a2a10880c19446a;
reg         [MAX_SUM_WDTH_LONG-1:0]         If0d55f861d4b3f0970c529024ca142d5;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib054f5d3f5cbb29a053d0e50c23cb3a8;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1d65e9f97e93de8cc2a5dd532f8e482a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3bdeab8c87325d46e45d9e2d44756934;
reg         [MAX_SUM_WDTH_LONG-1:0]         If9228f7ecf19c41f4bbd8dabd0d5816c;
reg         [ 0:0]                   If299d1a4e044acbc70bc3b7bce9f86e9;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibc0999e4d0b3cc2650f9348b8c204b14;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9e3edee214c4937d2aa462d3cffa624b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9fcbbd2e81b006b50e2d35ed2627bf83;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie16f3d50ad5e5581ca099549db7232d2;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6345e93f3fa7f5eb2008dd41742afc2d;
reg         [ 0:0]                   Idb373d2cf788f6a93a0e5df7f9179292;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2aeff1fb4b839a581acaf26f90f9113c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I698b93e10073b5d29357cde4bcac9dbe;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie7ced910d84655790823e6173a5a314a;
reg         [MAX_SUM_WDTH_LONG-1:0]         If6e3b6fd1810f6964e9024329d7cb3e3;
reg         [MAX_SUM_WDTH_LONG-1:0]         If1045908c6d7476bd5507e57d08c406c;
reg         [ 0:0]                   Ic73b8c8f76a985330d4ac1fa0cc28e7f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7d60d53f883f8187700c4e78b4c22f1c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4d4f6705ed77a16ff31b34bae0d8b6d9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I70a492396580ac1143d8a2f4b181e873;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2fade32b5bdf245fa15289620dae2670;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie0dc166f57fea074496241a32cdb6015;
reg         [ 0:0]                   I134dfb2c57d8cdffd2789e2f442c3247;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id6fcf4b7af4a37c854a12e2ae80851fa;
reg         [MAX_SUM_WDTH_LONG-1:0]         If6a2518891412caa6d6d507082501f1e;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic9912e5a838a377b26a19d22148a64df;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibc0fca22d16444bc17877106ca772c31;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie4291d233597d5d676a80fd62d9bd208;
reg         [ 0:0]                   I0c735e43be8030078ec10bdb6882e79c;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifa5e5f7d753964f14f0f16dbe552fd85;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifc13b798d76aa70ec1877c275fb31d36;
reg         [MAX_SUM_WDTH_LONG-1:0]         I57d6637f0bdab578a790e4a12ccaa16b;
reg         [MAX_SUM_WDTH_LONG-1:0]         If8ea04fe685b4f20cdaf9a84984d56fe;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie0c86f20c28bcbe410b191b90d29bf76;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3dc5d3f66726e15968a70cbf3d3b656a;
reg         [ 0:0]                   Ie9951415c1d599570af1787767caa2dc;
reg         [MAX_SUM_WDTH_LONG-1:0]         I900d471b087cf5a436c2ad66a84d8280;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id674686e7ac37fd6f63846f9a9cede19;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie2ed9668d13d219c60f2e0614488cd42;
reg         [MAX_SUM_WDTH_LONG-1:0]         I98abc995ff89934534543be93c6e3ffa;
reg         [MAX_SUM_WDTH_LONG-1:0]         I579cf9386ab7b08efa204d735335e462;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9efa4d729d10a6b7cc335fb765ed032c;
reg         [ 0:0]                   I2630f187d63ba9b0af52c77093e6b760;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6d1434907f0292ea2ee47cbc5b52bfb9;
reg         [MAX_SUM_WDTH_LONG-1:0]         If9191ebc8e88d4e75f0f35897ebb1421;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3511287cfe69d5cedc5a8fbcad708437;
reg         [MAX_SUM_WDTH_LONG-1:0]         I91812179d44cb675b90d477f33ec48ad;
reg         [MAX_SUM_WDTH_LONG-1:0]         Idb04a1aae91fdc477ca38ed66789ee88;
reg         [MAX_SUM_WDTH_LONG-1:0]         I566054aece562960590ee28b157e4a3e;
reg         [ 0:0]                   I83db667ace2f04ef4950e2c186e0e6a4;
reg         [MAX_SUM_WDTH_LONG-1:0]         I938bef7ba7ae1739d8e6a6a7c117a1b1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7b2ffb762cd9ef7aa8ba224efb75c46c;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id90bbb642b0f4434d8a148a28b6b2f65;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia4e297e35d484b15adce7e1d67f582b0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I84996b1d03b692f6f736fb04c7f91e83;
reg         [MAX_SUM_WDTH_LONG-1:0]         I83078cc7857fc17b30f640854a4d6be5;
reg         [ 0:0]                   Ie818c5ea3f3b879fded32e6cb06ca546;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6384a9416b2d1da01df1b2d7b16c5390;
reg         [MAX_SUM_WDTH_LONG-1:0]         I94bb467129904032736fb13dd636c600;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifa76758b50f439170ecd6d86ff898bc4;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9d831dd976e8cd5d8f6a6818601e6424;
reg         [MAX_SUM_WDTH_LONG-1:0]         I474774ae149804412ed4aaf1cdcaba88;
reg         [MAX_SUM_WDTH_LONG-1:0]         I964cdcb4e6b49a62d30c2a2540851317;
reg         [ 0:0]                   I3a67a175863091a52844aae6ad277da0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5097a79e7cf7a30d38ba198d1407119c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6df268bc9f85ce88674a9165664ea84a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I74fdcbe9f49f7bce1f5e31d956c5883c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4a1b8453cb7a21745d5f74ad05653ed2;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9c53b478b2011fac0615a152fe60d5b6;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id75dbed8f1a5befda32c60b994681013;
reg         [ 0:0]                   Ia3aba80aead67feab12e4800fef82322;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib113c26c8dcf49c972c41a938059a787;
reg         [MAX_SUM_WDTH_LONG-1:0]         I378a59323b74623c5524f854d6e11226;
reg         [MAX_SUM_WDTH_LONG-1:0]         I080bf885464a0cc948a4450e9f7d1d26;
reg         [MAX_SUM_WDTH_LONG-1:0]         If769e73adea227de1fd85c2e89d0ba08;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifa6a34b83225e9d9b28b14874c4444e3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I584b1d4d6fb7ee4f20ad9c96715cdf90;
reg         [ 0:0]                   I1181d42b560fca7bb5c924a81a5db1fc;
reg         [MAX_SUM_WDTH_LONG-1:0]         I970c4a25a8bce82a9d2846679029fcab;
reg         [MAX_SUM_WDTH_LONG-1:0]         I265f9b91fbb62164e589dcf96818c4f5;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3d59a47c88227734cf6fc0d6fd30db11;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6144b6df2c87ea0948d730343b42129f;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia7ca7400e36ea572fba8e19bcc81ecbd;
reg         [MAX_SUM_WDTH_LONG-1:0]         I302e61b49accf5db556b87517f2341f5;
reg         [ 0:0]                   Ie4e5f3d7c5d2df30653f5666d14567bf;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibe2af096ad2db26e54d8b4b3bb05175c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5d9af1abff6efe3a55c6568d936b6ec7;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8cde0aa611c476b5112edeb8f17f15bf;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icaa40ec40d6d26cdf70bb5ae7d492e47;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8346f15d822cacfeecbe5d75412cb53f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5ee364aab320ab40c0f65feda6f53b18;
reg         [ 0:0]                   Ifd9345cf219c58291c0b437aac093d78;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie48569c467fba0c1291f71d6080ebedc;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1f0ecba054900f96cd7100741191c5f4;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4faf2caf62966416118a54015908c889;
reg         [MAX_SUM_WDTH_LONG-1:0]         Idd0329980a36f87859150530ab44b52d;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie66bc10dde27f08813d4d347fd7cf6ce;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie1d8b3ea7c6603cebf2f9adb776910b7;
reg         [ 0:0]                   I4f2d7bb48918ce51efe6b3b12f9f8e65;
reg         [MAX_SUM_WDTH_LONG-1:0]         I90e7ded06617b49cdb8b5301fe9c6a20;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia37488e9a50cf5cc08de74ade676db96;
reg         [MAX_SUM_WDTH_LONG-1:0]         I08aa45211cab01d567cd5eb172fd2f0c;
reg         [MAX_SUM_WDTH_LONG-1:0]         If4ff0c63ec1deb46412858e496451a01;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ife7bfd15fc4c392b5d2288d9a4e879b3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I24ac26debafd03c7333d174e8725afd6;
reg         [ 0:0]                   Ifa612e6208151c616c3a0319182a96f1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4920014f5d017f4e840dc3b88526955f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I99d80ad68e2563d0f78a0e3bb82c5328;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9943733ef305983c629565c881054bbf;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7cb4420bc55c03a6500f5228d31fe43c;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic4d19dec464359c0a9fa75148fe90c73;
reg         [MAX_SUM_WDTH_LONG-1:0]         I44993416e1d22613dbd78402c37a934d;
reg         [ 0:0]                   I9cb28a0cc6358610854c8f8d1dd3c707;
reg         [MAX_SUM_WDTH_LONG-1:0]         I03b70553f1c501609400574ae7cd73f5;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibc9b94a9dea471805cb442ac6904bc97;
reg         [MAX_SUM_WDTH_LONG-1:0]         I917d9f9b144d3bffafc77bddae7fba6b;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibc91c6c3d56bb8a14e22909c43ffec51;
reg         [MAX_SUM_WDTH_LONG-1:0]         If7c2d3eddd96b47b6c2aea8b27c8c7f4;
reg         [ 0:0]                   I40bcc924f5cf1f7d587aa35267022261;
reg         [MAX_SUM_WDTH_LONG-1:0]         I63c9bf68b43ed66c51b0f4c0ed92e9ab;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4df093ed94d26b058e97db550e347e3c;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie90303b0326bee4ab203a8cf1e643da9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I19030d352fd059156ee42c66f9270beb;
reg         [MAX_SUM_WDTH_LONG-1:0]         I36767a902c53a384128ae1443cf88963;
reg         [ 0:0]                   I5238f7273b05b8b9f376314acdc6cc42;
reg         [MAX_SUM_WDTH_LONG-1:0]         If408dfead07757878cc878131bc7d6a3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I868dffa3f07407f7996bb5bc596939b7;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7d928be164d0dce8b1322ff230c053e9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I98be4971a8a9a08abb3ebe474d7f0c6d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I779e70dea33201e9237f29681ffd5e27;
reg         [ 0:0]                   I7137f56eeb4c4ae08bbc238db4cd3441;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia0857d63d309807789b6ff4f6028f1b3;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie2262914042172ab7e08599278f36af5;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4001323da8f7956cdd480ac2d56df929;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib1cd6731034887a0a55e405c9db3e8de;
reg         [MAX_SUM_WDTH_LONG-1:0]         I51aa496e8c03944c28a908102514e6f8;
reg         [ 0:0]                   I02335be013799e2560a98b6a82a0c528;
reg         [MAX_SUM_WDTH_LONG-1:0]         I53921b825c5e434b63bee0e1ecb7a517;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6415f3996318472532e161510ccc8ca3;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia11b671b59240988737979328c472812;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id4fabe0165a117a402dc14f2f3ec626a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I57238f501ab7278b308d76211ced8cf7;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9b257f8556ca4e5402637f01081b78e1;
reg         [ 0:0]                   Id327bb65156c8307901dfcb4184bb65f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5e68f84e123c37f19a03c13892c77e19;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2e093412a9fa3972cea01664389d8c27;
reg         [MAX_SUM_WDTH_LONG-1:0]         I17907fd8c6975c8c642535ff929221a6;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3c6577b04ad56d864bbaa2c048323c11;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6f0c341c05eaa8f35bbce4521f6e8f94;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib72ba950ecf9ae2668374f6633a67ca7;
reg         [ 0:0]                   I56331cb7b310613016958553732cdf40;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id5270b57c6fb4b18db3bbd0a523e467e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3d7c72d725f4563bb562e2992093cb02;
reg         [MAX_SUM_WDTH_LONG-1:0]         I813c881ac61a59041be3be78f6a466c8;
reg         [MAX_SUM_WDTH_LONG-1:0]         I866510e7dc721fa5aac312bc5ab5ba0a;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib4432359f97849dff6ad3e0f044157bd;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic86aa6eb1b4dcc2520309089b43292e6;
reg         [ 0:0]                   Ie3b00960f8af88a5aba7a2104dfca9a7;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3c18a84617eb21472d53e598700d7f4c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0731115afe5c15bcf131f7ef4f05802b;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib080b8fd34385aa7986dace4afd95267;
reg         [MAX_SUM_WDTH_LONG-1:0]         I134890b77451d0b78afc7402a6a28048;
reg         [MAX_SUM_WDTH_LONG-1:0]         I956da75f13433c1dd7a3cbd3b78922c1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I440b26c9f1b9ccf70f97c9d5f732d38e;
reg         [ 0:0]                   I7d1ef47f35b7a4c3ea2e4383732de398;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id36663e7a01fff3170833ecfecac1321;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5e3a441faca44bffc4368d96d8fb0bfd;
reg         [MAX_SUM_WDTH_LONG-1:0]         I21d7ba25247a87a1a9c245d0d1f553b0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I55aafa8162cfc4fccfae68cf78cd1c2b;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib99c25f0d8d6493cac4d5c816884c704;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iee7c9f0a0e8ca127efee008b4874edbd;
reg         [ 0:0]                   Ibb013f036fc42687a04bdcbe2d0bbd8a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8d3be15109c7007a79fecaac0d891626;
reg         [MAX_SUM_WDTH_LONG-1:0]         I17b4a3baae65161387f472037ffc6fc4;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie7b7b202a968fe73f6b1e02a044414c5;
reg         [MAX_SUM_WDTH_LONG-1:0]         I479ab5c0e483c36267d8248340006666;
reg         [MAX_SUM_WDTH_LONG-1:0]         I777bfe165e25d7fde4fc950f23db7b84;
reg         [MAX_SUM_WDTH_LONG-1:0]         I146d505a34ddb8d65e0a1769f623a7fd;
reg         [ 0:0]                   I77eae49d321f1d1e39dd7c75829aaedc;
reg         [MAX_SUM_WDTH_LONG-1:0]         I92169cc57291f20d336a479e392ec271;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia85239bddc04bf50bcf037ed2f76d7ac;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia7306bacf3c2b180d3261a5c1f0f4a30;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2018147b86e47af5842c4f29d047d157;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id17a85459845f8a8be694c4bf1fc29c9;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic012b15584d9d25af38f83d0526503da;
reg         [ 0:0]                   I420a4d69a077dc1996ddb4b715d63e15;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6178b220b469b40dac39168057023a1c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7f09bd4a45143a036ce04af11b9927f9;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ica32f94af6e6f3eaf2b724a2173fa463;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib750bb83ddfbbad2a2be8d1c8392b4ff;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3906ece39480f96020717c6243e8ba4c;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie68ce21ade07fa53c30ebf27216b03f9;
reg         [ 0:0]                   I652202a4dc8f102d29334b4811f5628d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I55342938216a0ea0889f96c2f6c05ce5;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6cc6fa167c0d2b4b62ddbeecea175ed2;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibddf3468ae7c27d5a4b1388e524aa9c2;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iadcb2b3acaac2e1bb505c65d3cbe4235;
reg         [MAX_SUM_WDTH_LONG-1:0]         I37cd96b8b0a4939d9a70098fd8bcf452;
reg         [ 0:0]                   I0e33e0cdf39fc4cc99f6696e9f2784de;
reg         [MAX_SUM_WDTH_LONG-1:0]         Idf28431c76a84a48dd895979d2b11a63;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib34b169dcc76daee2d1aa2b2a7513af3;
reg         [MAX_SUM_WDTH_LONG-1:0]         If36fc316d6ec7c7e09eae77807b37099;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifd214c332218ac5c0fe5aded4b952711;
reg         [MAX_SUM_WDTH_LONG-1:0]         Idcd0fc8f86e2b6f03606b818b8346e5a;
reg         [ 0:0]                   Ib9479328689dec62f900946e56ba0eb4;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1ef61124c8d62e8f6a82a729fb091694;
reg         [MAX_SUM_WDTH_LONG-1:0]         If486aa8ac2cfb46f936714812cc760df;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2d8e5b5fdbda7d599423c38aaace6658;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6d0878fb7ec75c0a26be4dbba62f80dc;
reg         [MAX_SUM_WDTH_LONG-1:0]         I16a16ff0e8a6685a09803634da429fd2;
reg         [ 0:0]                   I2728682c0f749d1a9e8afeacdf44bfb7;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib8bb96f0372323e6a8072ca56fb9396d;
reg         [MAX_SUM_WDTH_LONG-1:0]         Idb211abaa54ac26e7379c64a63f7d07c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I351205eb71acb31b59d2b4470f0ba28c;
reg         [MAX_SUM_WDTH_LONG-1:0]         If5660c495bf7690252783d888d1ad6e8;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3a5229cb8e44a15560b5c7bef96e65cc;
reg         [ 0:0]                   I07da3bb5f943db6271fe1867a358df35;
reg         [MAX_SUM_WDTH_LONG-1:0]         I432f74dda4f6b1cebdf5ad59c659080b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I889b9b0828e97fe44d8366c5ef71a8f2;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie23062e00e39ead706f5b6ead233747d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8a2589544c75ecfdc31d28912c639695;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5c21c59147e9c3a74c7cbbb6f2a23919;
reg         [MAX_SUM_WDTH_LONG-1:0]         Idacd78e24408e432abbbfb0c447fdde5;
reg         [ 0:0]                   I61fc44808c85a75909b9d9fd4035f147;
reg         [MAX_SUM_WDTH_LONG-1:0]         Idc689442305acd00f0f32416d8fb3773;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0e8b171fe5080485a7f4fef83f1f1528;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib22c2bd76e6c29cc2f1440885bf24b7b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I149559fccd9def4ec1ead1fdcff3c7fd;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icfa8fed3239748abca27a5fc17de79c0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2ff115fa483f080d93bada49a9566b33;
reg         [ 0:0]                   Ic5075ee0ad355c20dd45ed594f2a8c3f;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ida03738adc101c03c2229756bed2469d;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibee4f3cd2f516c29ab68e07a640ab65e;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie495ab560f59ad038992c573de7d2f5b;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibd812def78c3a9c02f9ba45cc0413711;
reg         [MAX_SUM_WDTH_LONG-1:0]         I98166634dc80201b0cefb01d9559c228;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic2f03a980b5f0b042853ca746abab22b;
reg         [ 0:0]                   Ic0a651f45a502ead495cf14f97d65bfc;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4d14c75f28f3e516c259ea288996131b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2807a88097d2683ebdb9e0e785e3af02;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8bebbb3a676c8506af0768516abcd740;
reg         [MAX_SUM_WDTH_LONG-1:0]         I31d380f34691c9fe9022035f233b77e2;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1ffb5675c98ab5b3c62b24eb23441473;
reg         [MAX_SUM_WDTH_LONG-1:0]         If56424546ec4f3445853538207ea864e;
reg         [ 0:0]                   Ic1c05ea22f708f620f626cc8c5ca309c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6e6cbbf430d57f347a0d70558af143d8;
reg         [MAX_SUM_WDTH_LONG-1:0]         I31a49be4a34d9bac2e0d815097439772;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6b96a2498078953e87de223aa2236d50;
reg         [MAX_SUM_WDTH_LONG-1:0]         I79bf36e298a85a42c7432f877055f0b4;
reg         [MAX_SUM_WDTH_LONG-1:0]         I90c070b9bde5da05e8a5d25d2de3ba6b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I28d0e4e6d772dd58d845d91952ada300;
reg         [ 0:0]                   I61a18378aadae4556da501ce997321b4;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib7487df45118e44acec6b9d07bbd5969;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7232b4e277acc6f1acefcb606ca24508;
reg         [MAX_SUM_WDTH_LONG-1:0]         I32da124c433c55f692ffa4734d0dc8fc;
reg         [MAX_SUM_WDTH_LONG-1:0]         I56e487db14eeb8d93f494d2f11b57a49;
reg         [MAX_SUM_WDTH_LONG-1:0]         I94d3c02bd5b8e84926d4b3c2f56efeac;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0c35b2e9176f9a06e26ca67d036411b4;
reg         [ 0:0]                   Ib1fc521709a1ce2198fd8df5b41d0177;
reg         [MAX_SUM_WDTH_LONG-1:0]         I492f382fea500462b3d0866240fb91b2;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia6ee7b70d0b7fe7c346760b1784e50b9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7ce57c278c683ad045526e49bcc47412;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie3d3e681cac0bb919946ac27057409e2;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8ea0a8cdd6506c982ad75f23136bcebe;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic812f8bc775c5ee6a83e2b9aeb22b2a4;
reg         [ 0:0]                   I1bb5511c9cda1a595c45ecde48e9ebc7;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3fb3ebddaf28efb56092d19a1b4695de;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0f0adf7fe957b9a68772bd8a1bc163d4;
reg         [MAX_SUM_WDTH_LONG-1:0]         If09562f8d82bc1dea7c38ed51523a889;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib0fd21d66cd89c4e5c95fbc9c7680b62;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5a2b2bfadc638fe3fdc31136a8f09a8d;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ica914d8c556285d6b90b35747065a6e5;
reg         [ 0:0]                   I4a29c37ed36b6e12f1f8e263c92bdbc1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I22a26b7f0b1c8c16b00597732ce2ab23;
reg         [MAX_SUM_WDTH_LONG-1:0]         I00c5d739bccb0ab6d05da70fe51aafea;
reg         [MAX_SUM_WDTH_LONG-1:0]         I18e448761bc014ce490b766183350312;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1b5920f488e9469bd416a6af3072a30b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I70b41ffed4b6d88ddff219c567b8e968;
reg         [ 0:0]                   I4bf02a07719402890405fb2e7b679ed9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2ac08a2d8c917ecb37fbaf5325cb0473;
reg         [MAX_SUM_WDTH_LONG-1:0]         I935e083b4561da7d015e98ca7f02854e;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iaca9ef263bf220d786242b88c994fd21;
reg         [MAX_SUM_WDTH_LONG-1:0]         I92169291959eb33452b79bfd32618cbc;
reg         [MAX_SUM_WDTH_LONG-1:0]         I126dabc3ebb9c4157adf62b57f217bd0;
reg         [ 0:0]                   I75bd82990cb60b6d7ccd7aa2982da7aa;
reg         [MAX_SUM_WDTH_LONG-1:0]         I50ff8f51e75fb9ce3db983c2a0f57196;
reg         [MAX_SUM_WDTH_LONG-1:0]         If4433b1ef2eb963cd301946958b69884;
reg         [MAX_SUM_WDTH_LONG-1:0]         I67ac5b9b794787b3c4738c3366689871;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4f022d70078c412bdbef158f750d3da3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6be6165385f6a77aeedb88f2baaa9cab;
reg         [ 0:0]                   Ia6d3e38249f8a1208540b68f54c46769;
reg         [MAX_SUM_WDTH_LONG-1:0]         I444bc340ffb7ef7b72d4d2e761d58872;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id1f7fe91547e158e1d39edffb1421ff3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7a51924134902612db53941390891245;
reg         [MAX_SUM_WDTH_LONG-1:0]         I45128b9e29dd2fdd94a78fc5ffdff2b1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7f1082408c8ebb5be18e8f71ff9510e5;
reg         [ 0:0]                   Idf548b72357ab28fd956791e84e5d65c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I039c6cac5830759529595a958b7f65c9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I655ebf19c2f4b3dde716668f9ce12e59;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibc9d493a507122d92af42d858cdc4c61;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib3d3103e5ee4feb160a97c7e26f7102b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6cc56b119e72175df3b7ce64dc3d9305;
reg         [ 0:0]                   I50b6f2e0ef2831535ac8c18cd7ca9379;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0584de7d919236ab138e288a27d08ff1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I57cf4a9378f1cdd94a1a5608dc57e05f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4160ab1aa18e8151c0a5c23b9edeb907;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia1f183f2d904d006e46399424e06c614;
reg         [MAX_SUM_WDTH_LONG-1:0]         If979702738671323995e56108bc9376c;
reg         [ 0:0]                   I4003a2515229ca8eb6fefa2bef289ca6;
reg         [MAX_SUM_WDTH_LONG-1:0]         I086402c82ec67ae09a9e6360c58904b4;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibc96fe0a6bf1f95036f97c7d44fab575;
reg         [MAX_SUM_WDTH_LONG-1:0]         I755a38220a693ba43701d30e7e9508ad;
reg         [MAX_SUM_WDTH_LONG-1:0]         I896fb82baa9647a14f4b5b1ecfa70a15;
reg         [MAX_SUM_WDTH_LONG-1:0]         I23d1c973d7a2048353fbb68e4a294c08;
reg         [ 0:0]                   I48672f8b83eef8c406694676746469e7;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1cefdc831c146187c77f861b3e2d1af0;
reg         [MAX_SUM_WDTH_LONG-1:0]         If9fd1e08af14f2fd4ca363383f48580a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8f3782f78d88a5c3bc93709564999b30;
reg         [MAX_SUM_WDTH_LONG-1:0]         I986d61d79ce31f4677f3293339db6ad2;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ica4d93d9fad21316002008ade5106a9d;
reg         [ 0:0]                   Ia14a60c9497c0faf3f1f448ff2abe553;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ida9c16ae57d17b6faee8a54838860447;
reg         [MAX_SUM_WDTH_LONG-1:0]         If77592d5d8bed32477fd690341e543d0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I25b70c6b830cbfe1b41d8f289c751924;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2a5d65eeffa18dd9af9fe36463dafd7c;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibafa6e10bd4edf5d224fdeb2f9adbf98;
reg         [ 0:0]                   I0ef3962dd323e8ec64c4a881bd4b3044;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia3b9fb112f39dd0ccbf7555659369efb;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifc25402bd879bc5c43b4945b60cd4540;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iec48da6882325d8a33e0e0e845eb18a0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0fd05e46862fdf8e614afaa3fd478602;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6253a59dca81842d9ab6e58cf204abbf;
reg         [ 0:0]                   Ie9b64c34e31dab63c03b3de4528d53fe;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib1bfcdc0c972aafc99116ed8c0511445;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib18d64bc58b354358ee6ac16785880e2;
reg         [MAX_SUM_WDTH_LONG-1:0]         I28689b693a7a5f761a1f252aa3ef3b67;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1a4e6d12f9776d5e61094e0b5edf71d9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8e1ad23b7ac662bb827a83d3709f0adb;
reg         [ 0:0]                   I5941476ded9f6dc25d7394f5d133955b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7adff505c50450a04f1717cac1adebe7;
reg         [MAX_SUM_WDTH_LONG-1:0]         I000ad2287813072cc18dad933758f2ab;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7bc3698b51b89ac38ba5f4b5428a0c96;
reg         [MAX_SUM_WDTH_LONG-1:0]         I78aea1705621e2845a331c3e61a8055b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0a31314c3580f5f9e61e79c133e5d794;
reg         [ 0:0]                   Ib46c78ff661ee6fb69c704d39235ffe1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I699feb4382974a02b21cb387c13f7f3f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0e274fd7bfc0388fef95a8ceb939ee91;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id6f39ddcb73d3f4ec081a365d11d1ef4;
reg         [MAX_SUM_WDTH_LONG-1:0]         I807770bfa86d160459d6ec3c0f4d6a0b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I31c89b8a11a3090bfd74b112cbc474bb;
reg         [ 0:0]                   Iadabc5abc7dfbc1dd747179ad7e37850;
reg         [MAX_SUM_WDTH_LONG-1:0]         Idc99c3b23e49aca3c98f0685ea34441c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I79b82cb1bfc72bd5a9d313b9e9c9203c;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib1046ae03c9a77fd2c0b3e9838e9af87;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic63723fd43cbbbde51c233a3cca15d3f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3abbb59abada1aec6941185f95f738bd;
reg         [ 0:0]                   I97a6b5f0976feceee3a5b5890d4d76a0;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib67318fa6954ec8f3247927d34e74f8c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8d5bd7039a77ce82ce0f6cbba9c2a076;
reg         [MAX_SUM_WDTH_LONG-1:0]         I527ad0b9382dd7b6e657dc1a32d8e472;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8de02f32e14e719f4930d99743c04a20;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7614dd5e9628c761dd9b2a512cb1da98;
reg         [ 0:0]                   I7217d4790fec9797a1eb8cab1ebce71b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8774ce3f11362915c4331d1026e452dd;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icae7efa4742dd0ad943ee1f67b0c9b14;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ieb1854b79e9a2bc6cf5aa1c319e8e753;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iff50b77f300183ca59a67ccbcc9573c4;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4868604f8178663de759d4c63dc6c4bd;
reg         [ 0:0]                   I3dd024db4130c105a6817e8a4935de0d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2392b2d17ffed6073875fbe8e92534cf;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ife992a151986c58df4cba79b6bc4ac0a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9ab973fb74d9fac5d78eb8fc2c7ecf36;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5ee7916e859b86a98538659401685016;
reg         [ 0:0]                   Iae502e5a5ae518fb7b817afff28b7932;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3a4f0d3e32596ef05477f494768d4266;
reg         [MAX_SUM_WDTH_LONG-1:0]         I48c284cefb8cfb5a938a8f23ce4d7f03;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5c1fc666b77a689478654dd29519f458;
reg         [MAX_SUM_WDTH_LONG-1:0]         I38bba98b59184c75ba3b27e1dcf52182;
reg         [ 0:0]                   Ib8b2b1d90204af5b100379ecad20fc0f;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icd08ff59cf6be3ba97698dd55703339e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6905b65403c16b0211643227ece536f6;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3ed34401bba9d5f229bc98480aedd9a5;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib4d05804277cddc7f00ac17ac14f5325;
reg         [ 0:0]                   Idf0e651d0b13e167df3c0cc40d149c29;
reg         [MAX_SUM_WDTH_LONG-1:0]         I985fb7ed22a8476ea322c9e3c2b3851c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I41babdca6d3fa462849592d37b0a7998;
reg         [MAX_SUM_WDTH_LONG-1:0]         I58cfec706dc929ebfdeaca6e01b00c0a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7efe3c5b2fc69840a79545e0399ce749;
reg         [ 0:0]                   I89daaca029498d05ca62c095db439eb5;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib985709316b1b0a9d3fa3c1eaf6c641f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I70e3eeb2b3966676d16a6aa4c85753ab;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2a32d545d1e7beecc7531174c7e8dfbc;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib8fb40e4ba0ba1f5e9f5a99d1271ed06;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ica792cb9850a61fa4a8bd8a4b6c6ca05;
reg         [ 0:0]                   I0fe5a34ceda936d0924efdd07fad11e5;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4be898887dff6e2cebe53f135ece131b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I779e5997c66649d6d54fd7f0514c47bd;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5aa578b0c2831453683fa44af1878cb8;
reg         [MAX_SUM_WDTH_LONG-1:0]         I735d6229ef1a4ecda0a1f1dbdfb53fc1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I62affd47512c5e8f0979244115624d97;
reg         [ 0:0]                   I7876cbb2b5d8aba3652ec8b218080dff;
reg         [MAX_SUM_WDTH_LONG-1:0]         I004db04f61fb57aba81e15cc015442b3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I14fe27afb3df5531b18dc9604e8dbe65;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib1b1626c84dad8ad13c058f921ffd57d;
reg         [MAX_SUM_WDTH_LONG-1:0]         Idf4a4bdddb88c21c5afe10a02373a6eb;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iadefc2a3d07ed4b2c3c46b2ab5dec252;
reg         [ 0:0]                   If692ff56ce90d22d7af881599c54df75;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8f7e3dfb2f728d4cd1e79b82b62b0406;
reg         [MAX_SUM_WDTH_LONG-1:0]         I19315957077b037ffc6415dbb06ef789;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1f9be09334407fc86c83a7c127e17bbe;
reg         [MAX_SUM_WDTH_LONG-1:0]         I28e17a5af7a7286a2643100d6d058dc0;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icb2297c397bfe56be251ffb6b249a020;
reg         [ 0:0]                   I18a7a4fe8931c79df3a69223af46c440;
reg         [MAX_SUM_WDTH_LONG-1:0]         I991054370345e61638ddaf81785505bd;
reg         [MAX_SUM_WDTH_LONG-1:0]         I64a48984527d660002f1f82c376c7a84;
reg         [MAX_SUM_WDTH_LONG-1:0]         I238b5fc70ce9f05b6322a2691b3a0207;
reg         [MAX_SUM_WDTH_LONG-1:0]         I00c16e7ad3821981032a42d5baa767b3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I42fd5b094da200b33036e6cb8c7d0286;
reg         [ 0:0]                   I8eec3538b8cc9c046954b6804cc656b0;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifa1f503965270d10e7a5c9a15576069b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I98b7e26a0e9ec9ad750ff87cc0641a73;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3ec904916870171bf837e162d1030052;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iedb11b97900b7dd769d31f8a89521975;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id0dceec6497c9f13ada07138986d4145;
reg         [ 0:0]                   I653767e659590c1676edf6c25fc0e253;
reg         [MAX_SUM_WDTH_LONG-1:0]         I24f773842a4742fb58d09cae45717b2f;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibfe7d9bac29b8838f20cdcfe8ef7da0c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4d6c95605595942a34573d6ed55eb326;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id6d8f32958dfa1a98958a84e7f1aed02;
reg         [MAX_SUM_WDTH_LONG-1:0]         I971cdf9ddd1bfff5664eec35f22da335;
reg         [ 0:0]                   I5ff863be142b92dff89f7916d0d088c1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5bac7e0d778a547a0ae764fe259b6f7a;
reg         [MAX_SUM_WDTH_LONG-1:0]         Idd8bc1412a0dc5f489ef253a6164ceea;
reg         [MAX_SUM_WDTH_LONG-1:0]         Idbeec36de0128e5924e214877c82bf11;
reg         [MAX_SUM_WDTH_LONG-1:0]         I50a9cd240979bc56421bf85011ae99ed;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6437095f6bad2d4fb2fbe0361f60bba1;
reg         [ 0:0]                   I49f9fd0e0719be527f2a54814dab83ea;
reg         [MAX_SUM_WDTH_LONG-1:0]         I255577ebee6768871df0224fc1db2db3;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie9b6eb3bbac26635aa00c38110958d46;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9f34e81e3ffb85539a6273babc2a732e;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id0a1ab8472d704001e0eba0317b117d6;
reg         [ 0:0]                   I945f2476eb599844cbee0cd89038e392;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia7fb4af3d3529a32f902a52cf5598474;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9e632217cd0561d8faa28e4b8850d995;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iedeb5b7b2fa8acf1ea083102678710ea;
reg         [MAX_SUM_WDTH_LONG-1:0]         I972431d1f5af0bdf4828e4f85591e358;
reg         [ 0:0]                   Ied0c5f8a9243cd9d93672ad6cc907d21;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2c98806141f064c9e92935b23a84ede1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1f41024b715d8312944ccbf70e95bb40;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia6bb5ca05f5d0af452c994dd50004e1d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9a1d1d1c862808f9a769cbdb3bc634e1;
reg         [ 0:0]                   I9134c7f579723c7615af60b4344efe76;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5680847bc8d224fa4ed93b2fc0d841e1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9734eb86f4e73ba217739baf5cb1b13c;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifc0fe00f86569956df72d8a960337e8c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I223341a807a1d555f759632f67815159;
reg         [ 0:0]                   Ie92388a9d1e71d73c07ed86e9bf6c887;
reg         [MAX_SUM_WDTH_LONG-1:0]         I365254279ebb10dd7ba0b3482d5e34cd;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6c1f5cdf5f2917118941f4af14d67fef;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie84e88fd1aa2a0b90aa1715fcd27a329;
reg         [MAX_SUM_WDTH_LONG-1:0]         I558f70d7039a8bb58d8ea3f72e43dac0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9924269ed3de12f1f2a28893c7f95292;
reg         [MAX_SUM_WDTH_LONG-1:0]         If1153befd1396be2798cc14535ddeb8a;
reg         [ 0:0]                   I6804fecdf59233c6cf14409bf2f1e430;
reg         [MAX_SUM_WDTH_LONG-1:0]         I57bf4ad773cc058ae1bb7b1911dc3174;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9bc447b20687fb3e7eff45792bd4dc3a;
reg         [MAX_SUM_WDTH_LONG-1:0]         If590520f01e452db9867a8d6d5dab29b;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id93ee7d283016ab9b0aaa21237237c54;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic1cf03baabaed466fe532e4db3a9ea78;
reg         [MAX_SUM_WDTH_LONG-1:0]         If3031f9aa8f6eba90eac12db7839fefd;
reg         [ 0:0]                   I9e777a342bf53eaba0280737ae404bc1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I57072dfb29c4a3d2e2b40e46e62f0d95;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0dc2708970ca2b6c092273b6626bacd6;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia58944aebf0b4f0a7d76a1444fced9de;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iedd8e69679d10e05f2889f1d71cf0e7b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I90f0d471914a2333b9dc14d6d01cf927;
reg         [MAX_SUM_WDTH_LONG-1:0]         Idceeb22013af64b6bb9f0d773e9ffe9a;
reg         [ 0:0]                   Ied53820aab06b5c3423b1d878c71948f;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id8cafb6f76321bdaba9711133be7be99;
reg         [MAX_SUM_WDTH_LONG-1:0]         If43574342e60a625fb6bee5a495e88f3;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id285f055275014d9f23d35f91879afa1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8c803ab08db372802117de4fa4e2a187;
reg         [MAX_SUM_WDTH_LONG-1:0]         I13ba48a6b360f3cff5f37ce60cb735c6;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4547cd1dad45dfd01e335e8cf20eadd6;
reg         [ 0:0]                   I24cceded372d782c67b33f3a78b16045;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6344e71ca2b0fd39d36caedd889c3085;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0a305655b815b0cc159ac1c5f4ce30f8;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3633737da6b74284b0ea9a06c3f5875f;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia949c1b338d1cba07cf6bb6572c3e322;
reg         [ 0:0]                   I2e78d36bca5bfb016af674c343f9c041;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0c99a68e0bed90afce18807acf7d55bb;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9a0185f8400159415bc0ad6c38284041;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3eeffe43e7deed7ee77a7f5a3bce3cd2;
reg         [MAX_SUM_WDTH_LONG-1:0]         I85af0c31ca7002ae569d9f5ce39943f7;
reg         [ 0:0]                   I17a9a995de58643dbbfb78604f26198b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1c95650979c86310ae2a949961c9db11;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3dfb8d2fad83fbd807fbfc6330c5b857;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic12be21bcba5fa49437cc44dd8a7f064;
reg         [MAX_SUM_WDTH_LONG-1:0]         I713a384d022d3012e3d0019f5c4ac077;
reg         [ 0:0]                   Iad642c4c62766e8f8bd5a1e9e73bdc80;
reg         [MAX_SUM_WDTH_LONG-1:0]         I04eaefa5d133e53494fc270b07be7043;
reg         [MAX_SUM_WDTH_LONG-1:0]         I80550019479d0323d0dd7e7d0f767d83;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib8a866f080dd997e0b6c93b6c844d1bc;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id542de206d736ee3769ea0bd037cb627;
reg         [ 0:0]                   I96f92481be1ac6cf985b8ab387d326bf;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4a64fa2412eb8058c2dfd9351d7b297d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I77e6cdb09c92492c3303d0213de9c291;
reg         [MAX_SUM_WDTH_LONG-1:0]         I788c33a9f94b26f4ce0f515891d06f90;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iaf7074c2b570a296fe2ea8a5a7097ca0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8964c6d3f8e02866a6ad86553ab05d99;
reg         [ 0:0]                   Ie03c09039ccafb427153d2347c1caea8;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie8bb2fcb752c6a33254963d1ebb4130d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2aa25edaca90c9dae8ed63b48d333c17;
reg         [MAX_SUM_WDTH_LONG-1:0]         I51a440917c7ae23339bec6f8a745c103;
reg         [MAX_SUM_WDTH_LONG-1:0]         I56ce875e4619d4d8d6ca2fa0ddee91b1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I80607da8f92f5a5d2e4798a62a7b1c5c;
reg         [ 0:0]                   Ie7381a8294b4cdf669b9c57cfe4012b5;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iac05b7e3ae18f948b72c356ccfb8000f;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic4dcaa520e26bac40b3876f02074f856;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3b2714d34081a3b6cccc47fa1638e72e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2db1d1ee8f546c00e512875ce2e13cee;
reg         [MAX_SUM_WDTH_LONG-1:0]         If80a6bb104ff3b2020e909103c104063;
reg         [ 0:0]                   I61c9e3f8e42f869f4c9c1386325100b3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I27da3f75cca6c49e55db90306aa68e94;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iadb72cc5444816fbd132256493930bb4;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3a8ec1ad07bfada3d2c6ffca88b8b678;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0aa042b86d9f68d22a49b4eb480a9088;
reg         [MAX_SUM_WDTH_LONG-1:0]         I89a387374771b68d87d7ff2dcc810829;
reg         [ 0:0]                   I24c5b2de59eb1f43fe1efe687231c4b7;
reg         [MAX_SUM_WDTH_LONG-1:0]         Idc7fed723190098341225fe01ba65ced;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2935b3d5c3bba4dddfc7ae03fa77b229;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4e0c0248f4aa97d263d64dfec36e3aa2;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia2871d7493b2727d2cb2fbab596b7e6a;
reg         [ 0:0]                   I43d43acde5f831fc32b7bf5f10b9b3a9;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ife9065805598960919ee4f14c3cc6fd4;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie57adae8873946d6c706074b52a49786;
reg         [MAX_SUM_WDTH_LONG-1:0]         If5ac85646e4b339a19af658f01d0a17f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1c092426f34be030b3e020f40517b0e1;
reg         [ 0:0]                   Ib06e93161fc8ca3be232f4261b04feb1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I717c5c2d6a2be61593492ae5f17a112f;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic719b72ad271bc7c077067518e6bbb98;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib87362230682c88d68a0ba70e25f3c20;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifcf097a102f8dc1f912022fed893d222;
reg         [ 0:0]                   Ia0dd00f83afc805036f2c6a0e38f725e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4c31fa8e6eb648439cdae1de1afe0d6f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I56483ca3fa550dc59bfa347780cfef7b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4aa9f61be376458185c3235442c8fda0;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id91fde1007d47258273299de80721390;
reg         [ 0:0]                   Ib0a0f924fe3757a1e0aade7017ad9277;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iead549a9af27f1fced7d9c36e7b5c3f5;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id58498c34aff2e1216c189b9df88822c;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib52e0c68caadcf4dd9636a84f5460e53;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie19679053b289bb5a0aad570cc81bd14;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8862c5ef45b723c9abf5d0ab6854a900;
reg         [MAX_SUM_WDTH_LONG-1:0]         I30db951a07af96a8ddf59360141b9a6a;
reg         [ 0:0]                   I1ca949071d734d230cdb8adda46c9d79;
reg         [MAX_SUM_WDTH_LONG-1:0]         I10422eb79364e7d0e21e1643d9060331;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4855a0a0c6426d33014ce6a4c96965ce;
reg         [MAX_SUM_WDTH_LONG-1:0]         I362e8db1791718290bd33a79b4fc0855;
reg         [MAX_SUM_WDTH_LONG-1:0]         I773f0508440fb71d73fd82a372cc0a00;
reg         [MAX_SUM_WDTH_LONG-1:0]         I792891cecae468d7a87e12f2da62a718;
reg         [MAX_SUM_WDTH_LONG-1:0]         I33303820ad094d7a0ab53bca722fc609;
reg         [ 0:0]                   I40170922c652fa7fa42abc6f580b5e3d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I914cb87eba8baa40cd515334e59f26b2;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iff98739de575e25104c0dc30f08912a5;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1952614b64ea451e9d0646dcce5dd1cd;
reg         [MAX_SUM_WDTH_LONG-1:0]         I49c1a7d1c20a25496821ad80c7eff790;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie2be17a55e79ca76350e033f227800de;
reg         [MAX_SUM_WDTH_LONG-1:0]         I737a5b06f848cacf0c8da4985c73c66b;
reg         [ 0:0]                   Ib1ad0b531ac9028971d68f533e7ae566;
reg         [MAX_SUM_WDTH_LONG-1:0]         I32ed679af4ab759901aee43c9d93eb67;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iab160609bb21501aa55b662d2010357b;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ief74f1a9d4a43ee5c9def7b83369bb21;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id144423f50751e661db3860a8487d004;
reg         [MAX_SUM_WDTH_LONG-1:0]         I623352a4f6705b21d461d6b32e85c12b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I28d1dc8dc594977b5058b5bb9f6bfc66;
reg         [ 0:0]                   I0ab0170c7ceffbb58377b65d2ad92093;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id376dfa5141402f4d41a8858180ed87e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5371a83bf9d6f334cf8d1c5b082527e9;
reg         [MAX_SUM_WDTH_LONG-1:0]         If1605d6646fd267e701668a7245b3b44;
reg         [MAX_SUM_WDTH_LONG-1:0]         Idf5eb1ac2c5bd92fa08ed935ae298255;
reg         [ 0:0]                   I9ac68f228a93bbf4aa4a559b1364e42e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I98a384bc62ee03f5ad7df20ef2d9af95;
reg         [MAX_SUM_WDTH_LONG-1:0]         I44ce30330c4d2d6033a0a970dd2bdd68;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic101b8f56ea1e25c6b752583a1b01242;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib7cf44e681881e55d2d353280a6319d6;
reg         [ 0:0]                   I375c5f7eac92d853e85e0606011f3fb0;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icfed259ca2bb2732d8e0c26ef67cd4cf;
reg         [MAX_SUM_WDTH_LONG-1:0]         I35690f724e964248dbb1e80fb1ea49f8;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5affa2759148a6baf5b9f0cd3122348c;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iaeea1f06ff0c6e9cfa43ba14420c3adc;
reg         [ 0:0]                   I94f9b1f2e63748c21ec7222c9641366a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I20861535c450d6e6bf11c45dac120454;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iac5a23266c3b038b4b54a916dccdf3a8;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icdfb7f52cc27b1cfcde90a100d29af13;
reg         [MAX_SUM_WDTH_LONG-1:0]         I71484d7e00efa02a08b54a1405f2902c;
reg         [ 0:0]                   I55500c1d85c4970932be67cc5cd2e023;
reg         [MAX_SUM_WDTH_LONG-1:0]         I013929385ad819ddfcfcc59c22902ee3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I68a9b0607e69e8b3dae64689eb288a33;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2598c48aad48072a7f216b2ab56ee532;
reg         [MAX_SUM_WDTH_LONG-1:0]         I796e3a193b1b66fa9a04ca60aee11ea1;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic96be7e69faf0f43b92618131cf0c98a;
reg         [ 0:0]                   I36b487cd1a57a3a503e587fdefbb19e4;
reg         [MAX_SUM_WDTH_LONG-1:0]         I34fffcb07fe82f11fe142f7c37f39155;
reg         [MAX_SUM_WDTH_LONG-1:0]         I648afe4114ce435bf1d13e0ad54425cf;
reg         [MAX_SUM_WDTH_LONG-1:0]         If05d7e30b4717e0a1bfd20b90d0539bd;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5fc356af8a62a1d739cb375fb851e90f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I22f4c5403fbe33d18f97cf21786cdd80;
reg         [ 0:0]                   Icb5350e8c55a2adb370078a7575e28f8;
reg         [MAX_SUM_WDTH_LONG-1:0]         I61ca60fde05ed88cce714dcd8c13b827;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9a1b2b9f924099f1e57fa501ba2e33ba;
reg         [MAX_SUM_WDTH_LONG-1:0]         If6253af4ebc430e4937269a5f4989b29;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0427d17423548dbb33cf792883b4be8c;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie539faf01ae85253e399308fef98afd6;
reg         [ 0:0]                   I8a7a31327c9e4cbd88ce39fea8971caf;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4907dd45c158dc7e0041c64f1fb388f6;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iae6e7c42f250cd9223f18f8830fb177d;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iff47ec1743b59d7f90e9042af7ce44cb;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1cf4a55ebab332defa32d2922b885285;
reg         [MAX_SUM_WDTH_LONG-1:0]         I284913858691ad5724073b73a820047a;
reg         [ 0:0]                   Ied069655ed3775819d0bcb722d6d0488;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2c8f6a9b9f655b317bb0af4d60fdbc4b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I35626ca53adbbf0a3a71cc6fcf43bcb1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0d74ef22d31abcec73c7c582310b1e6d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I15f4cf1aa0ad5ce2bda52df338e677e3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6c5ca5e68c8844bb1617a2288b5bbc37;
reg         [ 0:0]                   I78a5fc80d42e8db1b56cce5f4c97e325;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic7dff631559304ec59f0696c66436d62;
reg         [MAX_SUM_WDTH_LONG-1:0]         I44343a9491069c3c8ea4fbd6255a5a6c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1d8318b94d86e1fd28323a5e5684a37b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I825e83bd88575868f4fcc9a8b8729663;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3184a16c71cff80c8c90b40e45f114b8;
reg         [ 0:0]                   I3ade7e345432319c1a9c91d4068b3ec9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6a239d3e55b4a9a3be9989a85bbec545;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iae133550f8bad8357a73e7de1372faa3;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibccb4a43c410f698e0fff68553326a77;
reg         [MAX_SUM_WDTH_LONG-1:0]         I72dc7aa294a3af89101ea62a4223170e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I91eb3e70921e0b141a344bc57dfbc934;
reg         [ 0:0]                   I88aed46f6dad7a81006562a720670654;
reg         [MAX_SUM_WDTH_LONG-1:0]         I630f905e55f08e7d1569a08e937ad216;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1986f22f2269cc135c6ed28d35fb0bd1;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibef24017bc71de9c002aafa7ce9a784c;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ieae3ed78fa2c45507066f4e20d96e956;
reg         [MAX_SUM_WDTH_LONG-1:0]         I730fd25ffc7778fd4bb02d33cb3870d6;
reg         [ 0:0]                   I79e574dc9c7e18b695c9a2619b71b995;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8d13eb3669785c4279c685763d4f3fad;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9a32313f2911b797fb0848f7d97e62b9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6373e2d64fdb5dd77733b3e4bb405121;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib437aa67ab7c13b45d7a4d56ce9e79b8;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0cb5c7a759f4c75d4a675f9777f15c5f;
reg         [ 0:0]                   I800ef583bec1d46d3d4ffdea6b312ef9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I25a6f3de9a9a01cbbdd32ed848561aa4;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0ca91c1426ba14a7b47a081cb3becd19;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0737e0cc7453e328efab2277bb712ea8;
reg         [MAX_SUM_WDTH_LONG-1:0]         I456af863661122cc303fccb235f3c7a1;
reg         [MAX_SUM_WDTH_LONG-1:0]         Idc5916c4800e9f647d51c52444ab6fff;
reg         [ 0:0]                   I56cc5cd6d0a5a4e4601fd48e838fdaf3;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iba3dd4b2c2c85c4cfe770d9b52ef4634;
reg         [MAX_SUM_WDTH_LONG-1:0]         I57aca70e2b8d126c120736b2606ed333;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic6650a6d092b749b4498c08d69cf815e;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic2e3b8f91eb218650c7b9c515c7efe97;
reg         [MAX_SUM_WDTH_LONG-1:0]         I93a084aa1e6881ab8dc905dcdcdfd7ee;
reg         [ 0:0]                   I21047a3955b8b89bdb9013d571b2bd0d;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie1b744387b5200a504e4874e14d2f282;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8cba172573be52c5a90bd40e6f40a508;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1cccfd1516af59265731121dde878116;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia171bbefe2d20b4c058126c33ef28eb8;
reg         [MAX_SUM_WDTH_LONG-1:0]         I84bc44a5d53a8f66b985b70c7ec1ae7c;
reg         [ 0:0]                   I56eb529a34b484cd20e29958cd6878eb;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icf76cb69aedf4db01cd3444f4c4ba471;
reg         [MAX_SUM_WDTH_LONG-1:0]         I321b104ca3c818018d4b03adfe1110b9;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia79b8994da536c86634bf6f54a21145d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4df55ce80eec5fee295b5a0ae92bd6c8;
reg         [MAX_SUM_WDTH_LONG-1:0]         I46593a7956590d870fe680228081a6d2;
reg         [ 0:0]                   I74588df6399af2c1112e3fa557e89e17;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4857b5b50556c8e7fff4b2d3e08e4b28;
reg         [MAX_SUM_WDTH_LONG-1:0]         I906e9da31de73ae45579607a014e8b54;
reg         [MAX_SUM_WDTH_LONG-1:0]         If5dd1a1b9e3fc0e67a85da3183480aed;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iadfb1571c78c3f0c05e4ef498267df24;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icebb43b184c2745cc9da9d01b06bc62f;
reg         [ 0:0]                   Ic8eae1a92f46db040eb22d726c3a0e6d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0a1e9cf99f1d4725327615f50fcc3ad0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6e4b0489ec7333abf2245a1b72a8923d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I24ac5dd30526c1d3bc7b941103a66804;
reg         [MAX_SUM_WDTH_LONG-1:0]         I33681b2292c086fe536dae2aec70903a;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia373ca76c3b15a4148532b3822f82ba5;
reg         [ 0:0]                   I854a15bc7e9728b01c9a1960f6248dc9;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie844f4c446983ce381b0bc4c0e8ef7d7;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7d08adbaf66cea04be4891db610bca3f;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic09ed51b20f411683a801eaad61657a3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6a9af8c9009b5de47ebe9ee8b79d3831;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ife18e8a16d4437161b75a93e3dff1b5b;
reg         [ 0:0]                   Iae332cfd000fd0529684ab787041b5dc;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6067f47cccceea96ac46ff0d457b25f2;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0cde86532c8db1a32d9fbe38a40b91b8;
reg         [MAX_SUM_WDTH_LONG-1:0]         I49c8ec4cd33e6caed8ed7dab779e7ebb;
reg         [MAX_SUM_WDTH_LONG-1:0]         Idb86f95570587a0711d796aac7004c25;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2d1373d0b18992fa46a9607a86d21520;
reg         [ 0:0]                   I70148fe95244eebf7f0ec953703398de;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifd6fd1f3cbf8884ca7f64bc42278e4fa;
reg         [MAX_SUM_WDTH_LONG-1:0]         I30f26e090ab14551cbac41883ad8a152;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib1b4e41ab25733d1d6dd54e1fe81a419;
reg         [MAX_SUM_WDTH_LONG-1:0]         I146c0d5154a6de44c0536de873904ccf;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8eb9d4839a478a4e28b45a549b5682a4;
reg         [ 0:0]                   I24ee2d953e65fefdc73b3d3c4c0ddd05;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iaec9fd9e79371676bfa8ff14b4feae52;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2501ef991a59512c43693ba9d7db8571;
reg         [MAX_SUM_WDTH_LONG-1:0]         I38213f78fd4dc52f9d2c9b7b22136c1c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I49ce91ac152279af421bbc6c4d9b8087;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6a2b7bb2cb3ca2ab932c211a68dded55;
reg         [ 0:0]                   Ie3a5f8eec283fd4f682b5d0f909b051c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I500757c4eda5d3d899aee47b87da585b;
reg         [MAX_SUM_WDTH_LONG-1:0]         Idaae6ba9da8754615a2c34ef859492db;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icaca9fc70a3ec6c48c0e41f8168e2bb9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4f69b8ff834c7ab3194bc9390ce0f5f6;
reg         [MAX_SUM_WDTH_LONG-1:0]         I037cb596cd48c5533ed22bc32518d992;
reg         [ 0:0]                   I781d986d7fd6c2fec3a8cf3f29545174;
reg         [MAX_SUM_WDTH_LONG-1:0]         I47bf091b0fa74ad511a760bad9d2506c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I94a89577951de90edc4f73b281ad7364;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib7493a1a384aebaa7999ff1fb867fc6b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2ceb9e423696539135c5bae5cc2d8d98;
reg         [ 0:0]                   Ib4db8131350f8605e00907234aff901d;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia4c3d0cd9957f678880de5775de76e0d;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia6bbf236436b2ed22bbaae3b8849de6d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I33cdaee4676d546dd5507df4704ea1f8;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia44daa9ddc3e4d377267333813d4675f;
reg         [ 0:0]                   Ie093f0750b60d3aed75705637933f34c;
reg         [MAX_SUM_WDTH_LONG-1:0]         If5f957fa2f055b1c2c28e8d7cfe3e9ad;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie1f8fff3f43426d6bc39e45322a532ca;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4ee181895efc22862b6e85802a944095;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5c24ea83cabbb6be089ac084732cb9d6;
reg         [ 0:0]                   Id2fba7c1b3dc7a75a5e0d90494d56962;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3608378a5da8c66bef58528d56192530;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifee2342449a3b3d0036ce2ecbc9ae189;
reg         [MAX_SUM_WDTH_LONG-1:0]         I70a9a9b8f25066612a50e411ad68e6c4;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1870059af857c79d444bef948bb536ef;
reg         [ 0:0]                   I9ecee74c445711a376133636ef414666;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie6dead855e00ea0a8e6a9b7503aaebb8;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iafe61ab12e232a1090123a0f16eefaca;
reg         [MAX_SUM_WDTH_LONG-1:0]         I10ca809fe9a04eaf5d7784ba69314178;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7a1bd0a115b3a1f85cb9c54840f5bf9b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I986a564393d944d7d202414431c6d165;
reg         [ 0:0]                   Ifb3cf6b88835d27220df837682c4dc93;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3bae5e6862e003a8b9a476f72cc6858b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I464042aaa60a41c7e1faf3d16eeb121d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I34b9a0bf2b6b562fb36291022ddf5179;
reg         [MAX_SUM_WDTH_LONG-1:0]         I17dd8612b5c7f9dcc90f17e584aab2d3;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id77cf7c05844d83e808a694971145261;
reg         [ 0:0]                   I386fbb3bd550891d682e137044e8773a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4431adecba8be9e5f21bc6b3e1f8cb10;
reg         [MAX_SUM_WDTH_LONG-1:0]         I276c1155d766437253f12b25066b84e4;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id75b386d8076893cb73baca69c3eff59;
reg         [MAX_SUM_WDTH_LONG-1:0]         If62ddbe87274965cfd83189c6666401e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4f73a07452638a610b31e3ee52cb5639;
reg         [ 0:0]                   I7ede7d2e1c2730b3b71340b11e880f5b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I21c7a2885126d532d00484376588a469;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2a4faf3344d9bf4ee71da0be8994788a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7d7ad0cbb962a47e229fe9d8406e6fe1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I82988dc2dc83ac61380d2a5cb6551768;
reg         [MAX_SUM_WDTH_LONG-1:0]         I058c3a9848fd30010e4742d8682081ac;
reg         [ 0:0]                   I64c65fad4a7d958d625c783626808175;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2c4d7339ff2fe68d060dd8d961dcab8c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I368121c2534820a7147858c06e58b3fc;
reg         [MAX_SUM_WDTH_LONG-1:0]         I03d4541eeb1440aa72ee490c49977e32;
reg         [MAX_SUM_WDTH_LONG-1:0]         I75fdf5a355949a87b768b1e67db674e4;
reg         [MAX_SUM_WDTH_LONG-1:0]         I088f4a0af0239602d422324549cb9799;
reg         [ 0:0]                   Ib2e0cd0a2b51c3a265bdd20834c0ed2d;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iee518b15b067eec58cccfa37f7432ea5;
reg         [MAX_SUM_WDTH_LONG-1:0]         I787fe66b38237caf805ec14970d154c7;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icef176cff3ae503dbbe2af9ecfc4c859;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie0a66e4871bfe94f6716279ecc9ef21c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I474adf7a975b405c288058139a08be38;
reg         [ 0:0]                   I67be0b66c8d0680eb23290a4b3885af3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I42145be9c2a80288ba4a2edd91f661a3;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iebeadb39658f41dcf8719ed413e46144;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie018b0d9f05a86207ae09ca2efac54e2;
reg         [MAX_SUM_WDTH_LONG-1:0]         I51ee69807609fca0f332c8bc31afd632;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iee1cb471704b2a8718a68ef93fd2e356;
reg         [ 0:0]                   I01148401f7d058614dc1ae6ed3c8bd94;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9dc297ad41fafcda77f5347f331cfc25;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1731c0e3be86eec142c3732ee836e4d5;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id3b8c0ca32331f94fd98c8dae72bb15d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6a86b0a82441c6c14436a3e0af6b0fb7;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8c92ff598084da7a50f7c68da96620b3;
reg         [ 0:0]                   I3394319c370daf6102be00d938d55769;
reg         [MAX_SUM_WDTH_LONG-1:0]         I846700c79f30ca954cc2933fc94d355b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8bd1862e7bc2e83e9863389d532e6623;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8053269f8bd78a931878c8350693e1d6;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2ff66cdd7314276232715ef2361ad184;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icf541c76bfaf37fe6111de037d205f15;
reg         [ 0:0]                   I24d6a334dd15ccdea558f32cd029e6d1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8af96a91457316e49e3f7dd5e57c82da;
reg         [MAX_SUM_WDTH_LONG-1:0]         I68319c8b9febef9f564832429c91b85a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I127772614218dd7c50d3136b4f174d7a;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib8d1aea4ad24c6ceb44f2cc672e1ff90;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9ca26c8104bf15f48b19dc3256914544;
reg         [ 0:0]                   I3a41f68bca2d7edd1f5738c4fda8e73c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7d1c247500d7d32e406b2a5f7e2b745b;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icc76d9ffc3f3d7b410205eeb8232a33b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7fc4551d8a0445f79b87b4ba5f2ffeaa;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6b3c66c4e3fa0ef0cf0b52eaa4dac7a8;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie34c07af9f6adb9e4b636dce3d0682c0;
reg         [ 0:0]                   I9ef1784d165492f3482d14f475732451;
reg         [MAX_SUM_WDTH_LONG-1:0]         I66d85c030a8864505298919046056305;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib869a349250a765d2f8660e0dbdcf312;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1a4fb631fdc7b5454c266589962ff5f0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9de4e0e86e9edcf948d9eddf0401b94a;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iee7b4838986c962969c00a0bbe53ce0b;
reg         [ 0:0]                   I9d9378337a77515a4e8d04fb88938808;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4841257ae596d9d3e4eb1e6f886956b0;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id81b11a8ca1dd8989e36cef637ae6aab;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibe96deab015b799fe7f69bae8432952c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I986b52155cc1470299321a4933241ed7;
reg         [MAX_SUM_WDTH_LONG-1:0]         I04be63a04f3942ce749cc9bd7540e055;
reg         [ 0:0]                   If0e20ef9aa69b77ae0e58ca3dfc9998f;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icd6f7ec117f9ab4eda8c5eba41386ffa;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia7adea5b0ec86e9fcd427a5468d72b64;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie8990d8abd23f8f9f79d7fe38c57fa8c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9d2f90ddddbdbb525d5f070f32546b64;
reg         [MAX_SUM_WDTH_LONG-1:0]         I905256d73bdb63bf860e15687350795f;
reg         [ 0:0]                   Iec2cb48bb1b58f268bf164d5e8a8120f;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibc0498839d1d9b6dc853b8e5d7a88fa3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9adcfc18e4471209edbe9a379e996067;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3d7d048348bf833f744a9f73889b7802;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id619e8d4040014d0e415ff71c5e0591f;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iaf3de2ef283e03dd72002026e1299224;
reg         [ 0:0]                   Ia4ae7c98720d43a604f28dfc5dd67d50;
reg         [MAX_SUM_WDTH_LONG-1:0]         I142ebca7f155e287e38ddf45423ab0fd;
reg         [MAX_SUM_WDTH_LONG-1:0]         I64551529c0028ec145407be7f5dfef71;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5ebe580a943b65fb16ea722ba101fd05;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0921901599c43b27e701758026dd3ee1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6033532f27c26b2d42bb3ea128f80dfa;

reg  [SUM_LEN-1:0]                         Ieb085b219090cde5da2190093ce43730;
reg  [SUM_LEN-1:0]                         Ib325dab091dfc3a1a269adb3ea9c75cd;
reg  [SUM_LEN-1:0]                         Ifc045af19c3f10d92d2b0dfb4fbbde38;
reg  [SUM_LEN-1:0]                         Ib79e305e6f44a4a6ebef1db5c70246ea;

localparam I0c5eab3e4dfde17a8c7261f7827e941c = 50;

reg [MAX_SUM_WDTH_LONG-1:0]    I43864225be03ea8e9379eb28dfa6c599;
reg [MAX_SUM_WDTH_LONG-1:0]    I31cb0c699cffcd2fedfbed0e1b86490e;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibed5004d869a01005768ba694c2234d6;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia4b2db3d48f946b0bfd0be0e32d7518d;
reg [MAX_SUM_WDTH_LONG-1:0]    I4d908bbe633c193cd9fc93dd33c60bd2;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib14733d3585dbf7f196cfc068e9508f0;
reg [MAX_SUM_WDTH_LONG-1:0]    Idfcf7f3240d92bfc87d44833bc00ff9d;
reg [MAX_SUM_WDTH_LONG-1:0]    I1cff7306aaf303bb3342ea3d72048908;
reg [MAX_SUM_WDTH_LONG-1:0]    I26bdcc44692db066911c8d5b0a1aae0c;
reg [MAX_SUM_WDTH_LONG-1:0]    Id144785da9b171f1e2d0e9182d693e31;
reg [MAX_SUM_WDTH_LONG-1:0]    I6b7a8ba12de5b44817ec99faebe54617;
reg [MAX_SUM_WDTH_LONG-1:0]    I4a403449a9ba75243369032e1cca1a0d;
reg [MAX_SUM_WDTH_LONG-1:0]    If85d9a95c1c02ce2da1dc3486b53eb81;
reg [MAX_SUM_WDTH_LONG-1:0]    I8e470b68bf35c647af42b6e46201e570;
reg [MAX_SUM_WDTH_LONG-1:0]    I484ec87270fcc959a486ebce40a9a03c;
reg [MAX_SUM_WDTH_LONG-1:0]    I079932780612fbce79cbe9b58bb6c2b5;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibb157b97546cb19fa7c1c0a7c79b1d38;
reg [MAX_SUM_WDTH_LONG-1:0]    I45cb51c25c426c296f97a5d23a08c063;
reg [MAX_SUM_WDTH_LONG-1:0]    Iff1d4b06901796098f91e87a3c30f7a5;
reg [MAX_SUM_WDTH_LONG-1:0]    I16db9cab1981451a02dab21e2ca221b4;
reg [MAX_SUM_WDTH_LONG-1:0]    I72756ea6a4997bc4afd4bfde1dfb2d26;
reg [MAX_SUM_WDTH_LONG-1:0]    I2882ae2eb6d79a5b96d1ed937dcfd8bf;
reg [MAX_SUM_WDTH_LONG-1:0]    I1a632a3e06ad738d5865acc77e204f48;
reg [MAX_SUM_WDTH_LONG-1:0]    I4d4ec5540257040d10182ed478a71918;
reg [MAX_SUM_WDTH_LONG-1:0]    I8da7e01f56dc9a70eb6b3f110dc005c2;
reg [MAX_SUM_WDTH_LONG-1:0]    Icc5d7bcbd7fcdb5092e6d8e18f6de6ec;
reg [MAX_SUM_WDTH_LONG-1:0]    I83cec264bd378f1dc23f87e439e7310e;
reg [MAX_SUM_WDTH_LONG-1:0]    Ied7e494fb288f78d110ed06662f1926a;
reg [MAX_SUM_WDTH_LONG-1:0]    Idd5b362dab4f93bba0c39af78c4c5981;
reg [MAX_SUM_WDTH_LONG-1:0]    Id033e7adfcfb0420cc592a1fb6c297b6;
reg [MAX_SUM_WDTH_LONG-1:0]    Iaee91a5e94c3f174682f72a1ebfd0021;
reg [MAX_SUM_WDTH_LONG-1:0]    I0cd8a6e719305ee3fbe8228081993957;
reg [MAX_SUM_WDTH_LONG-1:0]    I9b8cfdb69b76453a3ac687a1e098417f;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic2159627df2efa5e677fa6f4498bdd31;
reg [MAX_SUM_WDTH_LONG-1:0]    I59fba74472ded0a985cb237104ac127f;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia526539cc0f844b802d412b7a17cb6a6;
reg [MAX_SUM_WDTH_LONG-1:0]    I5d80b7c7d102d2c2bfa73a68c73376be;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia92defa0ca87c7c30fbe901da40a575e;
reg [MAX_SUM_WDTH_LONG-1:0]    I8fb1602dcdcd2912ea8aec42e2b7848f;
reg [MAX_SUM_WDTH_LONG-1:0]    I0cedca0e2c589104d6f3318505910594;
reg [MAX_SUM_WDTH_LONG-1:0]    I54c260db5c1b2c76527c8fc1cee229fe;
reg [MAX_SUM_WDTH_LONG-1:0]    I3d700e050cb7f22b0e381f3c72a20124;
reg [MAX_SUM_WDTH_LONG-1:0]    I63c0c8bef1dea4e499a16ce01e781951;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia8abcb8cf8d9ecc17c27ff015aa0b71f;
reg [MAX_SUM_WDTH_LONG-1:0]    I3f59174b3764a0b0741462024be9fb92;
reg [MAX_SUM_WDTH_LONG-1:0]    If0c2d002c315b21e11ae776bb48c9338;
reg [MAX_SUM_WDTH_LONG-1:0]    I18e548b082364c75686f2b7ad2ef46ab;
reg [MAX_SUM_WDTH_LONG-1:0]    I5e0d6b44474a226ab2ce916a6d46072a;
reg [MAX_SUM_WDTH_LONG-1:0]    I0c53d8d6a5b92960e29fc31cf456c23b;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib16c6096ce80e2f15a5ccea145e28510;
reg [MAX_SUM_WDTH_LONG-1:0]    I0e7ca2d6470b9bfc6a1ca6143b468507;
reg [MAX_SUM_WDTH_LONG-1:0]    I4ba05e74c2f63e2f4c59268775d549aa;
reg [MAX_SUM_WDTH_LONG-1:0]    Iaed26e1c4a2578d16b111d15d31339d2;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic566fe27ccaf2220101cbc49fc187a6b;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibf9f6d7baed9e761b69fb41442761ac6;
reg [MAX_SUM_WDTH_LONG-1:0]    Id5b4ee69444e5b499476c05a7f1d6e60;
reg [MAX_SUM_WDTH_LONG-1:0]    Id6105518ade80c89d4f20222a2382efb;
reg [MAX_SUM_WDTH_LONG-1:0]    I26cf25e680483bf4e556d74efec35ee7;
reg [MAX_SUM_WDTH_LONG-1:0]    I8636f5c91b567780d3324e4b8a320fc2;
reg [MAX_SUM_WDTH_LONG-1:0]    I914bef0326cf82d350344317eb1359be;
reg [MAX_SUM_WDTH_LONG-1:0]    I7de222bc26e38b8b6543819701740302;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie3361a270ebc41698ef4651bb3548a49;
reg [MAX_SUM_WDTH_LONG-1:0]    I1240c9410b897a4d0504affca5ba139e;
reg [MAX_SUM_WDTH_LONG-1:0]    If17b4f86674bc5fb212a1f7751fb043a;
reg [MAX_SUM_WDTH_LONG-1:0]    I275f6334127640b2de3f0f87f54fd74c;
reg [MAX_SUM_WDTH_LONG-1:0]    Iec844d10736440b96f9d6c651e604efd;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie04ce30f26a4ef1ee5b34474368dbac7;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibfee0b4ad5cdf16e88fcf469c5e031e9;
reg [MAX_SUM_WDTH_LONG-1:0]    I3a4a965f22487553dec2a3e8e7836264;
reg [MAX_SUM_WDTH_LONG-1:0]    I2a2d014f94d7a3b9fb3024a3e9107a73;
reg [MAX_SUM_WDTH_LONG-1:0]    I5bab5ae46114c487f67b8e779d7461df;
reg [MAX_SUM_WDTH_LONG-1:0]    I45373bff54eccf8137da2931d841934e;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib9322ec1d3866ba3cb42e96b5ff5cfb2;
reg [MAX_SUM_WDTH_LONG-1:0]    I0a9cb91319cc0d0c1c4d0020cce321d7;
reg [MAX_SUM_WDTH_LONG-1:0]    I299b37fd45c6ee2031fb2c74caac73be;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic2f450f7ab60ba57dfc1406c92c0f077;
reg [MAX_SUM_WDTH_LONG-1:0]    Ieca5b21b91e150c9d509964bdcea500d;
reg [MAX_SUM_WDTH_LONG-1:0]    I48b39ee498563e23c3a4be079b6100d8;
reg [MAX_SUM_WDTH_LONG-1:0]    Iac8cb32c2d86b975f51a2ed605002e51;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic989dc794ce4356856b3916ab1889589;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie380b37a78242e6d45b659d568887457;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie43a7f8082f91c2955076a6373028b55;
reg [MAX_SUM_WDTH_LONG-1:0]    Iea765ae5e9c65b3186445b15c56f69e5;
reg [MAX_SUM_WDTH_LONG-1:0]    I74b55d2f94073ba8f948e4b02386867c;
reg [MAX_SUM_WDTH_LONG-1:0]    I015630502f5cb4eb27b2a673e810f1dc;
reg [MAX_SUM_WDTH_LONG-1:0]    I5085f161323433d8d38be2e4511b0c46;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie9fd8f7dc0c3849c0437a2a3d8607b4c;
reg [MAX_SUM_WDTH_LONG-1:0]    I9306d9ef7934ffe5902306b9783c351e;
reg [MAX_SUM_WDTH_LONG-1:0]    I70e68beb262fbdeba621b3794adf9f84;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie7bf11bab3d601fd0a6e3eb415e263c8;
reg [MAX_SUM_WDTH_LONG-1:0]    Ica3d4ebff001fb6ee69a66eb898eb5bd;
reg [MAX_SUM_WDTH_LONG-1:0]    I27951ef3d612004abdc639662807426b;
reg [MAX_SUM_WDTH_LONG-1:0]    Ice4f4ba8bb3381c8846941d5d5fe4534;
reg [MAX_SUM_WDTH_LONG-1:0]    I223151b6414d9979d71023053dd3f5e2;
reg [MAX_SUM_WDTH_LONG-1:0]    I73d2731c1b1ae5ef73ce0eb9c8995912;
reg [MAX_SUM_WDTH_LONG-1:0]    I5ca15c7da1f49580ddedd9ff8ba822c0;
reg [MAX_SUM_WDTH_LONG-1:0]    I8289bfc08a5d8979ec26825bcb6e3d18;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie3c88bc240576aa220f0f110b13bfdd3;
reg [MAX_SUM_WDTH_LONG-1:0]    I583c6d23506c7d7b84403bfe977ec1ec;
reg [MAX_SUM_WDTH_LONG-1:0]    I768afe193d9d79b136736abc6846d945;
reg [MAX_SUM_WDTH_LONG-1:0]    I277d7065150714e33d8ba64875d18190;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia5c77c9be26d62b026f24ee5a5e25fb8;
reg [MAX_SUM_WDTH_LONG-1:0]    I88a325547ccfe4eabf90792abd60e356;
reg [MAX_SUM_WDTH_LONG-1:0]    I21842d06e25948ef461d1fd03485f86c;
reg [MAX_SUM_WDTH_LONG-1:0]    Id65f22fa8fc9c47bfd00c796b63c9fa4;
reg [MAX_SUM_WDTH_LONG-1:0]    I288ff69a7395e74f7de8da5a6a7f9062;
reg [MAX_SUM_WDTH_LONG-1:0]    I2ba94ef71f97b9ba731b306d4a5fd02c;
reg [MAX_SUM_WDTH_LONG-1:0]    I26ae9e570a101c6f8237d7941285b924;
reg [MAX_SUM_WDTH_LONG-1:0]    Icb92c7c10f0bfc5d287228f98d8a235c;
reg [MAX_SUM_WDTH_LONG-1:0]    Iba4972a3b71a3101ab23190ed905dc17;
reg [MAX_SUM_WDTH_LONG-1:0]    I33703f538ec70268e6c00ad6eef6c4e0;
reg [MAX_SUM_WDTH_LONG-1:0]    I71b93abe4b20e6a17ff17e0f33ac2ca5;
reg [MAX_SUM_WDTH_LONG-1:0]    I91c2f3cdd7cc98a60090ec6e46d52ae7;
reg [MAX_SUM_WDTH_LONG-1:0]    I4254f2987cd014ed703ae18e9963e585;
reg [MAX_SUM_WDTH_LONG-1:0]    I9068cca0de6ecff56ca542d0998fcab2;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib3ec015a3d43d46e0b7142b21a81cfee;
reg [MAX_SUM_WDTH_LONG-1:0]    I8cb171677016e4309034dc5d83981a48;
reg [MAX_SUM_WDTH_LONG-1:0]    I2a4b3573ae7c3b38ec34591f20c1d076;
reg [MAX_SUM_WDTH_LONG-1:0]    I276c2ce5d3a1b7551c2790971071b094;
reg [MAX_SUM_WDTH_LONG-1:0]    I9dff504e40aaddefedbb7b0f822c844a;
reg [MAX_SUM_WDTH_LONG-1:0]    I4ed5da534afbfe9ecbc10ef4cc649a55;
reg [MAX_SUM_WDTH_LONG-1:0]    I618363a8ac413dd0ee52eb658940eaed;
reg [MAX_SUM_WDTH_LONG-1:0]    I54166b387c02e12374d6febc425bfb7a;
reg [MAX_SUM_WDTH_LONG-1:0]    I0b6cdfa1dbfa774fc9a12d856e61cddb;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic4af6c9097257c9b22a57ce4b79b40fe;
reg [MAX_SUM_WDTH_LONG-1:0]    Iae21bdea20a6266d3f69aa680b6b2817;
reg [MAX_SUM_WDTH_LONG-1:0]    I37e360420c7dd061de93a6647513676d;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia81c31ea4f4786136b539c9766987596;
reg [MAX_SUM_WDTH_LONG-1:0]    I5a4f0749acdc34fd0786e4b3d062f88b;
reg [MAX_SUM_WDTH_LONG-1:0]    I5529d6db17b6184c45cc4487e5a2c24a;
reg [MAX_SUM_WDTH_LONG-1:0]    Iabe5aea929c668c9b9728d073ffb00c8;
reg [MAX_SUM_WDTH_LONG-1:0]    I4fb3fe065daa2708e55c812e57c19fb6;
reg [MAX_SUM_WDTH_LONG-1:0]    I4bd98e902e805426fdd4606fcb5a5214;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia5e26c2417aba1005971749f4ab2f367;
reg [MAX_SUM_WDTH_LONG-1:0]    I0e112f1d4e9c934a118f79f3856744a9;
reg [MAX_SUM_WDTH_LONG-1:0]    I005e8b590924f9486cb23191d35c9797;
reg [MAX_SUM_WDTH_LONG-1:0]    I8c5f98353b5b082dc3cf056469945a08;
reg [MAX_SUM_WDTH_LONG-1:0]    I9aa11f30712f1779339b985212a7979c;
reg [MAX_SUM_WDTH_LONG-1:0]    I65928407b1d5447dbc815cd2d2e7b37d;
reg [MAX_SUM_WDTH_LONG-1:0]    If5b3850da967f6f3d7a71d680341ad1c;
reg [MAX_SUM_WDTH_LONG-1:0]    I0aa5522190c741b7df4c4d7d34e46987;
reg [MAX_SUM_WDTH_LONG-1:0]    Iff777b2c4a3939e330c4cbb36cbe1ac5;
reg [MAX_SUM_WDTH_LONG-1:0]    I2d839c10960739097d449efab58b9fd4;
reg [MAX_SUM_WDTH_LONG-1:0]    Ice8765807beffd3acf59fa137ee0baac;
reg [MAX_SUM_WDTH_LONG-1:0]    I529eaa7e5eeb6d0a1aba78df5d5a2fa0;
reg [MAX_SUM_WDTH_LONG-1:0]    Icb2805685607d5fedd0300c9d800f863;
reg [MAX_SUM_WDTH_LONG-1:0]    Idadf072247b351cf51d718f797c3b375;
reg [MAX_SUM_WDTH_LONG-1:0]    I6fcb3b133a6a654b69f41468a713d922;
reg [MAX_SUM_WDTH_LONG-1:0]    I77e1f5f504a794edbb89c66cf1ffcf66;
reg [MAX_SUM_WDTH_LONG-1:0]    I185085cbf8da6df921ba32442b28bcca;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibcb80df5bed66f8498561e3f3ffa4ec4;
reg [MAX_SUM_WDTH_LONG-1:0]    I2cf5304a672431888916e08b3c15f0c7;
reg [MAX_SUM_WDTH_LONG-1:0]    Icf266f710358631b7119ef526acb301c;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia209e5b03deaf4fcb8ae12b731a49e0a;
reg [MAX_SUM_WDTH_LONG-1:0]    Iffb7fe9c74dfc01a43e99a099c4e7e04;
reg [MAX_SUM_WDTH_LONG-1:0]    I43f52bcba1bd2e8ee5fac03320e4f19f;
reg [MAX_SUM_WDTH_LONG-1:0]    I9fdfe73e77c384d33196c0f2d2a2fde2;
reg [MAX_SUM_WDTH_LONG-1:0]    I546657528d591e8bb44c32fed7707af5;
reg [MAX_SUM_WDTH_LONG-1:0]    I6e4ae763dc4e8aa8afc4599de96c75d3;
reg [MAX_SUM_WDTH_LONG-1:0]    Id8c36004ae8e550569a491f6b514945a;
reg [MAX_SUM_WDTH_LONG-1:0]    I111ac0aadbdd3e4479ca0786491a7b08;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib83242b57ab050b0e5f9bdf91fa118fb;
reg [MAX_SUM_WDTH_LONG-1:0]    I7be8b2f8a9fe8e13001c2a1fce4a8a3f;
reg [MAX_SUM_WDTH_LONG-1:0]    If4d030e5858f325debc6f37abf4a7d6c;
reg [MAX_SUM_WDTH_LONG-1:0]    I627e4bdc8061c69e3fcac17535b9f1e0;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia443284a35e0873de59b3ae55b7f809d;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibafedcf9f2990ed9c1efa973a0b1d81d;
reg [MAX_SUM_WDTH_LONG-1:0]    I439c7c302b535bfd7db655c3c607d71f;
reg [MAX_SUM_WDTH_LONG-1:0]    I2133d362ba45ceb3dceaa84e95ace1e6;
reg [MAX_SUM_WDTH_LONG-1:0]    I67534b68fee8f76ac0c5e64cd02aba42;
reg [MAX_SUM_WDTH_LONG-1:0]    I8613cac4ccd4f956e8a0ae7b627f5be2;
reg [MAX_SUM_WDTH_LONG-1:0]    I8493e2dac01f009db1d2d5504b49d135;
reg [MAX_SUM_WDTH_LONG-1:0]    I5c278aad08b7c4b0237d68f88fcb3f3a;
reg [MAX_SUM_WDTH_LONG-1:0]    Iba75ff0f3b67c7e28cf627706733d528;
reg [MAX_SUM_WDTH_LONG-1:0]    I9164fa2a9a33da6612ea692cf3fa7d2f;
reg [MAX_SUM_WDTH_LONG-1:0]    I0f3c4fb63ef1e88168b4d28175a0b68c;
reg [MAX_SUM_WDTH_LONG-1:0]    I99d236d41be79090ca7ba1fb6faaec4c;
reg [MAX_SUM_WDTH_LONG-1:0]    I487b9b236d118786e475ccc5e4e56a6d;
reg [MAX_SUM_WDTH_LONG-1:0]    I6cb09ac924c3b3b44443263e08c3315c;
reg [MAX_SUM_WDTH_LONG-1:0]    Id924dafd31fd0af0b28c7e6b7e95ec37;
reg [MAX_SUM_WDTH_LONG-1:0]    I9184110e3e9b8614460fc0abe5fff2d9;
reg [MAX_SUM_WDTH_LONG-1:0]    If8865fee7dbf593b34ea54692d947f10;
reg [MAX_SUM_WDTH_LONG-1:0]    I4854ff71aa885da3d07acaaa24740d7c;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie8befb003fe83e774e8d1d01d4e2f4ad;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie7e196fbb66ba6bee51ef0064ca519c2;
reg [MAX_SUM_WDTH_LONG-1:0]    I685699f60c76b00df87c9c53e9a8e448;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib6c0e635e659f54724737f0cffd1b0fc;
reg [MAX_SUM_WDTH_LONG-1:0]    I3a8bcfdab631a268d21c87b98e9d1c49;
reg [MAX_SUM_WDTH_LONG-1:0]    I3faeba79f7af7a006ab5cd256352e2db;
reg [MAX_SUM_WDTH_LONG-1:0]    I02e672436ade3ee620c72c0d9ceee664;
reg [MAX_SUM_WDTH_LONG-1:0]    I65708fb59e90bb79b8107da619fe63eb;
reg [MAX_SUM_WDTH_LONG-1:0]    I840a1a7c0bf49f4f42499b33f32fa02d;
reg [MAX_SUM_WDTH_LONG-1:0]    If7543e2f5a158b1f3f3a4078ec54cab5;
reg [MAX_SUM_WDTH_LONG-1:0]    I98a2aa729628adde0b6047869bd12743;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibfb57f2b507c27759a3556759f23977b;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib20dec1346f227042c749ec1abfa4d39;
reg [MAX_SUM_WDTH_LONG-1:0]    Ifba318d4faf308168c5eac8fe92395b4;
reg [MAX_SUM_WDTH_LONG-1:0]    I95b923444062b4a98918c685c65996d0;
reg [MAX_SUM_WDTH_LONG-1:0]    I45a6ef43e6e42594444adcbda26700ab;
reg [MAX_SUM_WDTH_LONG-1:0]    I508cea40d87bec2672f980d145c89b55;
reg [MAX_SUM_WDTH_LONG-1:0]    I0ace1d51fdee91f8f3826a945c4e66a4;
reg [MAX_SUM_WDTH_LONG-1:0]    I99ff3922e018c409dc8ce5f3503e3c56;
reg [MAX_SUM_WDTH_LONG-1:0]    I6a3824a6598bbaa138e1e763ad85f5f7;
reg [MAX_SUM_WDTH_LONG-1:0]    I283107989a436e2c720123b8d9e335c2;
reg [MAX_SUM_WDTH_LONG-1:0]    I7b12345fe53174cadef6811fb8869b42;
reg [MAX_SUM_WDTH_LONG-1:0]    Iac6fcccf3a0cfe04edc0d998b60c2681;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic9678deca4bf44a7b99f853334f6a05c;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie40c90fdb38b3e4046ba89295ed77d7c;
reg [MAX_SUM_WDTH_LONG-1:0]    Iea4a7766d3b9d5d030ade1739859ef0d;
reg [MAX_SUM_WDTH_LONG-1:0]    I844b9a89ffb7a5e48979fdea546e244a;
reg [MAX_SUM_WDTH_LONG-1:0]    I656852be6f5b3542862e0f68d48be518;
reg [MAX_SUM_WDTH_LONG-1:0]    Id6551b6b053952162b90792ab73a1a49;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib7fde6a2ec1ff0a3af10bccf3012e63f;
reg [MAX_SUM_WDTH_LONG-1:0]    I989091b3586964ab598f166a89279d16;
reg [MAX_SUM_WDTH_LONG-1:0]    I9785922874bba479ce4a9bf1759e2933;
reg [MAX_SUM_WDTH_LONG-1:0]    Ifbaae8b3da03911a4c96d4efdb9283c5;
reg [MAX_SUM_WDTH_LONG-1:0]    I77a54091bc2c3d9006ecb3471b94d8c8;
reg [MAX_SUM_WDTH_LONG-1:0]    I9859b94cda465ceaaa5674eb19e94824;
reg [MAX_SUM_WDTH_LONG-1:0]    I5a7746e9fbb8c009f83ae57423296cdf;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibddcc2e26fba20dfe2a2d399be2bc45b;
reg [MAX_SUM_WDTH_LONG-1:0]    I8dbe6497a8deabcc60783bfe7548d0fb;
reg [MAX_SUM_WDTH_LONG-1:0]    Ifef870b405335975988b58b2273d4e1a;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic1f6842b4f246d624d91daa6ada10ca9;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibc8679379ddc43ee4bc508a1f577eb2c;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibdd9957b7f1a319b797c021933ff75d7;
reg [MAX_SUM_WDTH_LONG-1:0]    I041f9455435bfa375395eb330a34993d;
reg [MAX_SUM_WDTH_LONG-1:0]    Ifbe29365e7035c78af9f42902b0d303e;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic8759e2f58848b33082bd1b02acc9c0b;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie2e3d64640c339dc51512979dbd6a173;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib2c327648cce481482eaf0467e9227d4;
reg [MAX_SUM_WDTH_LONG-1:0]    I535cad8c919a4330257eb5b4bed61b3a;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib2afdf9534deaae465d99b7e377788bb;
reg [MAX_SUM_WDTH_LONG-1:0]    I6eaffd980e4d77fdbda5e63bad9489d7;
reg [MAX_SUM_WDTH_LONG-1:0]    I6e4786234b286b12c83e06e93c628534;
reg [MAX_SUM_WDTH_LONG-1:0]    Idcc745602c4b7b34df9c3d68f9a9d76d;
reg [MAX_SUM_WDTH_LONG-1:0]    I0fc42ce9cc31d781ea3013318c25a571;
reg [MAX_SUM_WDTH_LONG-1:0]    I4363ca6b3d9ca9863f70958aa7c23777;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic902e09b33db1b919c102f7971cdef7b;
reg [MAX_SUM_WDTH_LONG-1:0]    Icf4405d4a4063448a2be8ad0354ab1a8;
reg [MAX_SUM_WDTH_LONG-1:0]    I72108531a608f6d5e51a481c68d7b271;
reg [MAX_SUM_WDTH_LONG-1:0]    I6922b510e432e06d209095bcc6297e7e;
reg [MAX_SUM_WDTH_LONG-1:0]    Ief90f8a8efca2b06eff0d4cba1cbb342;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib5334df42ee8f1574e41cb30b903fae9;
reg [MAX_SUM_WDTH_LONG-1:0]    I535b29f7177b4fc009ee998f1f4f7d7f;
reg [MAX_SUM_WDTH_LONG-1:0]    Id0842da8068ee88d99af7acea50e7b77;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib6cdbbb765694d822639b7c8fbfc50c4;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibdaa6d215d34aa0cc27d5234da6fd991;
reg [MAX_SUM_WDTH_LONG-1:0]    Id769d4a92f5f6da262ce0521e5509368;
reg [MAX_SUM_WDTH_LONG-1:0]    Iaf3a0b5ea5d9eda47fcced9260922bc6;
reg [MAX_SUM_WDTH_LONG-1:0]    I03a8a458ee0942c35001cbfe8e589222;
reg [MAX_SUM_WDTH_LONG-1:0]    I25eb943ea517a4827efb1e797bfdc4f5;
reg [MAX_SUM_WDTH_LONG-1:0]    Iac4b8906947fc90bfe76cee2f1d4c4ab;
reg [MAX_SUM_WDTH_LONG-1:0]    I58a490344f87b4d5bb319e3e85ba9278;
reg [MAX_SUM_WDTH_LONG-1:0]    I9222c4c0eb2b110fd80547d46ba17036;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic1af7410a9d11c5324f3ee5b2e0e9dac;
reg [MAX_SUM_WDTH_LONG-1:0]    I9e0a36d0be66b4c02b03e5b75b686226;
reg [MAX_SUM_WDTH_LONG-1:0]    I1eef40a71c8d1e2da9802929a5347e90;
reg [MAX_SUM_WDTH_LONG-1:0]    Ied41909cd443432dafadba42672151c1;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib2c1636a66f6479d6123a038cbc668d5;
reg [MAX_SUM_WDTH_LONG-1:0]    Ica02d19b129c8b1d491ea4747a55113e;
reg [MAX_SUM_WDTH_LONG-1:0]    I31bf4597a3b776962f5c820378254065;
reg [MAX_SUM_WDTH_LONG-1:0]    I58361fb97f1b5aff0a2751d35c8da672;
reg [MAX_SUM_WDTH_LONG-1:0]    I8ab7efc436a0f2cc3efbc299a0ddf914;
reg [MAX_SUM_WDTH_LONG-1:0]    I3934ed7170967ff3852944cc39ba1de9;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic690477b1672dea4905a5e1c92b47366;
reg [MAX_SUM_WDTH_LONG-1:0]    I5eaa11e26f19b94dcb7eaee7f09d24b4;
reg [MAX_SUM_WDTH_LONG-1:0]    Iaf1d3be13e6441a7a9ab3f286a7dc21b;
reg [MAX_SUM_WDTH_LONG-1:0]    I61f5ebea2bbe443b644c95ee559c2234;
reg [MAX_SUM_WDTH_LONG-1:0]    I1fbcaf2f6be01b129ebc24dee8a65396;
reg [MAX_SUM_WDTH_LONG-1:0]    I1c0df8c2c64b688ae417a238263f33db;
reg [MAX_SUM_WDTH_LONG-1:0]    I4f169c2c8c0768f2725ed655a03acfc2;
reg [MAX_SUM_WDTH_LONG-1:0]    I96f65790e2cacf7b529ce5b88598da00;
reg [MAX_SUM_WDTH_LONG-1:0]    I6b5720d71a0b4cd10ea34affa6631a25;
reg [MAX_SUM_WDTH_LONG-1:0]    Ifc7eec6765af08463751db128f8818b3;
reg [MAX_SUM_WDTH_LONG-1:0]    I8dddcade21ad3bb330c1c25970c32b73;
reg [MAX_SUM_WDTH_LONG-1:0]    I74a7b85ddacad06ab1c6b0db9b084bd3;
reg [MAX_SUM_WDTH_LONG-1:0]    I2b0b168ce4fe8aa4a2e7cb69fe532aa3;
reg [MAX_SUM_WDTH_LONG-1:0]    I3e8d26ea83937cae01aadf1092c59bdf;
reg [MAX_SUM_WDTH_LONG-1:0]    I90a4190941651d885d04deb86a163365;
reg [MAX_SUM_WDTH_LONG-1:0]    I7d85b73e85379bf3a480e954c05516f3;
reg [MAX_SUM_WDTH_LONG-1:0]    Id5c9a9b9c34c8f9d56df0aa8d780c9d3;
reg [MAX_SUM_WDTH_LONG-1:0]    I21255a0ad20a9668c958faf68d53b2bc;
reg [MAX_SUM_WDTH_LONG-1:0]    Ifba1584d599da13b98a3b76b4db10974;
reg [MAX_SUM_WDTH_LONG-1:0]    Iad0f4602ec545dc6ef12aa34add00ed3;
reg [MAX_SUM_WDTH_LONG-1:0]    I8bb46c3eb9f54c5d1b28dc6aa0154358;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic09b4671e867144fe9f54a09e74c5519;
reg [MAX_SUM_WDTH_LONG-1:0]    I391a2f354262558ff17d7d80b8c39e8c;
reg [MAX_SUM_WDTH_LONG-1:0]    If6b40a030cb120fe017bf9d39e1a35d1;
reg [MAX_SUM_WDTH_LONG-1:0]    I490996026af34eba5bcd8d553af818eb;
reg [MAX_SUM_WDTH_LONG-1:0]    Icbc12ab47f586b12402ae5d4361c967d;
reg [MAX_SUM_WDTH_LONG-1:0]    Iee0e45914c52a357e1e32922299d6937;
reg [MAX_SUM_WDTH_LONG-1:0]    Iefe423653d454e21324a6857b52f98ac;
reg [MAX_SUM_WDTH_LONG-1:0]    I6d6a242cdfadfc97fe656510bef73adc;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib5c8d91204a2d313c9c23110a53cd0cf;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic9740baafb1c92e3a25f0a1e7bc46486;
reg [MAX_SUM_WDTH_LONG-1:0]    I6f69796a6fe6da57066319ec8210c1a3;
reg [MAX_SUM_WDTH_LONG-1:0]    Idb862697f62a6c678072de760e176096;
reg [MAX_SUM_WDTH_LONG-1:0]    I06e05a1ed002175a75d02b8b76f52c50;
reg [MAX_SUM_WDTH_LONG-1:0]    I1e110e27162231650875dd1152d96e64;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic46357bb77f6183329946f7e28294365;
reg [MAX_SUM_WDTH_LONG-1:0]    I8741c5cc763512d16cb1186fa3323f45;
reg [MAX_SUM_WDTH_LONG-1:0]    I30b5c7aadb5312ce96e833704bb3a320;
reg [MAX_SUM_WDTH_LONG-1:0]    If404a00ab81d6ebbc0dbdf4aecdce389;
reg [MAX_SUM_WDTH_LONG-1:0]    I19875f52f79482b477f1febaa7e97090;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic7855ca956651bd368cbdde7ec93ba6d;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic57a2627a194099105a2908a41feddfb;
reg [MAX_SUM_WDTH_LONG-1:0]    I4d1ba6ee8fb9505ba3b58b2b7553245b;
reg [MAX_SUM_WDTH_LONG-1:0]    Ieb7b388ff89e352dd239e0ccbe7b9ecc;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib1461f456ebc14f449eee77e386a4c69;
reg [MAX_SUM_WDTH_LONG-1:0]    I8786eb767f02164cdc32f14f41b5d0e1;
reg [MAX_SUM_WDTH_LONG-1:0]    Id6fa8ec5d1062fc3e09bdac65ff79f45;
reg [MAX_SUM_WDTH_LONG-1:0]    I83b77ad1a40dc102f28153f692516eb4;
reg [MAX_SUM_WDTH_LONG-1:0]    I55e54359961ef6e5a63f1c2eb0ad4aa1;
reg [MAX_SUM_WDTH_LONG-1:0]    I90001da8c360ccff128f637cd672ad42;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib38a46dc131d635b81fb7c196110fc4b;
reg [MAX_SUM_WDTH_LONG-1:0]    I926c049036f53f0a0a6ad369de116c57;
reg [MAX_SUM_WDTH_LONG-1:0]    Iac48d2ccf6c6e0c555e874ae77123f2e;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic6f40833f5f6284c9015304fd3fc00f0;
reg [MAX_SUM_WDTH_LONG-1:0]    I3f2507530dd648814af0964f7da11d35;
reg [MAX_SUM_WDTH_LONG-1:0]    Id9edc6ac95a260bf5af3de25f00e9e9c;
reg [MAX_SUM_WDTH_LONG-1:0]    I28fa295ebd90c2b7255d48ca9ffcfcf3;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia308e09137af1cb50167562efb5da628;
reg [MAX_SUM_WDTH_LONG-1:0]    I5aa85d9503b0e4ff46bbd63e873053ca;
reg [MAX_SUM_WDTH_LONG-1:0]    I7ea8fe50c45e213f3257060e2813240b;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic3e6e38a2986c7f14fd0db2246367a1c;
reg [MAX_SUM_WDTH_LONG-1:0]    I581eb136fdd08302e02c1fafb5d5c90b;
reg [MAX_SUM_WDTH_LONG-1:0]    I080832c25509f7003ed50d71210bc7f7;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib43383830037df764b48c637a28ab6b5;
reg [MAX_SUM_WDTH_LONG-1:0]    Iddf65ccb4396288264a400ba37cbb655;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia7673d73f0535906a99d6cb467892104;
reg [MAX_SUM_WDTH_LONG-1:0]    I8bc3210e86a523accdbeefe7e72ee4fc;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib63574478126e6ee30a388d9648cb548;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic4501a8a1fb34c30a97e18a0ab189e3a;
reg [MAX_SUM_WDTH_LONG-1:0]    I2b807c16cfc6d65cb2a7f28ffa837974;
reg [MAX_SUM_WDTH_LONG-1:0]    I0aa93075086164fdbab3814d60633141;
reg [MAX_SUM_WDTH_LONG-1:0]    I886750aaf8d2040c3f12ff113294f658;
reg [MAX_SUM_WDTH_LONG-1:0]    I103ec7cf279f527fc6e3648a19a12a8a;
reg [MAX_SUM_WDTH_LONG-1:0]    I9a57f2f03cf8a154c3a7d48ec089306d;
reg [MAX_SUM_WDTH_LONG-1:0]    I9d8f8c1792427975a9e7024041f59be9;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie8644d7edbadf19937c399cf275946e5;
reg [MAX_SUM_WDTH_LONG-1:0]    I2b32537c9178028493af165398a60875;
reg [MAX_SUM_WDTH_LONG-1:0]    If06a1563b9d7348de03a98d31bd85b06;
reg [MAX_SUM_WDTH_LONG-1:0]    I58a7c7b05b84d292cd06d68e96ecb9f8;
reg [MAX_SUM_WDTH_LONG-1:0]    I3fdec80112b3fc543b217d1c253406da;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia1aedd38250e76763aaee3de2f832b3c;
reg [MAX_SUM_WDTH_LONG-1:0]    I2087576fbc15119bf5d9e8afa2603b69;
reg [MAX_SUM_WDTH_LONG-1:0]    I7a6ab9e700bd94208ab6528af413f3a9;
reg [MAX_SUM_WDTH_LONG-1:0]    I4481555c402ba99bee05658ba6017984;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib849494e5087777f646ee0947b4f634a;
reg [MAX_SUM_WDTH_LONG-1:0]    I18d0dd7a10d6533f721a2392d4ad2d02;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib8603cb82ceb97c2f35bf8209306a457;
reg [MAX_SUM_WDTH_LONG-1:0]    I2418ae211f327ed45cc70c42078180dc;
reg [MAX_SUM_WDTH_LONG-1:0]    I6521c9167261db6eb37f50b66159ddb7;
reg [MAX_SUM_WDTH_LONG-1:0]    I920f95bb52cdc9b07f93afc3a6b5c009;
reg [MAX_SUM_WDTH_LONG-1:0]    Iad0ecc5208263d239e4a62c5563f52ab;
reg [MAX_SUM_WDTH_LONG-1:0]    I0c0be3347a7df9cc39997208b013f17b;
reg [MAX_SUM_WDTH_LONG-1:0]    I70dc03a46e1ac0da826388abd3bdc503;
reg [MAX_SUM_WDTH_LONG-1:0]    I452ba61d5fb5c7ead1824dade4bd7801;
reg [MAX_SUM_WDTH_LONG-1:0]    I8b5d10c412daccdcb07645bf239d61bd;
reg [MAX_SUM_WDTH_LONG-1:0]    I9b1390839ee2b9ba591e3873e967c8e2;
reg [MAX_SUM_WDTH_LONG-1:0]    I17e818b67440efaba9a5d19e7467bf85;
reg [MAX_SUM_WDTH_LONG-1:0]    Ifa67d343acc6f3ec50c2b01fc26b4374;
reg [MAX_SUM_WDTH_LONG-1:0]    If0676ef300628c4097565b13ef2d8854;
reg [MAX_SUM_WDTH_LONG-1:0]    I8d26e73fafa909f1e26e329828cf4888;
reg [MAX_SUM_WDTH_LONG-1:0]    If29fcea810adbdb1c4d8a4ace1d8081b;
reg [MAX_SUM_WDTH_LONG-1:0]    I0e3286fca6cd040758950259ab663df7;
reg [MAX_SUM_WDTH_LONG-1:0]    I696db0b98e27dcc4657dc7feb23a881b;
reg [MAX_SUM_WDTH_LONG-1:0]    I06c0921675f464807a63c7965796f0d0;
reg [MAX_SUM_WDTH_LONG-1:0]    If36016df78d833c80e1355151c038225;
reg [MAX_SUM_WDTH_LONG-1:0]    I0dbf900b4f430b4c1106aa86b640bb37;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib8664a2abe9d6326d6e45bb2a7ad59d0;
reg [MAX_SUM_WDTH_LONG-1:0]    I91893028c4409cfeceeb7976815b2d31;
reg [MAX_SUM_WDTH_LONG-1:0]    I2e14fb1e667e967ab4c116e0c7438aec;
reg [MAX_SUM_WDTH_LONG-1:0]    I0fb60c4f56f6d7b4007cf0dae39f4573;
reg [MAX_SUM_WDTH_LONG-1:0]    I24b4c998d19ae97f7178e37f75c77d06;
reg [MAX_SUM_WDTH_LONG-1:0]    Idb73eba1bd4ce25a6109e296f51e7dc4;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibc1a16427d8dfa5ee20dac15327a53ea;
reg [MAX_SUM_WDTH_LONG-1:0]    I0e52c25aa840402d944cbd81f73c1ffe;
reg [MAX_SUM_WDTH_LONG-1:0]    Id7619819e1297844d92c8bf3a1d61926;
reg [MAX_SUM_WDTH_LONG-1:0]    Idfa432a87877e1ce103e56891745b62a;
reg [MAX_SUM_WDTH_LONG-1:0]    I13b9e098622d90a1074f636d8f351aca;
reg [MAX_SUM_WDTH_LONG-1:0]    I78e1205de9119fac3ae8f43c72ac71f4;
reg [MAX_SUM_WDTH_LONG-1:0]    I5bbbc4eedb7c61516769f429a8498ea7;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia1d9dee7a9821283498d17de0cfacb32;
reg [MAX_SUM_WDTH_LONG-1:0]    Idd8643af2515f65fd9a1dfe66494ccf2;
reg [MAX_SUM_WDTH_LONG-1:0]    I1684820afb9d9cec38cfdfcd6ca8b36a;
reg [MAX_SUM_WDTH_LONG-1:0]    Ice8a82bdd966719098a8d5f2a826f73d;
reg [MAX_SUM_WDTH_LONG-1:0]    I338400586daa58006c0a3dcd82ea8f4a;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie467c5fde1d123da4e9587b5a56748a0;
reg [MAX_SUM_WDTH_LONG-1:0]    Ifc52604a4f9f9de392a35f2f9fe885b8;
reg [MAX_SUM_WDTH_LONG-1:0]    I20c4e393929b875521e5316f4d8e2d42;
reg [MAX_SUM_WDTH_LONG-1:0]    I064499f0315fbeec7b6cb50583388a07;
reg [MAX_SUM_WDTH_LONG-1:0]    I894ef04bfa1b7b39ef51b7c82f7686eb;
reg [MAX_SUM_WDTH_LONG-1:0]    I8d6927b0bcbbb318cf52987c121a07b5;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie0ce2826fd13b0e0b23c91e97787691f;
reg [MAX_SUM_WDTH_LONG-1:0]    I7dbd1aeba00bb8b257990b7bb294211f;
reg [MAX_SUM_WDTH_LONG-1:0]    Id5ddf5331aba567aaf5b7eb88b31a52e;
reg [MAX_SUM_WDTH_LONG-1:0]    I0f46a17f14ab18e6338aa3d06678b0a5;
reg [MAX_SUM_WDTH_LONG-1:0]    If1ec4241fd12255369f72b3f3310b6e7;
reg [MAX_SUM_WDTH_LONG-1:0]    Iedf37dac8b3a5331277ae4f0176968aa;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia422fbdf8f318ff3ddc049d1374e7939;
reg [MAX_SUM_WDTH_LONG-1:0]    I9cbe73d708c561d43d05945552d32dde;
reg [MAX_SUM_WDTH_LONG-1:0]    I7e36dcae438a712fca2320117b7e3356;
reg [MAX_SUM_WDTH_LONG-1:0]    I0f9bc36c9d40290f83489aac3d674924;
reg [MAX_SUM_WDTH_LONG-1:0]    I3a09554ca009781e28ef1b3ea70d39ad;
reg [MAX_SUM_WDTH_LONG-1:0]    I28ea268c5b51ac1d9249e96599bb6b0d;
reg [MAX_SUM_WDTH_LONG-1:0]    I1d648ed8f07f0743a6d616584270c513;
reg [MAX_SUM_WDTH_LONG-1:0]    I82a225237aeb1ceb31e8cd18b1e45c6f;
reg [MAX_SUM_WDTH_LONG-1:0]    I36ed1a0d0d618f90443fbea17b7c97ec;
reg [MAX_SUM_WDTH_LONG-1:0]    I612a41511db375f10f3c2b10d13edb24;
reg [MAX_SUM_WDTH_LONG-1:0]    I19032091a26dfdfffff60818041ec79e;
reg [MAX_SUM_WDTH_LONG-1:0]    I6aba8ca0e4b20a6355b43a70f19d9d8c;
reg [MAX_SUM_WDTH_LONG-1:0]    I839895c8614ff28df83314c44824900b;
reg [MAX_SUM_WDTH_LONG-1:0]    I8cbafa797ef136d7e50c909dc160deb1;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibac0851ce1a3c23f18b072d263afff36;
reg [MAX_SUM_WDTH_LONG-1:0]    Id58474582f209a3859f65a447fe99191;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic9e06a355beabfacc053ec48f17f49de;
reg [MAX_SUM_WDTH_LONG-1:0]    I77fd8001d879fc9e9117464fba27902d;
reg [MAX_SUM_WDTH_LONG-1:0]    I2a0dc4ed573a544cb13544e049514903;
reg [MAX_SUM_WDTH_LONG-1:0]    I71bc7271cc432bb3c5d0b7a416cdfc60;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib76e892d1a1271844338042381b5690b;
reg [MAX_SUM_WDTH_LONG-1:0]    Icb158c031d434cb419c15e0510511231;
reg [MAX_SUM_WDTH_LONG-1:0]    I563802213afb6abe2f6e8c6f4d1e5b08;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia5b779ef95333736b08f63770900e275;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic1120eb027841908cd64fe5c7274da14;
reg [MAX_SUM_WDTH_LONG-1:0]    I5160de2c5ce4782d8f8be10dc740694b;
reg [MAX_SUM_WDTH_LONG-1:0]    I5f7b6e6a30348ae86057f7e56f625846;
reg [MAX_SUM_WDTH_LONG-1:0]    I9de41d0b279b84366640880dbd18c502;
reg [MAX_SUM_WDTH_LONG-1:0]    Ifec9abca21cf476b70e0befa3926b46a;
reg [MAX_SUM_WDTH_LONG-1:0]    Ifc527b6af9486df7f52d7eb9637c671f;
reg [MAX_SUM_WDTH_LONG-1:0]    I31d94aae2e3721045fe850d84dd2225a;
reg [MAX_SUM_WDTH_LONG-1:0]    If3bdbb4c20efca0c5af78614b4271ed1;
reg [MAX_SUM_WDTH_LONG-1:0]    I4037f1b207aa101f354e59eddd7c9eb4;
reg [MAX_SUM_WDTH_LONG-1:0]    If4d63635a5f99c4dc9e5b57712830c20;
reg [MAX_SUM_WDTH_LONG-1:0]    I1f1f2fefd3381ee48ab0ec9c9301754b;
reg [MAX_SUM_WDTH_LONG-1:0]    Iba52b84e6e215842e0ca8e72c42ebce7;
reg [MAX_SUM_WDTH_LONG-1:0]    I597c3f5c14e235f90dc8c796bc3e931d;
reg [MAX_SUM_WDTH_LONG-1:0]    I397a69dab323c7148b620dd6fe0b0c51;
reg [MAX_SUM_WDTH_LONG-1:0]    I401ab1ad994f5018061a3f57d3a51ad1;
reg [MAX_SUM_WDTH_LONG-1:0]    I3a47540f34ce47bcfa1da66cc4e6e088;
reg [MAX_SUM_WDTH_LONG-1:0]    I18916d0023ca275d84c52af07dcc5ca2;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic79072d9e42dbc9974231f1d642b3f12;
reg [MAX_SUM_WDTH_LONG-1:0]    I1140fa91b5e22ba0c094c03295781e5a;
reg [MAX_SUM_WDTH_LONG-1:0]    Id2989aaee3930698cd374e6c9feedf82;
reg [MAX_SUM_WDTH_LONG-1:0]    Icda9a86a25dbe516a93b46fe487029e3;
reg [MAX_SUM_WDTH_LONG-1:0]    I53971b75cbd7ebc74b579776a6ea4778;
reg [MAX_SUM_WDTH_LONG-1:0]    I37e5c3118e8536e37bd797aeaa92476c;
reg [MAX_SUM_WDTH_LONG-1:0]    I9c68bfa3b888b6a6d41e38e674578284;
reg [MAX_SUM_WDTH_LONG-1:0]    I2c72d6c5fa6968dffa6517cf81219875;
reg [MAX_SUM_WDTH_LONG-1:0]    I9bb4d58b1fe80549451b00c4ed2b3885;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic488e78b5c73251b673301e84c4b5b0b;
reg [MAX_SUM_WDTH_LONG-1:0]    I8d07beccef519ab4ce4024d911ac2346;
reg [MAX_SUM_WDTH_LONG-1:0]    I7c191c2c2be09886d0f31e4368797afd;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia3bfd86e26efbef2cf6bb72be7ac1453;
reg [MAX_SUM_WDTH_LONG-1:0]    I4ae59dd2f57bda295e11b077e8668f1a;
reg [MAX_SUM_WDTH_LONG-1:0]    I3f6fad8bb0fba790fcdb1612b6fa7712;
reg [MAX_SUM_WDTH_LONG-1:0]    I58416287b268462d28f55c6c2705e613;
reg [MAX_SUM_WDTH_LONG-1:0]    I106d0e71b7378d110b0a624e5cbf0d6e;
reg [MAX_SUM_WDTH_LONG-1:0]    I59adad4fd84c1fc233dc58f70a12779d;
reg [MAX_SUM_WDTH_LONG-1:0]    I8e01532a1ab9534b8de0474549d41a2e;
reg [MAX_SUM_WDTH_LONG-1:0]    I80af3dcb716f3474a7257700aef89b81;
reg [MAX_SUM_WDTH_LONG-1:0]    I07d68462362d8453e83570cc793c55db;
reg [MAX_SUM_WDTH_LONG-1:0]    I9a2bba3f62de5f750dc8161a488dc331;
reg [MAX_SUM_WDTH_LONG-1:0]    I71da7e172b2b967040b6e6d02ef9949e;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib97b2670a6cd88b2327f07f62d887900;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib2963b82260024e1853d297798d88d3c;
reg [MAX_SUM_WDTH_LONG-1:0]    I0722ec4e9d400f8eaeacd060e42de79c;
reg [MAX_SUM_WDTH_LONG-1:0]    I1972375d51767f0cffa5395a354b3493;
reg [MAX_SUM_WDTH_LONG-1:0]    Ifb19d75cfa0051107b5fba57bfc002b5;
reg [MAX_SUM_WDTH_LONG-1:0]    I9d05dc0e39e85c23b62f343a8de12e64;
reg [MAX_SUM_WDTH_LONG-1:0]    I64ae3cd6f36b8bde29cd3e1fcba7bade;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia6a78664c080829664158f53ba330312;
reg [MAX_SUM_WDTH_LONG-1:0]    I2ba16a10a82c20d54c776a9804ee50e4;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie9a316de516ec4fb828a614c67e38b2a;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie945349d77442536992d9ad52ce84218;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic6a7a82d16e6106071934ba79d3698cd;
reg [MAX_SUM_WDTH_LONG-1:0]    Ide40b1bf9c0b642c49a5685a62af1c93;
reg [MAX_SUM_WDTH_LONG-1:0]    I79280400a4c9bed015106e5d006de757;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic6e3847f035738243f4c5f71f296da57;
reg [MAX_SUM_WDTH_LONG-1:0]    I45b64b2b963963d2d0a8318133941f1d;
reg [MAX_SUM_WDTH_LONG-1:0]    I1939152ddbede923cde577984e0aa743;
reg [MAX_SUM_WDTH_LONG-1:0]    Ifbcebda2bb0ce58a0e1764c392a816df;
reg [MAX_SUM_WDTH_LONG-1:0]    I6d0d098e6d47dea04d6d7be67b648a0d;
reg [MAX_SUM_WDTH_LONG-1:0]    Icaeb9a2ec8ec5822658fa85b88cca04b;
reg [MAX_SUM_WDTH_LONG-1:0]    I3cc30aaba3dcd3eda262a19e85e53117;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic0b2f9717b8aacb34325fd5aaf03a366;
reg [MAX_SUM_WDTH_LONG-1:0]    I002869e450d79649d27441ce00bfb575;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie4d20df6b1e7a42f0df9a3cc26b12ac1;
reg [MAX_SUM_WDTH_LONG-1:0]    Idd01d014f0469f893305057ae3f4cb2e;
reg [MAX_SUM_WDTH_LONG-1:0]    I79444eef1875b6ad1a0675b66392ff9d;
reg [MAX_SUM_WDTH_LONG-1:0]    I7caf8c7496dd96c1ed08e98b415f5775;
reg [MAX_SUM_WDTH_LONG-1:0]    I7fc6e2aecff5bd691872d1e10a39103b;
reg [MAX_SUM_WDTH_LONG-1:0]    I49321308413cb4dbe5e6c01ba5b9023c;
reg [MAX_SUM_WDTH_LONG-1:0]    Id27560fb44b4f2fda98d47e9f20d6898;
reg [MAX_SUM_WDTH_LONG-1:0]    I745187336b8a5ae4eac66e90539752cf;
reg [MAX_SUM_WDTH_LONG-1:0]    I772e844c41387e7079259875e0ba3fa0;
reg [MAX_SUM_WDTH_LONG-1:0]    I32c35da92922c5b477f8aba837fa6d92;
reg [MAX_SUM_WDTH_LONG-1:0]    I3bc01b072987a0c980615abbc2251e5f;
reg [MAX_SUM_WDTH_LONG-1:0]    If08adda7d796da7c7849e472a73282a3;
reg [MAX_SUM_WDTH_LONG-1:0]    Ife3bb8945e14d8746c82b66886293997;
reg [MAX_SUM_WDTH_LONG-1:0]    I45ef0ac486fe043f57e8a46aa91461a3;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic0ae1191869e636f9e4391efe93309ae;
reg [MAX_SUM_WDTH_LONG-1:0]    Id92d779518ae724b5fef5221372f8f26;
reg [MAX_SUM_WDTH_LONG-1:0]    Id0762ac7710c93249bc11c6ce4ae51a0;
reg [MAX_SUM_WDTH_LONG-1:0]    Ife6be241bc50560a14f97650e5cc2959;
reg [MAX_SUM_WDTH_LONG-1:0]    I1062442edb2bff727ca6283c8270bf28;
reg [MAX_SUM_WDTH_LONG-1:0]    I6c9ae8b8191507f908c27bbde53bf2d5;
reg [MAX_SUM_WDTH_LONG-1:0]    Iec936eeebd1f8c95307bd8705e6def81;
reg [MAX_SUM_WDTH_LONG-1:0]    I6332af145d560e3f22a4a88106749f98;
reg [MAX_SUM_WDTH_LONG-1:0]    I0c121fa3e9e6e0e2e8291a594d6b4ceb;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic3c59a5167cb83fd76ec6236572b1f3d;
reg [MAX_SUM_WDTH_LONG-1:0]    I3e8e280553edaa5c8555ace81ecc10e0;
reg [MAX_SUM_WDTH_LONG-1:0]    I3e466d40a4447a23953d96d2e6d61d47;
reg [MAX_SUM_WDTH_LONG-1:0]    I76e4c55148effeba62a4837cd19c5e51;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie335e68643fd2b0a53351f4bd45c3475;
reg [MAX_SUM_WDTH_LONG-1:0]    I89f75107ea95f207b9e664a1f4f0746a;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic8f0049e1298b14b4e039075dc0d5f74;
reg [MAX_SUM_WDTH_LONG-1:0]    I382153cec6f7d6258574e7c532186473;
reg [MAX_SUM_WDTH_LONG-1:0]    I351dc309e916f282cc1e19303eee4112;
reg [MAX_SUM_WDTH_LONG-1:0]    I9de5e90485b3f22e9003dc8a7b22a79b;
reg [MAX_SUM_WDTH_LONG-1:0]    Idc4171a40dd2470e852af37a461013c7;
reg [MAX_SUM_WDTH_LONG-1:0]    Ifae488cb68d95ea517376319eb11f1bf;
reg [MAX_SUM_WDTH_LONG-1:0]    I9cab38b69794ab661e12750cf69c822c;
reg [MAX_SUM_WDTH_LONG-1:0]    I24180fba17c21bacefa8a4514e4b685c;
reg [MAX_SUM_WDTH_LONG-1:0]    I83bbe6fa947f9f909e1a6785ab31901f;
reg [MAX_SUM_WDTH_LONG-1:0]    I202c385beeccee309104b66f8f096b2c;
reg [MAX_SUM_WDTH_LONG-1:0]    Idc549661d6694035874a3366704801c7;
reg [MAX_SUM_WDTH_LONG-1:0]    I778fbaea65beeb6de599490daf3b7e3c;
reg [MAX_SUM_WDTH_LONG-1:0]    I4fd45670f88265e5d7aa6582f3ad3ff8;
reg [MAX_SUM_WDTH_LONG-1:0]    I2d636a246d815a4d12c478794860dd40;
reg [MAX_SUM_WDTH_LONG-1:0]    I3319313fe1d2b4ec2626711b187b4a5a;
reg [MAX_SUM_WDTH_LONG-1:0]    I586aaa5c55efd37996b01febd3bc60a4;
reg [MAX_SUM_WDTH_LONG-1:0]    I95ccc219b5f5038641b38dff6db0b222;
reg [MAX_SUM_WDTH_LONG-1:0]    I5001118df37d08bd19d322aca8ff3996;
reg [MAX_SUM_WDTH_LONG-1:0]    I22c15857572603cc24d8a87cb47c33b0;
reg [MAX_SUM_WDTH_LONG-1:0]    Ifdcd91f925b63e0817798aa6e9200e50;
reg [MAX_SUM_WDTH_LONG-1:0]    I8435e69bc1ff06e7edfabbee7b9aa49e;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibeff607ba15fd8ef504224a9c1d102fc;
reg [MAX_SUM_WDTH_LONG-1:0]    Id15c3bdce785df234c68432ccec8f959;
reg [MAX_SUM_WDTH_LONG-1:0]    I25888aa2135fc403ca9eac4df634549a;
reg [MAX_SUM_WDTH_LONG-1:0]    I632ffd09a9091335b3aa91ab2a8f1cce;
reg [MAX_SUM_WDTH_LONG-1:0]    I283331db80e6d0891b13dc55e6a7d76c;
reg [MAX_SUM_WDTH_LONG-1:0]    I134a734d93e62f6ac6635015fe3a2096;
reg [MAX_SUM_WDTH_LONG-1:0]    Id66798f8ea67e74a67f264fe6b4503a3;
reg [MAX_SUM_WDTH_LONG-1:0]    If2ce7b8d2573494564393f7d426fa47f;
reg [MAX_SUM_WDTH_LONG-1:0]    Id59cf860d9f4aff11b205b8970d93df3;
reg [MAX_SUM_WDTH_LONG-1:0]    I75aaeab4f372e28a8e51453540f9c6b2;
reg [MAX_SUM_WDTH_LONG-1:0]    I2266afbacf1ba750ce18f296aba1181d;
reg [MAX_SUM_WDTH_LONG-1:0]    I69c2b063e61e14f5d49b907095ece00f;
reg [MAX_SUM_WDTH_LONG-1:0]    If077c67a062095cfe69f2260cee82833;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibc03a9b6115d0941ce9233df7ef2fa57;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia18bdb8d2f02b50281f0acd4a45ac973;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib88c884e54d6e6ecf5ac015bc304e4f3;
reg [MAX_SUM_WDTH_LONG-1:0]    If6f5efee5e1f9709d86bf28cfb741955;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia0caf6693d441ac622f416a86b665166;
reg [MAX_SUM_WDTH_LONG-1:0]    I85dd6a9634284c22027b4241551ea628;
reg [MAX_SUM_WDTH_LONG-1:0]    Id5cedaa397ebfc2567efcc2f8a648db5;
reg [MAX_SUM_WDTH_LONG-1:0]    Ica0a119af1728ae253c16cc3eb93f802;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie7274a7ffa053ced4f12a67986d3c81b;
reg [MAX_SUM_WDTH_LONG-1:0]    Ife7985db888089ea618413810611bfca;
reg [MAX_SUM_WDTH_LONG-1:0]    If49068db99aa9d09302eda27ab51fcb7;
reg [MAX_SUM_WDTH_LONG-1:0]    I2959f2dc554e599d675eb6912757e413;
reg [MAX_SUM_WDTH_LONG-1:0]    I898d1b59aab3d5d4adce8ec3c0e14a0d;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibb6e54edb9d277242c06d386a9a75a26;
reg [MAX_SUM_WDTH_LONG-1:0]    I51b1cd475d0e389326b182cbe680a402;
reg [MAX_SUM_WDTH_LONG-1:0]    If12366160fdc899bd71cb0de5bcfd84d;
reg [MAX_SUM_WDTH_LONG-1:0]    I44e5ce0cdf812c5b73e6e638da36e414;
reg [MAX_SUM_WDTH_LONG-1:0]    I4f38c3d620b72f21cf6d54c7df4ba816;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib66b897398ea0702b74bdd03774f3ae4;
reg [MAX_SUM_WDTH_LONG-1:0]    I0b3a936c3f7e0391111e696b2445803b;
reg [MAX_SUM_WDTH_LONG-1:0]    I10f045edf47784a91a5599494c2d3de2;
reg [MAX_SUM_WDTH_LONG-1:0]    I6a81b4485598387e4656c35e83866209;
reg [MAX_SUM_WDTH_LONG-1:0]    Icf7630b6002db2f9b59d5323d6cc8105;
reg [MAX_SUM_WDTH_LONG-1:0]    I3db0adb3457cb22c755f5d29a8fe7ed8;
reg [MAX_SUM_WDTH_LONG-1:0]    I887911fd9466f4d4fa7f50642d610d88;
reg [MAX_SUM_WDTH_LONG-1:0]    I9ae284c0089ae462a1bb9d168bde2fd0;
reg [MAX_SUM_WDTH_LONG-1:0]    I342a563de39175fe4a6eb7e3e1ccac9a;
reg [MAX_SUM_WDTH_LONG-1:0]    Idc758f8e6fabb6b31b0a7d9c0c590310;
reg [MAX_SUM_WDTH_LONG-1:0]    I72b4ef48363856af7faacc85eafbaf2f;
reg [MAX_SUM_WDTH_LONG-1:0]    I4ae2f2330a8ee7d5626499f2a030c7a5;
reg [MAX_SUM_WDTH_LONG-1:0]    I4aa98503fc71292d42dba1cab6db952f;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic35d5ac4dac46d47b2796bbac6452161;
reg [MAX_SUM_WDTH_LONG-1:0]    I32679702c19eab37b46d13bb372967ea;
reg [MAX_SUM_WDTH_LONG-1:0]    I6a86b03402bd2e35208d3fc74601f9cf;
reg [MAX_SUM_WDTH_LONG-1:0]    If8a259e0c4f1839e852abec6e1b904ee;
reg [MAX_SUM_WDTH_LONG-1:0]    I938dd59e4cdf3434086f60d000113430;
reg [MAX_SUM_WDTH_LONG-1:0]    Idc198bd5732ca5760d1a700a25273ce3;
reg [MAX_SUM_WDTH_LONG-1:0]    I9dfdffbfdb83572cc3205f674e5db753;
reg [MAX_SUM_WDTH_LONG-1:0]    I60520c850a95b893528569c4069bd677;
reg [MAX_SUM_WDTH_LONG-1:0]    If525ac3dc97e3187e036d70e9984939d;
reg [MAX_SUM_WDTH_LONG-1:0]    I0c1e4d400520935c5c78b792a9d554ba;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic7d5fe6c4b1dcb97d10ba3de2f95d1df;
reg [MAX_SUM_WDTH_LONG-1:0]    I8efad9622c05177563ab8a2747879044;
reg [MAX_SUM_WDTH_LONG-1:0]    Ied4ddedaf801fbd7238d8a55c17c8090;
reg [MAX_SUM_WDTH_LONG-1:0]    Ieb9720b6beb2363d651346ef0233cd49;
reg [MAX_SUM_WDTH_LONG-1:0]    I202aa0814e7e28a6bd21db116b652b4d;
reg [MAX_SUM_WDTH_LONG-1:0]    Id201f81bbd80a70006a10866b8efeeff;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic227f42a20219c6638ee3343ca445acf;
reg [MAX_SUM_WDTH_LONG-1:0]    I507e9bd0265d9ca6cd21a46fa21ba084;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie04e44d8e0756cdf34cf9ad53da76e47;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic92ab3dac1a151d6ff0b4e0c21003eb0;
reg [MAX_SUM_WDTH_LONG-1:0]    I3da241c7f221413abfbf1b4384bfca5a;
reg [MAX_SUM_WDTH_LONG-1:0]    I0807a826e91f92ef279ccf0b6512a428;
reg [MAX_SUM_WDTH_LONG-1:0]    I05aabdf73200996b7bea8db700fa8930;
reg [MAX_SUM_WDTH_LONG-1:0]    I03038b940be8bd21bd26b150b28754a6;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibf547f8a5e1059ffaabeb3f447904dcf;
reg [MAX_SUM_WDTH_LONG-1:0]    I2ea27544ba4cc14d0f7ccf7158a27a2f;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib2f34922b0d5346500de093275bebc94;
reg [MAX_SUM_WDTH_LONG-1:0]    Id2e223005a932987b6f60663773187f8;
reg [MAX_SUM_WDTH_LONG-1:0]    I3188d354c2ba494ffe210dcd89c00620;
reg [MAX_SUM_WDTH_LONG-1:0]    I09faa07bf38acd96c4e29afd8a5167e8;
reg [MAX_SUM_WDTH_LONG-1:0]    I6d4867d03d9187e95e27e99f7aecddec;
reg [MAX_SUM_WDTH_LONG-1:0]    Ifb09b84f9681c7bc28ffd562b633ffd9;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib55b0e4c45ebbdb605f0ba9d62bff21c;
reg [MAX_SUM_WDTH_LONG-1:0]    I4319fa23d59f4e690e31fb7e3a823d17;
reg [MAX_SUM_WDTH_LONG-1:0]    I4ee3f608cc8f8df27345949f1a3713a7;
reg [MAX_SUM_WDTH_LONG-1:0]    Iede5d56e52612e083407888da49470e5;
reg [MAX_SUM_WDTH_LONG-1:0]    I3b2739319710681986b9d3f8cd04f619;
reg [MAX_SUM_WDTH_LONG-1:0]    I850c257a0412bd9bd6001817bd9d0ee1;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib7875bf9d30d071e62a474c50d88ba06;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia92b76ee5b7d82a992a1b58147c0c0be;
reg [MAX_SUM_WDTH_LONG-1:0]    I2253b32e46200a23dba243819fce02f0;
reg [MAX_SUM_WDTH_LONG-1:0]    I1b01cadaac7d3d15007f0afe5c0ab0f2;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie96877deef8b1676138f814c4a720800;
reg [MAX_SUM_WDTH_LONG-1:0]    I8ce945d9f70bb317064a8d2d4eafd2d3;
reg [MAX_SUM_WDTH_LONG-1:0]    Iaed105b99eae5b078521e3a94d8a79b7;
reg [MAX_SUM_WDTH_LONG-1:0]    I05a812cd935867d1e417c64c26ea0952;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic0a580f94f3d03f72e3a487f84bf6612;
reg [MAX_SUM_WDTH_LONG-1:0]    I39d9044227c161f0163e58dd82aadc90;
reg [MAX_SUM_WDTH_LONG-1:0]    I5f607bdc9b276fdf07a17a11a20a6720;
reg [MAX_SUM_WDTH_LONG-1:0]    I12e8b8cf609c2fbdc72efce9bb5dabee;
reg [MAX_SUM_WDTH_LONG-1:0]    I6fdccefd034e8b4b86cfa997502512ae;
reg [MAX_SUM_WDTH_LONG-1:0]    Idcd5283cf7b42d403ee0e4404b5b311b;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia020344403aad35e050765a4b0cc42b7;
reg [MAX_SUM_WDTH_LONG-1:0]    Id11fd3a31b70da0e64138e71840cfb83;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie9c5e7c98281cd1deb6acc51590c9d9a;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia0e77e9544481aa0f56dfdb6eb253137;
reg [MAX_SUM_WDTH_LONG-1:0]    Iec0d7ea31e0f1a75b15121090dcf1e11;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia98bb3648ce3719b1c31ce0f41121c63;
reg [MAX_SUM_WDTH_LONG-1:0]    Id9c8055ef530f2cb8096cb7bb2af55a4;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib9081d438413a627f5b16f68c2eabb80;
reg [MAX_SUM_WDTH_LONG-1:0]    I9c5bf5451736358f8c84e150004fa5a9;
reg [MAX_SUM_WDTH_LONG-1:0]    I377933518c3807edb71f648c65ad5c85;
reg [MAX_SUM_WDTH_LONG-1:0]    Icec98d794a64752081fadfa74308fad3;
reg [MAX_SUM_WDTH_LONG-1:0]    I7bbe4d0a7d61d3f7da346de71b9a3a5f;
reg [MAX_SUM_WDTH_LONG-1:0]    I197c05f74bf7fb8d44124d40bd7c6563;
reg [MAX_SUM_WDTH_LONG-1:0]    I92acc55d81ec6e02880337b0a451ae21;
reg [MAX_SUM_WDTH_LONG-1:0]    I35c0ca76b28cd2f9355276b5d2f29ad4;
reg [MAX_SUM_WDTH_LONG-1:0]    I29da0e5661f29bd8493c19885c998582;
reg [MAX_SUM_WDTH_LONG-1:0]    I9426c8c1b4d988d5cd7d89a7aed4f8fc;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibd010f15e36194cbd2ce9f01c98a2b6f;
reg [MAX_SUM_WDTH_LONG-1:0]    I7e86ab53e6d9647b230a94e076831ba2;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia0ecfaedbc1d546d484978fd50096d10;
reg [MAX_SUM_WDTH_LONG-1:0]    I27098cbe2d4fdd634385d771cc290c2b;
reg [MAX_SUM_WDTH_LONG-1:0]    I5d7a0739e447775e00115799c52b11dd;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie95793e09085b6de1383a37cc7fc41ac;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib24b68cb35da39a743e1d90bba3f0836;
reg [MAX_SUM_WDTH_LONG-1:0]    Id4cdd72193e90dddd211af73d7f3634a;
reg [MAX_SUM_WDTH_LONG-1:0]    Iccab4c19a9190689f90a42160e2379de;
reg [MAX_SUM_WDTH_LONG-1:0]    I275ea08a3dc0600d8ccb6300eb7f2a6b;
reg [MAX_SUM_WDTH_LONG-1:0]    I1b53098a7240d2b5dc1f5c5c3b4bcc11;
reg [MAX_SUM_WDTH_LONG-1:0]    I278659ca1a0b093fc883d01987989dc0;
reg [MAX_SUM_WDTH_LONG-1:0]    If92e66cba66732798dd19f968a5ef8ce;
reg [MAX_SUM_WDTH_LONG-1:0]    I784c4e9fb75c314f271477e0621aaf7c;
reg [MAX_SUM_WDTH_LONG-1:0]    I3d3aafdd4d9d3e9fdab1f487c48a0ea9;
reg [MAX_SUM_WDTH_LONG-1:0]    Idb4c722992139f39914af7085378c6cc;
reg [MAX_SUM_WDTH_LONG-1:0]    I63c9deb7e6a4b400e0aff6887a09e647;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie6f67c6e4c5e2b8357c0a902979e8722;
reg [MAX_SUM_WDTH_LONG-1:0]    I1d7a4f99e3975fd01bfe5a9a1da84765;
reg [MAX_SUM_WDTH_LONG-1:0]    I059d847e09f5aa3f6a8147062f4b13bf;
reg [MAX_SUM_WDTH_LONG-1:0]    I48e5256ade4d061a3b5ba08a53252bc3;
reg [MAX_SUM_WDTH_LONG-1:0]    I635fb29c55e0fb5cff0b6f443c2e3de5;
reg [MAX_SUM_WDTH_LONG-1:0]    I088c5b971a2def57248769a33b7d2a2d;
reg [MAX_SUM_WDTH_LONG-1:0]    Ide22394fce1658f9e7002bdb30d03c2f;
reg [MAX_SUM_WDTH_LONG-1:0]    I9ff276a14d3205b98174a8a736f79774;
reg [MAX_SUM_WDTH_LONG-1:0]    I123255637493b9c7924e3a72d1b86ee9;
reg [MAX_SUM_WDTH_LONG-1:0]    I87e6ef84894cfc86b94e19c9d3065bc6;
reg [MAX_SUM_WDTH_LONG-1:0]    I4c32900878260a261bc5403e8abd6258;
reg [MAX_SUM_WDTH_LONG-1:0]    Ifc100357ae3f754fb0e3863334bcc764;
reg [MAX_SUM_WDTH_LONG-1:0]    Iefe9e5376010997c0ee52eeb28e57a25;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie6060acdcb16b6fa6aeeb649ed621053;
reg [MAX_SUM_WDTH_LONG-1:0]    I46c2b923860b0d1c01b9475f4467f280;
reg [MAX_SUM_WDTH_LONG-1:0]    I38b4eceb159ecb0dda3920290a21a02a;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic45561ffe1837c3d5bb42c695a377f82;
reg [MAX_SUM_WDTH_LONG-1:0]    I3e76abc721bf7ed186f4d0f8f4bbf4e3;
reg [MAX_SUM_WDTH_LONG-1:0]    I1afb4061458e9d2f5799afa1f2373bd2;
reg [MAX_SUM_WDTH_LONG-1:0]    I18bb9a781a4c314fe6bd990e4c275f67;
reg [MAX_SUM_WDTH_LONG-1:0]    I49d7342f105c4502377abd23db973752;
reg [MAX_SUM_WDTH_LONG-1:0]    Ieeb12d463444ca36af1ecf2e09504c06;
reg [MAX_SUM_WDTH_LONG-1:0]    I17525df1798fa2c1c4bbc4a1ddcdd0a5;
reg [MAX_SUM_WDTH_LONG-1:0]    I90c44c31fa7903a81826c1c568597362;
reg [MAX_SUM_WDTH_LONG-1:0]    I3997cf122743b612f49cd5dd125a9201;
reg [MAX_SUM_WDTH_LONG-1:0]    I1112c4267582ddb8148ee40d9529beee;
reg [MAX_SUM_WDTH_LONG-1:0]    I21c207af859b94634d3750482b42a2ca;
reg [MAX_SUM_WDTH_LONG-1:0]    I2ff2421bd86bf9ec110724460f1171e9;
reg [MAX_SUM_WDTH_LONG-1:0]    I6ba5c453b17e4b33c61caf5d70041c4a;
reg [MAX_SUM_WDTH_LONG-1:0]    I08318099725fbe033ab8d5427eb8b278;
reg [MAX_SUM_WDTH_LONG-1:0]    If36cb462cdf20b0b1758cd6417e524fa;
reg [MAX_SUM_WDTH_LONG-1:0]    I40e8463645b1122b7cb224770fa00447;
reg [MAX_SUM_WDTH_LONG-1:0]    Ide386e751e06dd5df0c042cd76f0f800;
reg [MAX_SUM_WDTH_LONG-1:0]    If63bb4681bf1116c0d1db3aa21bf52ac;
reg [MAX_SUM_WDTH_LONG-1:0]    I566c72342c69969892480fae41232c37;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia0f7deea6b1ce1050dcf97fa99de9178;
reg [MAX_SUM_WDTH_LONG-1:0]    I992b9876530d53c1b62d98511bf41942;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib8861f627f6273c0a031bf43e7812a5d;
reg [MAX_SUM_WDTH_LONG-1:0]    Ieb5bac4ef0f5e4e0b826cdc43ae71471;
reg [MAX_SUM_WDTH_LONG-1:0]    I3cd0883d9f0ba7475f474f1e318ef023;
reg [MAX_SUM_WDTH_LONG-1:0]    I5f8a41ab83a9257e534973e981e28e9b;
reg [MAX_SUM_WDTH_LONG-1:0]    I0e420136675d5f0d1aa027d589ee8741;
reg [MAX_SUM_WDTH_LONG-1:0]    I4aab6ff52e3fba90bb7417cb50766125;
reg [MAX_SUM_WDTH_LONG-1:0]    I1ba7f209cb735471073e8051026a148c;
reg [MAX_SUM_WDTH_LONG-1:0]    I711c5cf9fd8c5161bac36060b3443503;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie3591b22e0e127f04658da68d4846be9;
reg [MAX_SUM_WDTH_LONG-1:0]    I409129c0bf5d361e9916b6dc98e69a7d;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie4f4faa470f572da2081b63b6df6e392;
reg [MAX_SUM_WDTH_LONG-1:0]    I5011dfbbb0eccfebcff255e4a2c5e64c;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie32ca6b91d1c55883be8f63acca78764;
reg [MAX_SUM_WDTH_LONG-1:0]    I6c7965d39dc839a9df56e628c77a5457;
reg [MAX_SUM_WDTH_LONG-1:0]    Ieac9cea5f36bd82f87105b530e8fb614;
reg [MAX_SUM_WDTH_LONG-1:0]    I79657595561eac53237215fb4110f09d;
reg [MAX_SUM_WDTH_LONG-1:0]    I9b46463a6c54c3668e76190d942b7b38;
reg [MAX_SUM_WDTH_LONG-1:0]    I3ff883ad434cd5153b67186b6b21418d;
reg [MAX_SUM_WDTH_LONG-1:0]    I92abaae6fb89206885616877cca1e25a;
reg [MAX_SUM_WDTH_LONG-1:0]    I33668b0ef7defef974b7a4c0f87689c0;
reg [MAX_SUM_WDTH_LONG-1:0]    I338daeacf82ad288b14c6b5bd4099870;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibe085a39ecb07a8dca62002afa38df93;
reg [MAX_SUM_WDTH_LONG-1:0]    I1f88dddf05f255942e2749891a7733da;
reg [MAX_SUM_WDTH_LONG-1:0]    If1d0be4e9b995ec98c346e8392b9518a;
reg [MAX_SUM_WDTH_LONG-1:0]    I56a4443759b3d786bc9a34a0dc32abf0;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic826d371f2cfc503f5d9e43dc17481e1;
reg [MAX_SUM_WDTH_LONG-1:0]    I5502f383dff392ef1be4cbbf9dbc3c2f;
reg [MAX_SUM_WDTH_LONG-1:0]    I96e6f1dc0cd451da6ac9170d5f83976d;
reg [MAX_SUM_WDTH_LONG-1:0]    I10cd840a369d3e25556a41beede2be27;
reg [MAX_SUM_WDTH_LONG-1:0]    Id85c2285fcc45211f0fa6963b74a663a;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie0bdfac78159144aa65090028931a3bf;
reg [MAX_SUM_WDTH_LONG-1:0]    I28fa30cd1f3b476fa6a354863108cbcf;
reg [MAX_SUM_WDTH_LONG-1:0]    I7a927f4f266cc5253ec30f5c127bb17a;
reg [MAX_SUM_WDTH_LONG-1:0]    I7571c7c306861230de71a75fca79c5dc;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic79811a48840357d0b6303e7b19413dc;
reg [MAX_SUM_WDTH_LONG-1:0]    I0f29300446f020dd23cf847d3e3d3530;
reg [MAX_SUM_WDTH_LONG-1:0]    I802bd5b13c183c37e842f7e9278f35a9;
reg [MAX_SUM_WDTH_LONG-1:0]    I0297905b35f06697625420b7fc2434f7;
reg [MAX_SUM_WDTH_LONG-1:0]    I8487a819dcb61016798cde56f9662fcf;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia2904a5d5db43a209bd4b358ace68c6a;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia8b29ca047a643f47bd3a0ffb50bf8cb;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic45d0537b94bc30713c0a0ee07b1ec40;
reg [MAX_SUM_WDTH_LONG-1:0]    I337231f0dc7eb85f7d950262e0adb724;
reg [MAX_SUM_WDTH_LONG-1:0]    I530cf1f747d1df44b913f49eee90c079;
reg [MAX_SUM_WDTH_LONG-1:0]    Ief52461e4a5ddb128be5e439edf34862;
reg [MAX_SUM_WDTH_LONG-1:0]    I46d86bfa6de26f3cfef9d802549ef2ad;
reg [MAX_SUM_WDTH_LONG-1:0]    If6a3bd6f002d91e0773c4ab9caaaa01e;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib33e1c6d57e5e6fc465dc9c9a7cf29fa;
reg [MAX_SUM_WDTH_LONG-1:0]    Id92a319da408be46970faf524513fdd8;
reg [MAX_SUM_WDTH_LONG-1:0]    Iae182ffae6cea89363f0ccc8b5679561;
reg [MAX_SUM_WDTH_LONG-1:0]    Idfe6aecb694385ce8c3c1544a4992a20;
reg [MAX_SUM_WDTH_LONG-1:0]    Idfbc5726963cfa31bb4324143ffd08c7;
reg [MAX_SUM_WDTH_LONG-1:0]    I205d5fdeae55fae7be2f06f11c949244;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie667e1755ae1561a2eefae9b63845dec;
reg [MAX_SUM_WDTH_LONG-1:0]    If7348fdbe0400aab92e8fd6a7cf6c267;
reg [MAX_SUM_WDTH_LONG-1:0]    I143b91852fddcdcc30bf1041332c4ed7;
reg [MAX_SUM_WDTH_LONG-1:0]    Iee5e74945ba15220f0f707c9c1927ba1;
reg [MAX_SUM_WDTH_LONG-1:0]    I4d1c47569b0bc8c651c897ac8e88bd1f;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib9d6c5be487a434fbafcda25ca9351dc;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib0d033ba28e8c606ed92207049c76884;
reg [MAX_SUM_WDTH_LONG-1:0]    I300d9f403e33d860ff5dde9f91bae11b;
reg [MAX_SUM_WDTH_LONG-1:0]    Iebfe0fa45e4b34e142e82ddaa15243cf;
reg [MAX_SUM_WDTH_LONG-1:0]    Ieb778442bc855e93e11c9b13f1a7ae06;
reg [MAX_SUM_WDTH_LONG-1:0]    I57a393cc9cc9e1abc7962aa2cc840a7c;
reg [MAX_SUM_WDTH_LONG-1:0]    I0ffb8b65525af38861280645ac310e3d;
reg [MAX_SUM_WDTH_LONG-1:0]    I30fb41a57460a0b1f21065b4b97ddd42;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie8298c5c8ff538a3e37af46798f6d753;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie7dc322fee8ca0b6b9659e5183e0d6d6;
reg [MAX_SUM_WDTH_LONG-1:0]    I91bbec0523f77fc52a88ebcc49267e9c;
reg [MAX_SUM_WDTH_LONG-1:0]    I38ae79956762380fadc94f8126dc1c90;
reg [MAX_SUM_WDTH_LONG-1:0]    Id55a1ab9d158ea509e5f57286a3d1b67;
reg [MAX_SUM_WDTH_LONG-1:0]    Ice615e7e18356ae4c3f615dd997be943;
reg [MAX_SUM_WDTH_LONG-1:0]    I57b40c72004f2c3072cbdefbeef72b7c;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie38351e19bdc4f2ce9caf75fc3937dd4;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibba6269b560db9d4913e1e515ed8270d;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie392719059587a201c0148138ba2a2d4;
reg [MAX_SUM_WDTH_LONG-1:0]    I4852d6bacfd82fef6fab4502d61e9a37;
reg [MAX_SUM_WDTH_LONG-1:0]    I9200526d94c38e638370e9a2d7fed75c;
reg [MAX_SUM_WDTH_LONG-1:0]    I15b8aa7d973edcf3b2365040f5570d82;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic3f8e77259ee3eb5be80e11b607818bd;
reg [MAX_SUM_WDTH_LONG-1:0]    Iabf228f57ac154c417389f6711af1950;
reg [MAX_SUM_WDTH_LONG-1:0]    If37de611ce4fa330c4fc9dcb87d4d95c;
reg [MAX_SUM_WDTH_LONG-1:0]    If3c44eb85217da3b6bddb5aed97a9bb7;
reg [MAX_SUM_WDTH_LONG-1:0]    I8c36318c45dabe6bf540381373f09fe5;
reg                           I3931f8f1df3ef8a71a54685fd9eccd76;
reg                           I3c62d5bd891bd3750b7bd1d32612f589;
reg                           I699819696b0299ab80e7233d054ec590;
reg                           Iac11baea9832d6493626d2fe40fd385f;
reg                           I92354deea988f3beb25bfba90735c6ac;
reg                           I6d3acefe6d7dfb94a5d66dcaa1bbbb76;
reg                           Ibd047e2643dc68affb5b4f25b82ded31;
reg                           I65e382d77592c7d1af308d171b27ff3c;
reg                           I7d4dc5e91ba3d952184d90de12f67bd3;

reg                           I86a86d41a29fd0d7596d668e79aca825;

   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
          I3931f8f1df3ef8a71a54685fd9eccd76 <= 1'b0;
          I3c62d5bd891bd3750b7bd1d32612f589 <= 1'b0;
          I699819696b0299ab80e7233d054ec590 <= 1'b0;
          Iac11baea9832d6493626d2fe40fd385f <= 1'b0;
          I92354deea988f3beb25bfba90735c6ac <= 1'b0;
          I6d3acefe6d7dfb94a5d66dcaa1bbbb76 <= 1'b0;
          Ibd047e2643dc68affb5b4f25b82ded31 <= 1'b0;
          I65e382d77592c7d1af308d171b27ff3c <= 1'b0;
          I7d4dc5e91ba3d952184d90de12f67bd3 <= 1'b0;
       end else begin
          I3931f8f1df3ef8a71a54685fd9eccd76 <= start_dec | iter_start_int;
          I3c62d5bd891bd3750b7bd1d32612f589 <= start_dec | iter_start_int;//I3931f8f1df3ef8a71a54685fd9eccd76;
          I699819696b0299ab80e7233d054ec590 <= I3c62d5bd891bd3750b7bd1d32612f589;
          Iac11baea9832d6493626d2fe40fd385f <= I699819696b0299ab80e7233d054ec590;
          I92354deea988f3beb25bfba90735c6ac <= Iac11baea9832d6493626d2fe40fd385f;
          I6d3acefe6d7dfb94a5d66dcaa1bbbb76 <= I92354deea988f3beb25bfba90735c6ac && ~converged_loops_ended ;
          Ibd047e2643dc68affb5b4f25b82ded31 <= I6d3acefe6d7dfb94a5d66dcaa1bbbb76;
          I65e382d77592c7d1af308d171b27ff3c <= Ibd047e2643dc68affb5b4f25b82ded31;
          I7d4dc5e91ba3d952184d90de12f67bd3 <= I65e382d77592c7d1af308d171b27ff3c;
       end
   end

// `include "GF2_LDPC_fgallag_inc_all.sv"
// `include "GF2_LDPC_flogtanh_inc_all.sv"

function reg [MAX_SUM_WDTH_LONG-1:0] I29b4fdd4c13c96461c76660df767ea73 ( input reg [31 :0] I8e6a6a3bcc7726a2e71298c75b3fc8da);
     // `include "GF2_LDPC_flogtanh_inc_inc_all.sv"
      `include "GF2_LDPC_flogtanh_inc.sv"
     flogtanh_sel = I8e6a6a3bcc7726a2e71298c75b3fc8da;
     `include "GF2_LDPC_flogtanh.sv"
     return I0ef7780b478bfb05e8c9bf2fcea00183;
endfunction : I29b4fdd4c13c96461c76660df767ea73

function reg [MAX_SUM_WDTH_LONG-1:0] I2bcab411f9bec1541259751bcb9e0823 ( input reg [31 :0] I8e6a6a3bcc7726a2e71298c75b3fc8da);
     // `include "GF2_LDPC_fgallag_inc_inc_all.sv"
      `include "GF2_LDPC_fgallag_inc.sv"
     fgallag_sel = I8e6a6a3bcc7726a2e71298c75b3fc8da;
     `include "GF2_LDPC_fgallag.sv"
     return I7ffcaba1b7d64b619b19a68a22aa495d;
endfunction : I2bcab411f9bec1541259751bcb9e0823




   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
          Iea07d1adf9016a29cffd61d183e268d0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If92db65b39a83e1c699e4cc6d7f9e57b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8f2986bc015fcc64ac5e5395ac6dd851  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I355725a804e0df68b4acf96ca98f2448  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I78212ae965ab2dcb2eed0b060d6b253f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0b56aa7a1b7549c91dddd3a06ecbaacf  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I71412803cc5229025487255aec62ec4f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I32fcb28a27356bc6f403528836ea4c1f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iad354d876cb9fc72fc0143e6f7da9357  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If6e745bb85abba7282dae1f6f701225e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I93bb43c1b89d4c70a57bdc019d64fd22  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7a2e554d07bbea291f2cfc18694fca3a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3e59b2419c7dd1553b792d536208514e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I46894c6526983bf1ce4b503159131b41  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6404d0df952b5bf8292c753e4c6f35d8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8522c402e654d007abffcb0e904af5e6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5ed85845c39337c37791f16e718069b4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I89013d61c1ea8da8b1c6071cc21c316f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4102100fa5f1dd299af0190862efcc42  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4939f69abb1eac56d5021e06406a93b5  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iadbd245bf842aebb456417579a3e6296  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ifc8ece44a4e68c3117eda9e65f3084d2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I91679dfab57a372eddc7f9b94a231edb  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2213c1a2b831f421707a261f5a58b1b1  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic53b875b2ddcba11406eb2ca39354757  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I634484f00590216c0f74f975c9c83400  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib3b1db2d8b669988c887ed780e439b26  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I735db8b0ee0ec98e4cce0030b11508da  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If1607e907e626902ee26d15020a64c21  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I081b38dbb37d4c14a6a9fd3fefa13daa  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibac5e7b6d4bf5cd6926358318f0c418f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iadfc60386481092ae85cc148a2c40abb  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie0ee5445c56a5f9b41640b57422206de  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie5f8620371236cb11c9e88c16b509ee8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8d7c1fe2e33bbd45379b0325a3c5e989  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4fbdc4ee57a3be42b62d9bd43078d6ef  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5510b88bfd65811b3200adf4ef975b48  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib57ef2f577cca54713c16717cbbd1ce9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I15943aa74e9fbbaebdc0d54eb6a3bffa  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6ac24c46319a787daa5c545de8c6eeea  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I52403a0454e5fa002e79eaab7ea497bd  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I634f0ce28934600a1a31ab0d8e59b4a9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7103aa739616a39c03e675ea0efb0335  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0296d01fd3f9a269a617efd4beea9b8b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I065a81ba25962785215583e7ece27661  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I631a3300cb6685f47da7781940ec5d27  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8bbe1a2ace8f51aa22cca5d9fc66f136  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I38c3e3e136acb79c8a0ff850bcc55f16  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I35b2c7e9cdc53a98913e1c16a3a47b37  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib1a2b31d49ae476e2f1fb9acba2d5af0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic72f41f9bbf470aee3c9b9b8787b31c3  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3ea4c33a9419820ed54460eb64134dff  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia0d940e16c8cbd4f7544f5a5cd7d83b2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4a8abfa0896ce414d9b98093ef84455f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I680be647bf2a62e0ee9b5d379dc87b4f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If4d75f83299a21802b6fbe136913489f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibddfda6413e3dd2f483c3174ea836b6a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I33bddb0adcc2af7b12a83bf843036385  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I529f92b82248efe2cf64f7da0ec8283c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2f34af0036985cd94ade9cc905bec065  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia1a0d8d7dfd6e877f15cce773f85f5b7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5dd29fd1a73df5662d2b636e7285bad9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ide530e6f4622c8a7b101b6dce9650e42  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibaf00a6780325882067a79f0c4d693d2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I16e3559c63ebfed83d6698fc9a9cd93a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9747a02384abb1c2dd1f52b3a5a999cc  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iceb7a1d4c23806b8f5824016779ad129  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I40ef50004a60ae58aedc49eb5e6797c9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I753f92da60980736440aba814a156f1e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4ac79b67a8904b95f7912d24af420585  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iad44c932cfa5c249c5e59f8c706173a8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I10f14b6433498e3b9e9bf021b60115e8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I96008f47b9f134c9c4274cfcfb28e550  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id0344146d1a53d418add6d2b185377dd  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1eede74f12d37331b399eb7136bc621f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3e4754acc31d99bc71525789bdee0c1a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I11c1fc94a3bd6dffa17e1571cc6ae97c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5395ee57418c31e11cf847f0f514ec19  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iff125392fa39afebae1637a19c4e23ec  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia6308e16fae5428f4ab6560f5b21479a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5ea02b5349cd4d99ccbcb6b26f0cfdd7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I21de4f6194dec9e3c401934db92c25e7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I57d0920119f8901bd4dea2d5f8fb5d90  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I89537301987d6da0dbe6cff3caab3ff4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iaf0bbbe791bb71d0f557dc71caa5fb87  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic7ff9cde71054c1ee9eef81eabdd7061  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I88c10c47ae424fbdcb852fbf1e94127c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Icd2e75e47cab1d539ba9ff1b6e1d7155  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I37e6bc7aff363ed0ed1f84b23c5f3e34  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I733605337bf6972630c089d32fd7f98f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Idcb1d8bbdeaed6768c2a418c3048e6ee  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia89da2f1890524ad3519ab403dd0686c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie33a780b0221084898c9fc5b237b244a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iabbd1668e0014df518ede5216232834c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibd89458312687610aa166a9538968851  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Icbaf92a8e9875bcb19a1d074779a9ea5  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I80f3c8559da8e97bc5397bb8b621a0bd  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7a0eada108891aba06cecab5071232c9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie21a2c9b22e7bf8425fb5c0f33e5f4f7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iaa5b2807e5cc2403c5787eeb3d10ca6b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6da2b3a481ee71b85f3087b36b399288  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I11094e852295755925c3c61f1df81643  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9c633aa620cca127b0ff8cf882178e76  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I694d471fd353eb54aae08a2afa7b645a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I816704585ad393f685731104ad3ec64f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I85d95015a9ce27a18ccbf73bbbcdbd70  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I992e7c551b4aa818606c3465d33eb798  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2ead0e9941e2280309ab53535b1e1ac1  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I56873feb8418005b5661c7382f2dbeec  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib6ea4a822da2ea32e0abf6cf8a33d295  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id1659ccdeaea3e59eb2d3f65a65ebd05  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic2171967791a0329f3e39fc19d0a6bc8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7d5041a6796c00188f74936d283defe6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iba7608ee0a01af103e022bcaf564bf6b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iedbe9d0e48bd36064f59faea51afddb9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic3871325d57b310c95ca02fcaca529eb  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I42f9b1f8ef24ad56c10086852678b456  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3ed5d0fca86f35b3d4b4a89c6147d0cd  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib0126fb335e32793c400a97c5a4a337c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I20590d8fb97ec0b2164ffe17826136a7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3c128efc9f80c9b8334bf7b61de71b43  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic7147944f8835e26b9838fdbdc18ca41  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I698b1dbc9d8664d1c86c7a763d97b3b7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I508bbade361787127e1a2e8687ec884c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2afeb2a7b199c0c6738938f156ae4274  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I86255756ddd1f88b74e070b19f8c3bfa  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7d4924388dc5373ad7936dca76797473  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie317e5ea2ca4ba2060d0f491290af96f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I56ea52c50a188ec47e48740839a031c9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id9b9a8fe43992ec0793845715dd2226c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I93b69bfb228db4b569a6772179d603be  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I71afab29cdb962e1f1ca21b61dfb50c6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9905e2686b350e8a6e7f790563a91294  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I524e78ae6a4204e17ba4532dba047d4b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I71228fe4188ab1d9796081184a422094  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie19b39200436b0bfca13502ad36c21b9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If6657f90c84ca5e2ba08ec705f34be03  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I60ec7459bbe99fce295406bee1f2af46  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I29ab844f80c105d247c5c15faa35863c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I856fa68463aa5ef1ae53442699d38b33  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic3d00a27f15f8983a120395082854d6b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6b1d01c3cb8fb51e43cdb788b89816be  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib74a56900c1f8b159ad381f61acee801  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia5eba52d169755c507b9e0094e467fab  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0899e8fec1a7209cd94757c0b2f87c9a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I08ece7cd684e593e02321612b7a88cee  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I691c84d81c60a462e28e2b2bae3ea845  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I58dc9cce6384160c0a85c6efb3319cdb  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I56bf74b5890ec67090f499afdc0a9c88  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibaf2f1f8bda2f6b932dc30f8369c0e1f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id9364a29fd79b52d0442e18dc0227854  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ica3a41ace27f7d94377981079952f4f7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib57795a63d642a73456324bab41384b6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iabf572c97b48c6a7dcc19e56676e3a82  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iefd370d0df1a93639af482f78a1e8706  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I995d2809ffaf0ecda6a004d01cb9c8c4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4e8ebc46bc068c3f9889d970db131112  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7b561638da1b4a45ff59be81243e4471  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If0a3b88a66a816b25f17ced5d0e8f775  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0374ada4fe50717f2158468b7ad205d4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I357137b41bb91e0659b1ac6ead9b5c12  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5d70bc64cf7b3d3ef4180e082e533237  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7d9ad929660cd212387d893266b681da  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I34be4b353cf75603301372840c2f91c2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I14834fc8e6489775359bcecf5a37ff4d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I633a74e4dfa841c9fd13dbb6564c8493  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I157bd468200e63385583b9045758d81e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I918c46173eebc5b2a95e041cfd91d958  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4f8792c18bd07b23e82bbc44b4ca947f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8d0a1ae4c47edf1f2b99d1175aaa7197  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I734e601f5f9d568a44a48834559e04db  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie421da1dc5aaea57c50d0c7d9c5a2717  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ief5cbddfbfb98fce4812a676849b9a98  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id113cab2dd1949d32e3c1c15273185c8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Icfe1a689e33b2b9aa9dba692d6d610b9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia4b671f3360f3ce55db0dc0e4d78ddbe  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I60cbd4369e7ba9b6532f279e5c59084c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ifb6c65a00d9a2c31d8b1119b949828d8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4a777f0dd62b19dd340ad31517c4e789  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib75747cb32130d44b338ed8c8af8ca11  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic7e35cf8d5cd230b94c40714f16e2418  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic51bb9184dfd103703cd0c6ad6edff4b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I103f1449c78c47396d6a54dc1c810934  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I56b3a97dc3037f0bb2eed93a9482c813  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I51e98035b35a35fdc52f5bab8f19c152  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia6a7f9beaceb08d81012f0e72171252f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I21b062856ced09cb9131c01b5e166f32  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4f1221ce7880729fe584b42ef3afe6b2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie7f3f1d6cee7f02ae1b17740ed54c049  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib196f5bcf9152703dc32c5101076600a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ide9ef5a16d8fe32353c2c2a30e8ee3b0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iee6f2484a381bd42e441ff072ec582e4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I53121a39de0bcba91a4d0438be2ae958  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iff7950f24f0a6b0073942c37fff49d37  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ide86f019e9573706c25bd8b4552396a8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2370042234b0e93bb66e44b97fca3e43  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If9efe7a1c359ec03014a52870ac13aec  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6a6eb62960b616043415406ebfc21346  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I06c7728ef64be8311f48d10d766d0c44  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9fe11f6c8147391aa4a5afd1a4e4f731  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id50edc56fce48130247fdbc42eeff9ea  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If3e5161254eb9056914c46263b865c10  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I58703e8b6d04f8c69ac38f5fcfdc4efc  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie1f41720e296ced1b74cb325b666d88f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5d5701435c96f1078e741921b56e3c65  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id96e744d9b10dcddd1ae0115ea57a76a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0c0060fe260afa3cdc72f35ffb6938ff  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iaec1f186cb4a65da21d41e637fc628f7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9c15a6a5c0db11ede80ff6d04c9a56d8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8922487573e02d684a3d71448c3828f5  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I47f17afcd5871fc3ac378316fd3d7ae9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia9642d79bb50567348083b4435c7d66d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2b2bd845428c49346ef8e94e95b618f8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib730fdb59198f23d1e590f6d6039e96a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I644e83f0a7d432fba38ffb2d99088eca  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I97f2b15ce0a74e68d5a4438111adcb0a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I84c88b631bed5311cb6e99e58941149e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I45c5e6710240685bf54b73b0d7a64271  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5827bc87b5db1801b7db16e1e61515db  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1c85c8f73ef80a6808c6aec0c8eca8ab  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id13c99b7f7500c8195b54627efbc4232  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4636821315d702a677dc93113872e647  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9c981b0614a29386ca5e8ebc06a17f15  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4df3d4dac24877b14e6d361bafc1a800  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I913d818403024510c55b65b56a38dd89  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I57015930f5b09a6c6b030ed01dad2177  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib54d55a70605119e37e9898b940ff636  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If7e146da4f3bd255b8457fd6902005f6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ied00d87af99ae55144fdde41ebfc1357  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7774313f1ae5a2de98855aad572b3676  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I679baea452c3c6d04c53baa88edd8eb3  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If4132b39ddb92aa02d8d0346fb0e6691  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iba70e737d52e6812a67c159520e5192f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib9ceb8315f0cd848f861bab677c2c694  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7846bc2cc11e08d05f7c853c4920d555  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0865623d3350645e63fa6e6c9b78ac57  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0262b30a4efa9f1cfb11d1c3940de9e7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7a2e79d42779ad235bca6ce3757cf588  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I09e9a3cd4c12d204f760758e873a177b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I30b0b1d54912c1a41a02a25ab238bb54  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I49fb0909ddf66fc0073e6400f1a07844  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9938397dc94002481984f5b560fadc58  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4378d139db4b710e3587aa72df22b70d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ifa43d74fa91b7b9884969f575ef9ca8e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7c19a79f441ecbb73685db5a505e7479  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If2af8106efc1f7dd02c074af68278b3d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I89a3f8d5f760d1a650f85814cbfdc017  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ifae345c79662c3df3dff0fe68ad68746  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I88a61cf72347d695489909d0819332ab  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9aaa036a6158d11c235bdc8406d79f4c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie8df350430970b5f1229cda772440f85  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7d77ac9b64b2e8cae21c6e36947e3ca2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic1faed76fca5a9ceb7db26c2f43623d9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3ca2b9b77ed8d78a10aff42a07a53b07  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1f00849ea055a7893df386aed162a7b6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iaf8a19fde3de660c3fa925593bebbe0c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Icd1da43a4d95230e79dbd35a7ae41066  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ice9079fb6e08d629f8c0c9ce332c8f11  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I15fafe2baba4d2f28037023a81ce0a81  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If4d5b48882e9e628cf51ad2ac2f38c22  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id0eef1adba01447c14a6f005782dd9a2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1d1a7c5928982c278d068ebd262254da  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6354a0e638340378124e4df7f3d145b8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0236c912c6d684bf4862b725be9d5951  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6f3be51d69b2b64a04e55b8946d5dd56  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Icde3e6dbcf985682041f30903ad95572  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I46ee30b46020d91707689f3468f00e26  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2605f078c1a9006c93855a9a2b0cf6b9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4d226dd2f0bfcdbea6a2e6a6613c1b64  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5c942076b173cf527e1be2ddb8560e84  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic95191bccb18e26c10e56be395ca6b1a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia284f974dd8a526f31eb81ed71a06e94  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Icc93450a007cee4c0a42717ed7600528  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9ec9f389d0489908d497487e44c6edcd  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If8a527cc7f06a9963a80a880d225d34c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I39ff4663007dbc89b403f3b08a69bb6c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9590eb28a81c730b83b92ef7653e71a1  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2ba1acca919bddcc22a41a28d43a4e3e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I62d8efd4227cb3dc88aa08b6585fafc8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I749e987266a20840bb8a4b1a2a2fc5b0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7607af5d98e8070e3d15cee23cdf877e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2e11a697d7f17ac30302eadb500de72d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia0886ce792e062e22d0c224158cdfb7d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6b3cd79aa87235ff174c0299b855dd3d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie4ae993ddb776bdffec843db0def2f5c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3ed2da9b53daac0852a06ad1acfad21b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Idefa29d4d4e2a6e9147f84893520096f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id1fbbe0594dae272856566522633bb3d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8070a3b7d8b1a7ae90c1a2d27aed09aa  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie88285ce2b9c71de02ebd62e8f44ca72  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ica1997c6c569c1d1f45224fbaa4e6b59  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iaf08bcaaeb15bb0c971432f7f8b16d0a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Idcb37cfc357cc088c775409fb9225b51  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic419255414995e7168afb97b051fa64f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iee6da3120d73373627b25ab7c0dedd28  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I56fc99a22960232b305d6e683c66fcc7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0a9a09b0ab43d2a0f1d1d01e13f0333c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibc73d07e0c97a6fcae791e04106cb082  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I224bbdf94ac86c5c376d1db4f4d4e060  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I43f2b69c6b427de3095c44d4166b77cd  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1e50c90010a3df1a8ce1cff811cc7a0c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie1817cbf3a80dae435a5571dfbd2f5ad  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0052d562fb3182890c8828e52d437b11  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1eedecb1d8ff505c75be7787199afada  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7ef544597a185b1de63b4ffc4a1d44c2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iadeedf3870f0b1eae98d0f7dbbeff04a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I70ae07db9b44d530be220f06401d3d3d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7992ea31927b4f0e268462a3b0f18c5d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iadf927d18644a232ad1f1eba7db82934  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2a9c673cdd7ded79e09ada38c0f47e6f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia86740e870d8063f0266b68ad6d7481d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6627bcdbaa8afb115123777abd45435b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I96fe3eb633eff6958ac575b997460bb9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iefdcb71f2903b11f5cb0b8857f7a1727  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2eb90278aaa54b9c8212b3b4af7c3617  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I43493f70f0336453d77caf7f27503daa  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I26a7fe395eb583258c1ac58aaaa3234a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I21668ff77cf75570cae97f575cbcf644  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie48be9e6b6fd63baa104d0a6a4561a1a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I05370777439b01811fe7f750d2f724f4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Icdcd83341f6b5c404f91ec7e97d0550c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibba4e82d1510ddc16eb4ef64893cec02  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ifb00ae47340bc99669c71da34cccc59e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I75a4cf2948bebc58e12bb039ed273ff2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5a9fdec7d7ff99fe33ad6cd8afd9e059  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I47b1695a74e4d27389b97543415dcc67  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ieb38fa62119a5a77c060d6634e051298  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3459d98131faef5a5040a03847890b55  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie9b9221b2122087cd5f309570b6d31ca  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id4451722e8e2393d627dcd0175dc9903  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic10356f9069e3651b9c045c906e63512  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic3a431f39c678b7175ed30fde1fa6424  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib01cfd833a63500e03333f263805db3d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0b7b4c0a8503c751229edfe0237cc903  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iace01234164c8a9f7c98eeb83268745b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iace8b3b3a4c16763132b5aaa6b24212d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I80a89644e278e96b1cd1c4b7f764dc34  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia92d2276a8a23521ad1b88df7c27bc2e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I39bbec42c442d1e8c818f46ad9c096a8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I88f1b5c12759a5efb2d2ded8483c9ed2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iaf4ae293c576af16f5f43a8b86c1aa3d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I68b575fcbc5321d4d26a22bcdbb506f6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Idf600b93ee1018ecf969ed7944b6bc7b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1cd93172cf5996bc870063aa642188a2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4af080cb4e5cc525db95e5f401019e8c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6fc8044eb226a14ff1a786ddc96d2414  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I27fd0073dbcdee599fbe85cf48806efc  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iaee6d725a8b2653eeac6d5acb91f8f36  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4afdeba4fc2a12a6cbe3567a519367fc  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib42816335dd8475dcc78662c4c0786c1  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I343c9efe71164c01e9c7d599e032864a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I108c269ceec4adcff9afeda01101b838  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I761983331fb6e3c6c437b3f1660f0b6b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I70d32affde22f9dcb2d77430fca39069  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic08e85346f61da036a15345a13ac12f0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If5dfdadb3868ed5a495007362f7db648  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia1ee5579358b564de06c08ca418a9bf4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9bb81dda8102b829441be46460eb8900  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8eef6ca0a61a21882ea28b3d63735228  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I438522d92cce6f7010246424746ca255  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I92496f68b44a94565af28a2c28d6fbae  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I66528f43f614f0edb715564eba3c77c1  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8cab9fba615b94fd4bb6934325be8ab8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I92d9fec22d36b1baac8bd78abfc1bbd5  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4eadce87f47df6d8f0e4acd057de5a09  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I73203143fe37933c16fff873c1abf512  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibed2a63af723a7abf96dacf1951e5266  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id667c80003b5541de9f84d3b8709c828  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I02cbb4255db2b21ea32140f9e9ddb36b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I65354f2069de0c25bbe7cd50fbe892aa  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic279867ebf3055980f3d813d5dc8dec6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5c05da8a222ad5effb9815cbf3ec25f3  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib8bf21f32c0e8b9cfa42a53807bfe3a3  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7208256bb198bfce1be71390b01bc028  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I49f2a06ceb3a59773c65b19f54ff362b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I86e495dc894d2aace15c1aff89798bf7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0d53bb5344cabe5fa5ce3ecf7122a260  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib2f5f5fc77ea8b529f2471c54388f2d1  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Idcada1bfb3c0d1f2a09aab58a2071a57  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I814b62120953991f9da055f118967e05  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I123a212546a8ac394051425db4924812  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie95f1a7e0effcec0aa423dc803056a13  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I106deaff50b8480eac31ddbae2ec7c61  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I68528be9951f5b8805411711cd11ea59  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0f034a8f077b0ab231727b6298e366d8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If9c12f8662333fb54a45cfa1bc5da487  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie1681d905517daafcc7584725cd6014c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2ff3edcdb6158f1e3c9a555aeefc0850  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I43b380be6df7df0d354223d0a0d6d6b6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I23eb1dc4d1c992f804dd04a2d823c778  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7f90f96c0260560ad5e6dc7448b2670a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I07b417cdcc99eaea3413f563e26ddc73  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2f3ab9654e515a54e22e73d6c130ccc3  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iebdc41368d57498a04fa73e30b10a966  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5b4305bef5b4350c1d7ae143667afddd  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2795d21d343b83a69146314a2407cfa2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic6386d7d8813731d612e24b715740275  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4c366a57920ff090a98a2cb8b9caa00b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I14cf5d43fc9864820a8a25efcc5c6d86  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I33b99994abbb5ecf8eed4de39033e4f8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7c3291f0250d13ca94802b0b071a95c6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2c926fd9d306e9ae13364e07c4b0395b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib23edc35fa5bbfe0415fcf0861a22d9b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3e0e682047f7cc36142e668828cbff1e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I99fb9030e8361e57818c07511479a9b8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic87c3d7762a18772972552162e1d1a8c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7e393e6c1d1bc44daaab120d55f5dd59  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I448f126fd3932d5065abbe7bb2d92c56  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ifc8c6df8904b97674f2970ebc95b523c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Icd0622a90782b9c451950e7ab0399567  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6493b3c087d4685a6b3f98c73dc2ff49  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I20c2057240417146df144b518b43d052  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ied029d0bdea3bf134744c99426fa72dc  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Icb82c9ff4cb58159a1c3115c6fdd5f8c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia3450e134e4086c35acbdee1e6042396  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5a0f27df5158309f32f0df31e8ae3ae3  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I17d9e19854cef197fd3267618617efc3  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2993acb61f1abe529f8a60c94a438550  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic8be2c94235fb40f78da33179ce4873a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib3367565e4456da15e7c2315dccdb5e4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I15a1671def323cd294591564ae6ef8b1  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic512effb493a06ece58a2af155135004  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2c72248cbe49ec0a0febac2437b8a6dc  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I964e17c41a134c080e9c43412a514f3f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I94f1724740defe5bb7e40041d0e266a0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic19486b6ab0373b9c0ad8f7597782d8f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I31243de90dc2a1656ca9d5e03bdd78da  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I242a30bdc8699d8ff550b25dd53d6c59  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9d15f76bb68b214057566cba4b511214  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9cc16a00912e7dfc05fb505a9db23cd8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iacf9640cbf486411d6ceb8fe1a2fd5c9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9015033ab0caf3fa41dae4de43f24a82  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia630e59cbce82a570ae3890a6c0221e5  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4904ab14b19fa1b6befc218bc7be3842  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I282d2eb4e74e034694e33273b9cb19d5  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3f33901c407a87e10d86c13c83dd52eb  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I43f41bf07836cee48069e9890c1de2a0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id88480a0a350bb5fcf01ed5fff0bbd4c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1d9b9ff357667a362f0442f19986f451  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ice73589836da9028def6efb24a04dbbd  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Idb72c046c5996fbbd80b706666ffbd92  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie5757e7b1647ab7d43cdbcf98cbb77fc  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6072331f838d82329a07a4ffa340c7b6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Idf6875955525d80dc660ce956f4a84e7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia96955d9c0a8a587e0afab37c8415d8c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ifec374bce7f5507438f550df22d61a01  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ief67e897e57b96e2ec200e82bbc7caeb  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ide604e9bbe35cb55892a4602e18b2527  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I262f2390e77ec486ccd3a6ed05816e2d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I280e20c20c0b4f26278b3de9b2ff84e4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib3a0307176d424a4733720416d71069d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I76060709de3ea188748849f043c59ac0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8be20605d26d218911e80a883a90d085  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ieafa9d74d4a61d28ac4a913db460bf33  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6fd1b4395af175eff85b3bfeef4c329b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I39e6d3fb468aa40ea73535e81556ea65  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iae449b74e50e0907feae9e60f2329426  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iebf769a6bdaf214c1006c55c608d4eda  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia030c08757123aae947f86ab8bfb6d94  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8c35c5b343b552c22000e194c517ca12  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibf80bb564263ea85bd886a8617f09bb2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib8dfd9b8badef282ca00a4f793c3c868  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I596ad7e132f272cb196b74faa8c75aa4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Idc629414f6d0236ce0714cfaae23f065  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I157fdf8775206858c08682db3039b084  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iacbb4daf5ce5c7eb1a2afe30d0cb5382  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4e08021c0235fafb60200aab97827a8f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I730634ea15ac94d241f3ad2d6393a227  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iee367c535d9c39f872d2ec043e7e7b33  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I68bb1f26f878862f288c1f57049cf58b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia9b5d9ede006c56a6d83905529c77b7b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1487170cb1f3370ad45efc801cefc8ab  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id88568dd34fbee42c9cb8cc15ac5c31d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia30539545e66c4cfc16828140149180a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Icbfbb37bad6344005dd233b3605a784f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I91a6408a11fab36a8ba3dbd3f895a803  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I47b878f27c30f79a37e97e022307e9e9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie76b0739aec66f8860870e66e87a6445  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I50383e3d7c172eedfa00aa50a9faac4c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ifeaa99e03bda8ded058f98387de3d49d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4255ac1af4367c321567c4e46b06ab25  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia445bdc7def7d8c1eec31ab892c25c41  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic3b4752136ac08e343933ccc3a4ec47c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ica6707efd6d44ba6bbb87c0593a3d828  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I739267bcc50c54b8a685cb3c6afc5cc1  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9160d11439c5140c0109b5190eb82e6b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6ff7b86cd7f63f9243646f1be10b2577  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I165653ab165cfafe2b74cd441331f9e1  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I08a8cd6965c23af6650568b654831b20  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9b6a674dbcbfcf65f1ae0deb8fc3566d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie3a336de822ac7baf8486b1618ef1126  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5fc3c26d6c5aa893dfd5caa0f677233a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie22b94121b58f17af14c75bfb27f96dd  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0d9f8c99194d9d6e187b4ad02fcce8b4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I71e101962e766a4d1484b3235359a4b5  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If2539da6722562bbf31786fd0036666a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I22c8ccd4a9018ad1c129aa058bf579d8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I83330fef69470d2f5def8e6d7d9c50d2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0539d598bbe3d50940329a282c801328  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I202f88fdc946494d55fc8831c2e8a34c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3ee10f6a7785a236db317515fdd23a2d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I453fdf4fbb5af5bd28a20d7643da9eb2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic4a6c02880a9aead7353332708e3f388  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7fb3b66cb48521f8715f66bf5642cdb2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2fd872df07f50688486c0d602cfc5549  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iccefa45795486757515d95e5908b306a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib1357cb20f471f1670ac2448f964f8eb  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iab953a8974a1eb619dc0f074c003b5f9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6e37582849c2c98fd15ad92d22c222da  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If004de0cac6e5f7701a1fce48c6936d5  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic1efa395cc1fd2c5a1d1559fb169a5a0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8e96c69e7d872be23229353808c34953  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib6aded6c73a8cc3cb964b0ae895b859e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I939368b76d98b43826c68c7f468a5632  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I544f6263f16cd5e0b7cf28c511a8f6e3  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I484545c4d2c869d79eb17f51e11070a3  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I39289e6385a9bc378a9b8dd440249a7f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie9cce5746a83479a567bbaeac6dbf497  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic044d7419cc43736d278c2df33b4a3cc  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6714551e8885ef5e4490673fe1b2dad1  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie9ab3c88ac62369e3d92d110165a94a8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If38feb4f76f761dce6145731ad235d7f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6359856a1843d8c8b65dc478bccb3acd  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If6f3d91c3c7a43622b9a522492cd83d3  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id023a6298e65da1f4da3831f5136afc2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6b24690f394792edb0d82b3b9e110851  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5b55c285f7e3e78447fee68532ab9f7f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I32701d9e4b96853c53f0ab651a6a4ba2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I82f266e5792cdb6e7ebd264e246161f5  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibfacfe5b83819afe7fbd4bffa2d6d4e2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib8e68a77ad8b9e7cf415bee17645c3f9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I644ee0055a55f54ab3544bb532e39c61  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic5467e42aa377c6ffd8f70673808774f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic57eb4a034247a4c952d8224ea9f2bac  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia642db613c0ec1ca4e69afde7a14a839  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I432aa7cb844286c442356954f8814260  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If520c1cd27f9d4bc52d0d029f693b660  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie87075ac979410cc11099a356966b8a2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6fab46b1766878b26b53f352fee98223  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ieaf14683f40374c4531326d228cb43c3  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5149125aaaad943d891df6a3c2be93a0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I770dff588ee1f52f58bea1921cb23383  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8f0a90e761111a613d2488285534a500  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I765a8825e42180a6c63f7b33703bb483  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I512cc8f6519aa08aee18225b56d47c9f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If08370fd0e8af818c6db20f43e74034d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0ff382edfc8051459657ffa3899f5f73  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9d2864024148337277523ef7fa2e1600  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1c85a2d1df6749a194072eb731506bfe  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3e3ce8b4ead150a6eae2e5c701c7b598  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I45bc13ae0e0554a79c62cd9c6aa8f2a5  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I92678f5b52c9c55556ff7f17f0f607b7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib4bdc9069d0c08655f5e87f705943eda  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Idbf9094c94c931f16fba468b9dd59a25  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1c3c4ce44610e04c5eef2fcbc2ea5114  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie84be0ae8311d906eff08f7f5b214943  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic90b98708faa8c8b75d4bd9a52c292f7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8eba6f14f42701d22859fbea94bd1871  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6d83efa9f988328f487e9232bf2633a2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic23e01562c8a753fd70c343297be288a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5669856f88f5e2c98f64df696db76414  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic3a608b850709286ea0ad2f67425d9ac  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5267fa34449e6eebe891017fc32d0749  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I599d01cfe6e54d8e45d64446c446818d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8f94dbafaac589ac9f14b56d4556ff96  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I754563caea429d3d0e22df5d193b84eb  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If7f373506cac70f8ba1222db135c27e8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I69f563e7b7ad483893ac9c4684349769  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia0a02781c674fe5d769206448d475245  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1b7a401bc11741e6f011fb9895b5c797  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ieb528d666fdb708279184bb59eac25d9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic3ff7ce12c836bf0693252b9a7a7cfe8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I19bba6a58ad3ef959b33701f82761984  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8acc93b34974c1e708b0e1591f7b2d3d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib60d4ac0fcadcdfce5a14fb92f58423f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I039f05d5be891a37e04556f1eae674d2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id0f75e19b94541ed5c5c352d13390d2d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ife1190f76c2e251704c2960c23330a48  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id3e0c98bff2636e216b4d3a0ffd51054  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If4d3b31b87c0f723241d35ce7e854eba  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I72369dedfe36cb22269033cc305b730c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iec71fe7fcebccf1ae0d10a5d187fcc44  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie11da10808c4ca84f399535df6261307  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I280fa9d114e227cd649bf0e55e845651  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I94c4e11670b4233fa072517a8f19c901  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4dca2dd40a7127ce44f83b430a34c738  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1a24e98165afa62bd14986911a36fb6e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ife1164cad7cda4aa9a08d94dfe86add6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8d8d95ff26f33f69a182b32ccde23905  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2508854bcbab37bd09c9465c377c06aa  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I140078292f7209eccacd53a8bab18016  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I141fb1cbe09f9abe282cffd4de815d25  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If79d1d378f7c6fd29fc3335ec5f5c51d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4a41999cea9357a85c73a0af509eeac9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8e517c401d62dbb10dcc96ab536f6afb  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8ad3627f171eadcc960a688ac0afcbc0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I85c4d3d6c8408c6f38741257ed177ca6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id66c47fd69c175a4393e975a269cf053  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I37dca40506d61bdeab1255ed4892ca20  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I340c98b886123c541a1b8d9fc8a6d48c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2dc64c3b06588542b027f997437bee63  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id92a37c091100e9df08e24498ecb4022  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I74a4b9365391fd20c34588002ad40547  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I461195b7ae78743e09ee50486ad6ebe5  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I356d747600182675699a2d2634d4c5ce  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I87d6a5d30c3e4202cf51f33c7a770c51  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I960768a84aec9d5b8bc7c1c523024a25  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I09b5273bb15d48a7fd78559930fa6d1c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5814a85c45fd0f7be21ed325235fe4b7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib06b60cf9933dd8952206c5f3ccced8e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I67347c413b5efd8ff9e0d5bc7ab2a047  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I72b1bb104bf2843f161448baf7aab44b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib23d889edb5a6d9f27de977d3b1a2616  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ifaff9dd032cf96487be819c59b03000a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I028ce03be0618b816e0ecdf43d4cd6e6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6ae2523095237282533e0b5f1c26b488  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5aba6218461e8d571be03a3ef041ebaa  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6ca8a1fa2c72b1c61d11dc7d1ba5f37b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3ec5819176ad4b0895a9118d90ab22b5  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I49b64469d298012dbb131d879bff38d6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I95361d5f524ccb9feb42811af5c482e2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9c4b34b5fb1d59c132bcaeb6258675df  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I613d4b1e3b9e812b785c9cf14fefdfe6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I848ed394bd4f0b199d11c0ff458394a7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie65a0634454381e24bb3223a333e3ad0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iad166146f7df5e8068fc6efe4d3e4141  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I63e45abd4d27219bddcef06108b72021  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id1bacd13718f7c29c26b63c239d04dd8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia3104c69fb4f7abfb5efa3874169a7ad  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie1b7257c99831ec5864f65958ecf14fb  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4accbad1b451ed2b622e15ef9ae16d13  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5ce8b2f633011e89356243a1a71edeb6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3e5139f24e3d082eb31b0e61ea9fa1aa  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I61cc8a0f49e393721a62a776e4793deb  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie631e40caade823a196370fc3358f042  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4c971e714427664c59c6371e14781bae  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I36ca732e811d67cd742d24fd4cae887b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I354fdd241d5d07f0d8380fe8924e0a8c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id38b705f5d2863a020a475ffffc8afd6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id6e5d67e7bb7c4b999459374ea80459a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I05341013abd4206eb66fcddfd63bfe26  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I15da71a21f5842cb65b543d9bc3e267b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iccf255fb3422c558465e45226068a16d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1c2674b2e6b269ed539827412c5199a5  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6a3f405bb4a0c4448d9b9d3dd95d036c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib528bb7a64cce4f694081d151fa6fa86  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iaa40bd3abf668a21e0f87c7bda7b3f69  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I919d36a7f6ad42c4bbc23222beb73106  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I648d2a279dd1f587b1e45eeb35f2fa90  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I194a64bef92ecf6714141eaa5d41c9d4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id332e7f482524adeac7f7cdafcf5ca46  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I226383d68f89db716cfd8d08b837865a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2bdf5d319ba9089a4da34b108f5c5ae5  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia91800792941ec7cc60415c3f844e4ed  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id7c507d96098ee7a955af8a48ee5d72a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie15e4c1bcdb0e18085d4b320ac6a925c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5485d9edcafc6202f6e5f0969979802f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7fe364f9f537cbef782e7007848a1c10  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I52dcf5bace9cadcf8a895aaa6a8c1da8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I13a9eec6175e695ab8bc4516cf57d6ec  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iee73a7c685a4cee03f33d3ef379b1c8a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I740dc91716e3906ad078e2c7cc3c925a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I514d2dc697e9b39ba027c418a6df6cb9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I782726e317a2aada9e755bcbc4b0d3fa  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I11eb26cf0f0b3a334e8f7317bf8d9eb0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I26cb63ba20245b2c332b09e25c4409aa  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Idd7691d31f8d0c09ee988116d574ec59  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iecc02842a2d2b9b9e8187f2d39e62e05  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5551342f1751fc64f32744a46b9649be  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iff7c29299f005c1cd5a16b64601e727e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I17a5446e942bcc1dc2c96930e0a87a70  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I719b67f84e07e90dfd29a8cd5d94cf39  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2c835dfb3596b8bf057a7cc21122c81f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib71b3d357c98dcdfae5c777ca3082275  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I086bf19f620c8a8f6888e775cb1ed7f4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I802c554d5b04af6b949677819a4966ed  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iceefb06cb3715e1b41e6f7d89420e5ba  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I56948bc48c0220893d68004615a6ebaa  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iec1368f034655d61354ab5b5e94d7d89  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1e43c0aeeb8a2461d208eba24967af30  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia6eb85b127cf9c1a437611556296b967  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ieba89aa901e61218074af53a2484a74b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8b3b875c6c07bd97ba598a5139156fa4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7b33ddad346077928620344542b9481e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I11d967a5c5d14c88b5587d4cfed1d05f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I27458d76b3ac6520fb379405c6b2956f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2525111a2fb5f10d64bbd16e148653b8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7b7cbcd1c6d2a2eeaaff474536a69eed  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id2a7f0781d18dccc7c4e0b383b7cddfa  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If8bc141d98ebe1be7fa81cde5c65868e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8645e1326c66f5efef4b9c923599d1a3  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0426ef66185128dd1ef4dbb68dcda585  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iddd954df5bae9b4240e0512f746669a9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I29e940970d87e8e09b26ab1b0b8f2286  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I488f6d9676aa85a55d030bf12e8997a7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I99d761b75ade1fb2e8afbb1a77752609  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iac4e3d20178049f9c59abf374752dccc  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I618d33f26badabfa578908903a613bce  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I822d7973afe090b2764335f1b72dfd0e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I12c1035353e553b3b6a13bb174ce6020  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia6d61947d36fc128c689808c82db80f6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie9b042f686381739b9ff219041f1e0ce  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0c4268c01aed70ce4fc71531bf4bb862  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia34e42f8de91fa4861b0c6cac5dcfc29  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib7c5850b4f7cc77be2048d114a2128d9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I32bb50faa2b246b2d3b462a79be597c5  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Idc6d40a49f05c5422758cee50f787eb1  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ide1d7dc22a4b271ef764df14ac22366a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7ace6778ac86b3e05939a3fcc716136f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I044e01e8d2df46e03f00a0af2beb0bf5  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I45a7ddcda2662e36b7617dfe64514346  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Idada779a1ac7b844867571d77054b657  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ieeba01b18a244ab8c0ac263c138fabcc  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie4c9797a955778694dd8615219cb51e7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I28a5ed4c239e64c76bb6e566b50cfd23  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I79a705ee1e414fe4a5fb14e9b3ce9597  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I04f90a907f10a7fa1ae3591b48094d5c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I31d25b1b49e65216e90b39aa27acd6be  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1f6540c5f037d861dee2c0091cba01ec  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9632bb500b7faaaaeb649d74c21cbe8c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Idd0217a35c3adc8abc7bb581a5df7a2d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic05b46168884322644db4e331d37d759  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I53c88dc237bb2cd02d50fd7f0a168a48  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7450d4ab3ef0227e93a02bfd620d047b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2b16e5b4e279bb29c3c675b72083e5fe  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I70c92e8ada46476d15ef4b3c620d2601  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib193b07804d6d5f111b06bda487bfa5f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I885433b0ab16c6d87abe45af13c9e529  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I198c055930cb89d0390c336eda8fed4f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I688a2c72e69b217d2673e8da75146a83  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3b6fde4ed14cd68af1468ae1d4cc1a22  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5d3df1e7563630311f56143ee6d97a8e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I90a7ea789d3bf7f9126c786474a56da0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5029424c9d9fe923eeb858b1e62cd758  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1e805c70d50c2765b4a03ad2982dc421  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iba58175a7fd5c5da650222193caff0b3  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7401a0501ba69c5559fbf00c77e58dc5  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Idd9f7ea657ea9cdcb45a7e4b573b9d50  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I53f275395dd6be17961a5edc3e8da7f2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Icab010d78cd66b02e089c74f04bf4e75  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I376a48b7e0195a5aacc76a0ad8bd14b2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I241622b0367dde514f96ece55c8c3964  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If94a1abfb972f63629d07e64dc23863c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I07b9b1f4fa01b16cc69356057d3b6154  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2288a6ad3b748b716249f4adc42d52c4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I022df337bcc05ac5648b8ae2e42f3a76  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I60d9a7f95fb8623753002ecaf9a4efcc  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I23a74ea5e7174d95e6d16a5e85ac236b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie697d28d757df82b3901564bda43251c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8572aedc94f7243ce5eacb332c81eae2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6734123aaf6320da75638b212812732f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7f6dc6f0f403c58f9aaaa70c2383a666  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I66391978843c39b6acbdb4847a01050a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4f756e4125c8af5c412944b273e01cb0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id2c9f7ac95de07148c54803f69347f56  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5061e13a179d27e1ba5f89ce8ee0fd4a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0f7c32fc1548fb49b8041f55c157498a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I89ffab735ee30423c82e079ed98216c5  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9494921d8487ee0b314f75cf0380fd2f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If2b3e7d1541cbd8ffc2b4cfc3ad13a57  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Idf3d79da44f2d686f5bd43c3c1427430  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If8125ad3c9e7f0a2b84106064d320996  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic9018b88fa91fb638bbab0613795ae13  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iad4ea0196eb32f9a152c9e6fe5059e46  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia8ff29ed728e7f2ae4213f00328b495d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I70717726200ec02929f679ef05496455  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iaf1e4c7dae6ad89567836877c08f57d2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Icd09aa81e9b43528af73e23b2f0f80cb  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6ebb2b94f0f80425f8401ae823d92a1d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4a2c3204a6a9936d4a215b46c0ffd045  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib02c0694762c4815448b2c8d3df767c2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I98cee6efbbe565d3a4de16703189782f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibf981c01a9d44cbea3c6d8ead92bc2ab  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I864c33e8ea204d20a9baef4584f22d4e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6ad3228e0e2e1f19648d73e83ba5a229  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie099210a99a4899c53baf39559592690  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ieeec71d9df4613555fade2ced7b3baf1  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4931884e3544af182bcda9061091a42d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib3fb10da528d450251764a9b9ede0dba  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Icdc9e676957b2223d60c413331fa982f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I381f6051282c062ccf53866830344cd4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Icfc21935c007fbbceb2a67ebe1a68a0b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I120d597a80158374726e064fb0f099fb  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2520aa556aadf851f58f0b1820498730  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6203f49a08107f7185ebadeecf2c16b0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia706fb593b63cebbee0321c154cb859b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia4b5f2b07556629673fc6576bc49a5dc  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic532c6b85b156f821e0742f47239a65c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
       end else begin
            // Id66554a95b5375bec1ec7c8e6bbfea7d and I8fee031b61092657fa6474c0ef478763 I55f195813a158d82e2934cfac569575d I12de3a4dab98ef8a7d67aace8150b540 Ied2b5c0139cec8ad2873829dc1117d50 I51037a4a37730f52c8732586d3aaa316 I05531b19bb846b18c09f979eeb429ad3
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib0973b6e90e7678addcb064fded7ce0f != Ibc0871b3c992fd278815fdbefcd2bac0[0] ) begin
                    I91679dfab57a372eddc7f9b94a231edb  <=  ~Ifeb14203f4daf31c7701a6a742be57cc + 1;
                end else begin
                    I91679dfab57a372eddc7f9b94a231edb  <= Ifeb14203f4daf31c7701a6a742be57cc ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib0973b6e90e7678addcb064fded7ce0f != Ibeb5edab51cd6aedad9c2ecedaded6f5[0] ) begin
                    Ic2171967791a0329f3e39fc19d0a6bc8  <=  ~Ib581c19864deecf01268595049268b19 + 1;
                end else begin
                    Ic2171967791a0329f3e39fc19d0a6bc8  <= Ib581c19864deecf01268595049268b19 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib0973b6e90e7678addcb064fded7ce0f != Ib0bf69cc797f330fb2546eb46d2d6f76[0] ) begin
                    Ic7e35cf8d5cd230b94c40714f16e2418  <=  ~I661d84af541e30828bcbd962d72baba3 + 1;
                end else begin
                    Ic7e35cf8d5cd230b94c40714f16e2418  <= I661d84af541e30828bcbd962d72baba3 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib0973b6e90e7678addcb064fded7ce0f != I5686b595177e07dd5bf231a35ee41659[0] ) begin
                    I679baea452c3c6d04c53baa88edd8eb3  <=  ~I1c6928cccb4bf7ea7dfd74e425b9624d + 1;
                end else begin
                    I679baea452c3c6d04c53baa88edd8eb3  <= I1c6928cccb4bf7ea7dfd74e425b9624d ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib0973b6e90e7678addcb064fded7ce0f != I33a6ffad80ddf99a4d316a049078244d[0] ) begin
                    I75a4cf2948bebc58e12bb039ed273ff2  <=  ~I6eabc5c074fb1e2183a5f1ecee87a518 + 1;
                end else begin
                    I75a4cf2948bebc58e12bb039ed273ff2  <= I6eabc5c074fb1e2183a5f1ecee87a518 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib0973b6e90e7678addcb064fded7ce0f != I72a2f42b727a0503d43332c0f22d5ae3[0] ) begin
                    I9d15f76bb68b214057566cba4b511214  <=  ~I0107769bbd7c239685b4818731334437 + 1;
                end else begin
                    I9d15f76bb68b214057566cba4b511214  <= I0107769bbd7c239685b4818731334437 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib0973b6e90e7678addcb064fded7ce0f != Ic2580cbeec8c11a19bd1e2ebc29d255e[0] ) begin
                    I8be20605d26d218911e80a883a90d085  <=  ~If723180430080198d18a08d6775ab208 + 1;
                end else begin
                    I8be20605d26d218911e80a883a90d085  <= If723180430080198d18a08d6775ab208 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib0973b6e90e7678addcb064fded7ce0f != I6f5c991e5fdcf56d582c6f80eb6731df[0] ) begin
                    I08a8cd6965c23af6650568b654831b20  <=  ~I44abc734d6acf92a8e8209186d7a1676 + 1;
                end else begin
                    I08a8cd6965c23af6650568b654831b20  <= I44abc734d6acf92a8e8209186d7a1676 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iee06707670e19a82d911c1750bcfc811 != I8695e1e94cbfcbe4b9eae315b042529e[0] ) begin
                    I065a81ba25962785215583e7ece27661  <=  ~I72aa55988d58c664f3291b5786fc8ceb + 1;
                end else begin
                    I065a81ba25962785215583e7ece27661  <= I72aa55988d58c664f3291b5786fc8ceb ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iee06707670e19a82d911c1750bcfc811 != Iceb64ab2ff8a2e0dfdb74803811d4cfe[0] ) begin
                    I71228fe4188ab1d9796081184a422094  <=  ~Ie69528583db8155917ab3d32a446de04 + 1;
                end else begin
                    I71228fe4188ab1d9796081184a422094  <= Ie69528583db8155917ab3d32a446de04 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iee06707670e19a82d911c1750bcfc811 != Iec7404bc79c58d4d2538fcdf659e9134[0] ) begin
                    Ide9ef5a16d8fe32353c2c2a30e8ee3b0  <=  ~Ib22b47d95b72871e74069fe80a191680 + 1;
                end else begin
                    Ide9ef5a16d8fe32353c2c2a30e8ee3b0  <= Ib22b47d95b72871e74069fe80a191680 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iee06707670e19a82d911c1750bcfc811 != I9c0b88a0be66d62f8ab061aeaee7e60f[0] ) begin
                    I0865623d3350645e63fa6e6c9b78ac57  <=  ~Id9451e945bd26b8dcb4cb83ab4ade73b + 1;
                end else begin
                    I0865623d3350645e63fa6e6c9b78ac57  <= Id9451e945bd26b8dcb4cb83ab4ade73b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iee06707670e19a82d911c1750bcfc811 != I980165c1147ac5ff86619c841c6031dc[0] ) begin
                    Ic10356f9069e3651b9c045c906e63512  <=  ~Iba4627d3d3ef91f168068ed128c04113 + 1;
                end else begin
                    Ic10356f9069e3651b9c045c906e63512  <= Iba4627d3d3ef91f168068ed128c04113 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iee06707670e19a82d911c1750bcfc811 != I8b8b9c4777e6df3eb2b9313e69ef2c8c[0] ) begin
                    I43f41bf07836cee48069e9890c1de2a0  <=  ~I39bef4d462b0a3f88ce1485a58d66da0 + 1;
                end else begin
                    I43f41bf07836cee48069e9890c1de2a0  <= I39bef4d462b0a3f88ce1485a58d66da0 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iee06707670e19a82d911c1750bcfc811 != If79ed5ee2b8710da0608c1e245d07d55[0] ) begin
                    Ib8dfd9b8badef282ca00a4f793c3c868  <=  ~Ib95e457d5ae9fc89e197c249414abbcd + 1;
                end else begin
                    Ib8dfd9b8badef282ca00a4f793c3c868  <= Ib95e457d5ae9fc89e197c249414abbcd ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iee06707670e19a82d911c1750bcfc811 != Ia5cc3055ba3365e64cf59c4d4fd3f093[0] ) begin
                    I2fd872df07f50688486c0d602cfc5549  <=  ~I2be28be47a38e9ca9d3b9167327d3d59 + 1;
                end else begin
                    I2fd872df07f50688486c0d602cfc5549  <= I2be28be47a38e9ca9d3b9167327d3d59 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Id8d5df9e869aaeb107a41a6bca3b89bd != Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[0] ) begin
                    Iceb7a1d4c23806b8f5824016779ad129  <=  ~I2ee6154b613d0d86c2354604e93a9a57 + 1;
                end else begin
                    Iceb7a1d4c23806b8f5824016779ad129  <= I2ee6154b613d0d86c2354604e93a9a57 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Id8d5df9e869aaeb107a41a6bca3b89bd != I5b7caaeb34c43e66e8d095a859e708fe[0] ) begin
                    I7b561638da1b4a45ff59be81243e4471  <=  ~Ia7479d4940b575cf918cb8421f041e44 + 1;
                end else begin
                    I7b561638da1b4a45ff59be81243e4471  <= Ia7479d4940b575cf918cb8421f041e44 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Id8d5df9e869aaeb107a41a6bca3b89bd != Ie1cd04c7668d3f450c387a6c1ad778c7[0] ) begin
                    Id50edc56fce48130247fdbc42eeff9ea  <=  ~I3c5b1cddd608ad869e0182ad68bd0494 + 1;
                end else begin
                    Id50edc56fce48130247fdbc42eeff9ea  <= I3c5b1cddd608ad869e0182ad68bd0494 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Id8d5df9e869aaeb107a41a6bca3b89bd != Id88b9265ff08e0730e6a41abe1f80a32[0] ) begin
                    Id13c99b7f7500c8195b54627efbc4232  <=  ~Ic4425ae997c479e05e12347a803213dd + 1;
                end else begin
                    Id13c99b7f7500c8195b54627efbc4232  <= Ic4425ae997c479e05e12347a803213dd ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Id8d5df9e869aaeb107a41a6bca3b89bd != I19df055705f322292a3601fa63f0e5f9[0] ) begin
                    Ia92d2276a8a23521ad1b88df7c27bc2e  <=  ~I3a0518d0d382758ae579acd7e6cd634a + 1;
                end else begin
                    Ia92d2276a8a23521ad1b88df7c27bc2e  <= I3a0518d0d382758ae579acd7e6cd634a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Id8d5df9e869aaeb107a41a6bca3b89bd != I4a16e8e7946d9a8220304fc1be3fb362[0] ) begin
                    Ia96955d9c0a8a587e0afab37c8415d8c  <=  ~Ifd28c1cd286b7a483891bdd094b70db1 + 1;
                end else begin
                    Ia96955d9c0a8a587e0afab37c8415d8c  <= Ifd28c1cd286b7a483891bdd094b70db1 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Id8d5df9e869aaeb107a41a6bca3b89bd != I9497bbb4f746969a95cff948a3ee9ade[0] ) begin
                    Ia9b5d9ede006c56a6d83905529c77b7b  <=  ~Iadf7734be049c645819d9d023b58c4dc + 1;
                end else begin
                    Ia9b5d9ede006c56a6d83905529c77b7b  <= Iadf7734be049c645819d9d023b58c4dc ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Id8d5df9e869aaeb107a41a6bca3b89bd != Iea7da1f43ba202d753b0edb0be8b3fcf[0] ) begin
                    Ie9ab3c88ac62369e3d92d110165a94a8  <=  ~I5f23af0d0853ea6de084ccf77702b78d + 1;
                end else begin
                    Ie9ab3c88ac62369e3d92d110165a94a8  <= I5f23af0d0853ea6de084ccf77702b78d ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I507f8602a99a1096e4c293ba3c235bbb != Ib58043c04b5c4c86c1c67e57cc66dcf7[0] ) begin
                    Iea07d1adf9016a29cffd61d183e268d0  <=  ~Ic5c99c42e9ebe5dded369ac78a1bedb5 + 1;
                end else begin
                    Iea07d1adf9016a29cffd61d183e268d0  <= Ic5c99c42e9ebe5dded369ac78a1bedb5 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I507f8602a99a1096e4c293ba3c235bbb != I61f0c04673dfb262ef6912eb2df39120[0] ) begin
                    I37e6bc7aff363ed0ed1f84b23c5f3e34  <=  ~I4f2498bec0e96802b82f0419d97c527f + 1;
                end else begin
                    I37e6bc7aff363ed0ed1f84b23c5f3e34  <= I4f2498bec0e96802b82f0419d97c527f ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I507f8602a99a1096e4c293ba3c235bbb != If511a6ea6aa5cda5353658d8e192791f[0] ) begin
                    I47f17afcd5871fc3ac378316fd3d7ae9  <=  ~Icaf86e0abee612aa972388c0b6f90763 + 1;
                end else begin
                    I47f17afcd5871fc3ac378316fd3d7ae9  <= Icaf86e0abee612aa972388c0b6f90763 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I507f8602a99a1096e4c293ba3c235bbb != I6330943c9295298c53e889d47c7904d9[0] ) begin
                    I57015930f5b09a6c6b030ed01dad2177  <=  ~I478c4f13c05651605a2045bb5fd6b60d + 1;
                end else begin
                    I57015930f5b09a6c6b030ed01dad2177  <= I478c4f13c05651605a2045bb5fd6b60d ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I507f8602a99a1096e4c293ba3c235bbb != I3d50cfeaa4b69c09bb648b8873a6bc24[0] ) begin
                    I26a7fe395eb583258c1ac58aaaa3234a  <=  ~Ide67911b52687d67ef0c25f2aadf14c5 + 1;
                end else begin
                    I26a7fe395eb583258c1ac58aaaa3234a  <= Ide67911b52687d67ef0c25f2aadf14c5 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I507f8602a99a1096e4c293ba3c235bbb != I07930a807994815de45864af579902c4[0] ) begin
                    I15a1671def323cd294591564ae6ef8b1  <=  ~Ie9e7630af25f39a0e820181918edd029 + 1;
                end else begin
                    I15a1671def323cd294591564ae6ef8b1  <= Ie9e7630af25f39a0e820181918edd029 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I507f8602a99a1096e4c293ba3c235bbb != I651d700a00d7004d8728bc7356f30926[0] ) begin
                    Ifeaa99e03bda8ded058f98387de3d49d  <=  ~I0e1f07f30cfe36f189e9dcb4e713b5c8 + 1;
                end else begin
                    Ifeaa99e03bda8ded058f98387de3d49d  <= I0e1f07f30cfe36f189e9dcb4e713b5c8 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I507f8602a99a1096e4c293ba3c235bbb != I872f61d20baf011e867b44dc5539fc37[0] ) begin
                    If520c1cd27f9d4bc52d0d029f693b660  <=  ~I31cee5e2a93635987776b0ea477e6211 + 1;
                end else begin
                    If520c1cd27f9d4bc52d0d029f693b660  <= I31cee5e2a93635987776b0ea477e6211 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ibdf2178bd18783c4797c21e642388d16 != Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[1] ) begin
                    I40ef50004a60ae58aedc49eb5e6797c9  <=  ~I84721f2bc5ae10db78d2e7e07cc28d94 + 1;
                end else begin
                    I40ef50004a60ae58aedc49eb5e6797c9  <= I84721f2bc5ae10db78d2e7e07cc28d94 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ibdf2178bd18783c4797c21e642388d16 != I5686b595177e07dd5bf231a35ee41659[1] ) begin
                    If4132b39ddb92aa02d8d0346fb0e6691  <=  ~I6c6d057e910da53aa47441566f95153e + 1;
                end else begin
                    If4132b39ddb92aa02d8d0346fb0e6691  <= I6c6d057e910da53aa47441566f95153e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ibdf2178bd18783c4797c21e642388d16 != Ic2941d16ae6a5cbce70e8546a18ca4ff[0] ) begin
                    If2af8106efc1f7dd02c074af68278b3d  <=  ~Iecbf70768fbaaab8da98eaa9a2b956ee + 1;
                end else begin
                    If2af8106efc1f7dd02c074af68278b3d  <= Iecbf70768fbaaab8da98eaa9a2b956ee ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ibdf2178bd18783c4797c21e642388d16 != I480a0f6d6c3eb936de10a72749f6cd3f[0] ) begin
                    If8a527cc7f06a9963a80a880d225d34c  <=  ~I71b8492d70b423e95938995c07395def + 1;
                end else begin
                    If8a527cc7f06a9963a80a880d225d34c  <= I71b8492d70b423e95938995c07395def ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ibdf2178bd18783c4797c21e642388d16 != I980165c1147ac5ff86619c841c6031dc[1] ) begin
                    Ic3a431f39c678b7175ed30fde1fa6424  <=  ~Iae469bcbba9598bb46aa7ccf9fa06a37 + 1;
                end else begin
                    Ic3a431f39c678b7175ed30fde1fa6424  <= Iae469bcbba9598bb46aa7ccf9fa06a37 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ibdf2178bd18783c4797c21e642388d16 != I0e0b15868b02ca52b260f17f150d237e[0] ) begin
                    I4af080cb4e5cc525db95e5f401019e8c  <=  ~Ie2e854376f4b6509ec41507401173269 + 1;
                end else begin
                    I4af080cb4e5cc525db95e5f401019e8c  <= Ie2e854376f4b6509ec41507401173269 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ibdf2178bd18783c4797c21e642388d16 != I6ebab438dc55ccf6c1600313891d9c38[0] ) begin
                    Ic6386d7d8813731d612e24b715740275  <=  ~I7b1401c3c2c389d9bf05658c88ff6b40 + 1;
                end else begin
                    Ic6386d7d8813731d612e24b715740275  <= I7b1401c3c2c389d9bf05658c88ff6b40 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ibdf2178bd18783c4797c21e642388d16 != I07930a807994815de45864af579902c4[1] ) begin
                    Ic512effb493a06ece58a2af155135004  <=  ~I88ee95aeb6c744eca0e127e8497b5dc9 + 1;
                end else begin
                    Ic512effb493a06ece58a2af155135004  <= I88ee95aeb6c744eca0e127e8497b5dc9 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ibdf2178bd18783c4797c21e642388d16 != I6f5c991e5fdcf56d582c6f80eb6731df[1] ) begin
                    I9b6a674dbcbfcf65f1ae0deb8fc3566d  <=  ~I5573e18ade3430ef3eff5e6d960e44eb + 1;
                end else begin
                    I9b6a674dbcbfcf65f1ae0deb8fc3566d  <= I5573e18ade3430ef3eff5e6d960e44eb ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ibdf2178bd18783c4797c21e642388d16 != Ieb244944e7ee8236a207924f56fbc689[0] ) begin
                    Ib4bdc9069d0c08655f5e87f705943eda  <=  ~Id6260fa8a9be077673e82344c736b1c4 + 1;
                end else begin
                    Ib4bdc9069d0c08655f5e87f705943eda  <= Id6260fa8a9be077673e82344c736b1c4 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I2c690809d9b9e3482fe5a133b5c00afa != Ib58043c04b5c4c86c1c67e57cc66dcf7[1] ) begin
                    If92db65b39a83e1c699e4cc6d7f9e57b  <=  ~Ic052eadb342350c52d89e73d5fea80bb + 1;
                end else begin
                    If92db65b39a83e1c699e4cc6d7f9e57b  <= Ic052eadb342350c52d89e73d5fea80bb ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I2c690809d9b9e3482fe5a133b5c00afa != I9c0b88a0be66d62f8ab061aeaee7e60f[1] ) begin
                    I0262b30a4efa9f1cfb11d1c3940de9e7  <=  ~I98b8d024432fc54ebf2f15d99968f2e0 + 1;
                end else begin
                    I0262b30a4efa9f1cfb11d1c3940de9e7  <= I98b8d024432fc54ebf2f15d99968f2e0 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I2c690809d9b9e3482fe5a133b5c00afa != I8e29ebe9ee25ea8ef3e52ff56fc29157[0] ) begin
                    Ie8df350430970b5f1229cda772440f85  <=  ~I98f54ab8454940141a484332f2a05369 + 1;
                end else begin
                    Ie8df350430970b5f1229cda772440f85  <= I98f54ab8454940141a484332f2a05369 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I2c690809d9b9e3482fe5a133b5c00afa != I50976b0051e84b6a42fc1dbabd7d20ae[0] ) begin
                    I8070a3b7d8b1a7ae90c1a2d27aed09aa  <=  ~I9d94ad2da06ac1fef4da7dcc56abffca + 1;
                end else begin
                    I8070a3b7d8b1a7ae90c1a2d27aed09aa  <= I9d94ad2da06ac1fef4da7dcc56abffca ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I2c690809d9b9e3482fe5a133b5c00afa != I19df055705f322292a3601fa63f0e5f9[1] ) begin
                    I39bbec42c442d1e8c818f46ad9c096a8  <=  ~I51262e3abe460148e3c2d2b74989c2b8 + 1;
                end else begin
                    I39bbec42c442d1e8c818f46ad9c096a8  <= I51262e3abe460148e3c2d2b74989c2b8 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I2c690809d9b9e3482fe5a133b5c00afa != I3c0b6f53f0a5cda5b6758b2ee2c83b92[0] ) begin
                    I9bb81dda8102b829441be46460eb8900  <=  ~I560583680bb2f5a0b5ede42ceaafcf8b + 1;
                end else begin
                    I9bb81dda8102b829441be46460eb8900  <= I560583680bb2f5a0b5ede42ceaafcf8b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I2c690809d9b9e3482fe5a133b5c00afa != I2fbf89398a148c47810456812dbee5a6[0] ) begin
                    Ib23edc35fa5bbfe0415fcf0861a22d9b  <=  ~I389f83346ffaffe8186fb0074d71f43c + 1;
                end else begin
                    Ib23edc35fa5bbfe0415fcf0861a22d9b  <= I389f83346ffaffe8186fb0074d71f43c ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I2c690809d9b9e3482fe5a133b5c00afa != I72a2f42b727a0503d43332c0f22d5ae3[1] ) begin
                    I9cc16a00912e7dfc05fb505a9db23cd8  <=  ~Ie89c2a1b3943d12197bb972bd12595b0 + 1;
                end else begin
                    I9cc16a00912e7dfc05fb505a9db23cd8  <= Ie89c2a1b3943d12197bb972bd12595b0 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I2c690809d9b9e3482fe5a133b5c00afa != Ia5cc3055ba3365e64cf59c4d4fd3f093[1] ) begin
                    Iccefa45795486757515d95e5908b306a  <=  ~Ic7be56919976a2d1088114c21c3c1ffb + 1;
                end else begin
                    Iccefa45795486757515d95e5908b306a  <= Ic7be56919976a2d1088114c21c3c1ffb ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I2c690809d9b9e3482fe5a133b5c00afa != Ie9b2be4c32334220e134e041ca8dfc06[0] ) begin
                    Ic3a608b850709286ea0ad2f67425d9ac  <=  ~Icb5dab0df062ab46bd3d1a73e85ef4c2 + 1;
                end else begin
                    Ic3a608b850709286ea0ad2f67425d9ac  <= Icb5dab0df062ab46bd3d1a73e85ef4c2 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I369ffa98995ba0834f8029ecce705c56 != Ibc0871b3c992fd278815fdbefcd2bac0[1] ) begin
                    I2213c1a2b831f421707a261f5a58b1b1  <=  ~I27a568cfc2df13cf689d366a25e5d05f + 1;
                end else begin
                    I2213c1a2b831f421707a261f5a58b1b1  <= I27a568cfc2df13cf689d366a25e5d05f ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I369ffa98995ba0834f8029ecce705c56 != Id88b9265ff08e0730e6a41abe1f80a32[1] ) begin
                    I4636821315d702a677dc93113872e647  <=  ~Ia6688964078f1ea87b742352877aac45 + 1;
                end else begin
                    I4636821315d702a677dc93113872e647  <= Ia6688964078f1ea87b742352877aac45 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I369ffa98995ba0834f8029ecce705c56 != Ic3742290179b27b9865f9d1f88d66266[0] ) begin
                    Iaf8a19fde3de660c3fa925593bebbe0c  <=  ~I180deab4fe0d03104cf2ee035f6a9b8c + 1;
                end else begin
                    Iaf8a19fde3de660c3fa925593bebbe0c  <= I180deab4fe0d03104cf2ee035f6a9b8c ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I369ffa98995ba0834f8029ecce705c56 != I82e0e091fba6f79cef97eacac4b43ecb[0] ) begin
                    I0052d562fb3182890c8828e52d437b11  <=  ~Iff6cd034bb64d13c21910c11bd92266e + 1;
                end else begin
                    I0052d562fb3182890c8828e52d437b11  <= Iff6cd034bb64d13c21910c11bd92266e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I369ffa98995ba0834f8029ecce705c56 != I3d50cfeaa4b69c09bb648b8873a6bc24[1] ) begin
                    I21668ff77cf75570cae97f575cbcf644  <=  ~I7c34057a77f2bdda93c422506959818d + 1;
                end else begin
                    I21668ff77cf75570cae97f575cbcf644  <= I7c34057a77f2bdda93c422506959818d ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I369ffa98995ba0834f8029ecce705c56 != I8e591d83170c8ba46d31c61935311b22[0] ) begin
                    Ic279867ebf3055980f3d813d5dc8dec6  <=  ~I7ff7d3fd63fa67cd72d1591c1a373180 + 1;
                end else begin
                    Ic279867ebf3055980f3d813d5dc8dec6  <= I7ff7d3fd63fa67cd72d1591c1a373180 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I369ffa98995ba0834f8029ecce705c56 != Icac5a9001ee113e612e3457b4b49ee68[0] ) begin
                    Ifc8c6df8904b97674f2970ebc95b523c  <=  ~If910e75bf10cf02a5b414cbb4fad1304 + 1;
                end else begin
                    Ifc8c6df8904b97674f2970ebc95b523c  <= If910e75bf10cf02a5b414cbb4fad1304 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I369ffa98995ba0834f8029ecce705c56 != I8b8b9c4777e6df3eb2b9313e69ef2c8c[1] ) begin
                    Id88480a0a350bb5fcf01ed5fff0bbd4c  <=  ~I266697a6eca2b73a76fd375a0ad72a05 + 1;
                end else begin
                    Id88480a0a350bb5fcf01ed5fff0bbd4c  <= I266697a6eca2b73a76fd375a0ad72a05 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I369ffa98995ba0834f8029ecce705c56 != Iea7da1f43ba202d753b0edb0be8b3fcf[1] ) begin
                    If38feb4f76f761dce6145731ad235d7f  <=  ~Iba188abd7715fcbdad3b1f3d985c6fc3 + 1;
                end else begin
                    If38feb4f76f761dce6145731ad235d7f  <= Iba188abd7715fcbdad3b1f3d985c6fc3 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I369ffa98995ba0834f8029ecce705c56 != Id6f07dee3e47f39e3b43329c26f690f7[0] ) begin
                    Ieb528d666fdb708279184bb59eac25d9  <=  ~Ic60c640562e3e45c89a1de78af509b6a + 1;
                end else begin
                    Ieb528d666fdb708279184bb59eac25d9  <= Ic60c640562e3e45c89a1de78af509b6a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9ccef4c47ae7cfab43584de0f2e193d3 != I8695e1e94cbfcbe4b9eae315b042529e[1] ) begin
                    I631a3300cb6685f47da7781940ec5d27  <=  ~I0456494b33e4ec852c123cb3003b9886 + 1;
                end else begin
                    I631a3300cb6685f47da7781940ec5d27  <= I0456494b33e4ec852c123cb3003b9886 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9ccef4c47ae7cfab43584de0f2e193d3 != I6330943c9295298c53e889d47c7904d9[1] ) begin
                    Ib54d55a70605119e37e9898b940ff636  <=  ~I2ed7c217fe3e21fcb27e04f68b95dd6b + 1;
                end else begin
                    Ib54d55a70605119e37e9898b940ff636  <= I2ed7c217fe3e21fcb27e04f68b95dd6b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9ccef4c47ae7cfab43584de0f2e193d3 != I9ef21ef20099af28d9a8c794f70d45a5[0] ) begin
                    I49fb0909ddf66fc0073e6400f1a07844  <=  ~Ifda5780b42bf451a7ce834f17b3fdd20 + 1;
                end else begin
                    I49fb0909ddf66fc0073e6400f1a07844  <= Ifda5780b42bf451a7ce834f17b3fdd20 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9ccef4c47ae7cfab43584de0f2e193d3 != I04302edb2671c5bc0ca2673cd53935e1[0] ) begin
                    Id0eef1adba01447c14a6f005782dd9a2  <=  ~Iadca92fd39d1fd6032feb8415ca5246f + 1;
                end else begin
                    Id0eef1adba01447c14a6f005782dd9a2  <= Iadca92fd39d1fd6032feb8415ca5246f ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9ccef4c47ae7cfab43584de0f2e193d3 != I33a6ffad80ddf99a4d316a049078244d[1] ) begin
                    I5a9fdec7d7ff99fe33ad6cd8afd9e059  <=  ~I613453382f19dd7eb9bdf51e945a33b0 + 1;
                end else begin
                    I5a9fdec7d7ff99fe33ad6cd8afd9e059  <= I613453382f19dd7eb9bdf51e945a33b0 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9ccef4c47ae7cfab43584de0f2e193d3 != I02b62fafd371de339f299f8aefec6c43[0] ) begin
                    I68528be9951f5b8805411711cd11ea59  <=  ~Ideafa683e6a3a38848fb8bee22eba11b + 1;
                end else begin
                    I68528be9951f5b8805411711cd11ea59  <= Ideafa683e6a3a38848fb8bee22eba11b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9ccef4c47ae7cfab43584de0f2e193d3 != I9461e92a5880cb9e04fcece2ef4674f0[0] ) begin
                    Ia3450e134e4086c35acbdee1e6042396  <=  ~Ie4226e7e17c7971f07aaf0cfaeae495a + 1;
                end else begin
                    Ia3450e134e4086c35acbdee1e6042396  <= Ie4226e7e17c7971f07aaf0cfaeae495a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9ccef4c47ae7cfab43584de0f2e193d3 != I4a16e8e7946d9a8220304fc1be3fb362[1] ) begin
                    Ifec374bce7f5507438f550df22d61a01  <=  ~Ifbbfa268bd4c31c7eed45cd43fe6a405 + 1;
                end else begin
                    Ifec374bce7f5507438f550df22d61a01  <= Ifbbfa268bd4c31c7eed45cd43fe6a405 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9ccef4c47ae7cfab43584de0f2e193d3 != I872f61d20baf011e867b44dc5539fc37[1] ) begin
                    Ie87075ac979410cc11099a356966b8a2  <=  ~Ib2d99d95f7a31e4745211c5ff96f851c + 1;
                end else begin
                    Ie87075ac979410cc11099a356966b8a2  <= Ib2d99d95f7a31e4745211c5ff96f851c ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9ccef4c47ae7cfab43584de0f2e193d3 != Ic7f04c065f8ff82c2288f1de77d37189[0] ) begin
                    If4d3b31b87c0f723241d35ce7e854eba  <=  ~I692c0a91b415b400a3640e2d9a40edad + 1;
                end else begin
                    If4d3b31b87c0f723241d35ce7e854eba  <= I692c0a91b415b400a3640e2d9a40edad ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ief31fe169c1b360d5933558208dbb602 != Ibc0871b3c992fd278815fdbefcd2bac0[2] ) begin
                    Ic53b875b2ddcba11406eb2ca39354757  <=  ~If8c4dc70212e8873167e1cad8e8e5692 + 1;
                end else begin
                    Ic53b875b2ddcba11406eb2ca39354757  <= If8c4dc70212e8873167e1cad8e8e5692 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ief31fe169c1b360d5933558208dbb602 != Iceb64ab2ff8a2e0dfdb74803811d4cfe[1] ) begin
                    Ie19b39200436b0bfca13502ad36c21b9  <=  ~Ib2f75e91bf9e1d32a3f170fc85244139 + 1;
                end else begin
                    Ie19b39200436b0bfca13502ad36c21b9  <= Ib2f75e91bf9e1d32a3f170fc85244139 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ief31fe169c1b360d5933558208dbb602 != Id88b9265ff08e0730e6a41abe1f80a32[2] ) begin
                    I9c981b0614a29386ca5e8ebc06a17f15  <=  ~I3606dc61f24567cb1ace443cea62a43b + 1;
                end else begin
                    I9c981b0614a29386ca5e8ebc06a17f15  <= I3606dc61f24567cb1ace443cea62a43b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ief31fe169c1b360d5933558208dbb602 != I9ef21ef20099af28d9a8c794f70d45a5[1] ) begin
                    I9938397dc94002481984f5b560fadc58  <=  ~Ie402c9f793b7306323efb8fe23533250 + 1;
                end else begin
                    I9938397dc94002481984f5b560fadc58  <= Ie402c9f793b7306323efb8fe23533250 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ief31fe169c1b360d5933558208dbb602 != I6ebab438dc55ccf6c1600313891d9c38[1] ) begin
                    I4c366a57920ff090a98a2cb8b9caa00b  <=  ~I54652565023310e2eccfc4cb87c56b43 + 1;
                end else begin
                    I4c366a57920ff090a98a2cb8b9caa00b  <= I54652565023310e2eccfc4cb87c56b43 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ief31fe169c1b360d5933558208dbb602 != Ic2580cbeec8c11a19bd1e2ebc29d255e[1] ) begin
                    Ieafa9d74d4a61d28ac4a913db460bf33  <=  ~I616b7a5987edbc001e0ae1b638f25a39 + 1;
                end else begin
                    Ieafa9d74d4a61d28ac4a913db460bf33  <= I616b7a5987edbc001e0ae1b638f25a39 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ief31fe169c1b360d5933558208dbb602 != Ieb244944e7ee8236a207924f56fbc689[1] ) begin
                    Idbf9094c94c931f16fba468b9dd59a25  <=  ~I06604bac478ee906b3fe8ff307cdf046 + 1;
                end else begin
                    Idbf9094c94c931f16fba468b9dd59a25  <= I06604bac478ee906b3fe8ff307cdf046 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ief31fe169c1b360d5933558208dbb602 != I4267622319ca65909a3b40484dc74d3a[0] ) begin
                    I8d8d95ff26f33f69a182b32ccde23905  <=  ~I135dd8a85aca863db660f2ad4f80ca2e + 1;
                end else begin
                    I8d8d95ff26f33f69a182b32ccde23905  <= I135dd8a85aca863db660f2ad4f80ca2e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib8c0317dafcfb91b3da5eb5afae1f2e2 != I8695e1e94cbfcbe4b9eae315b042529e[2] ) begin
                    I8bbe1a2ace8f51aa22cca5d9fc66f136  <=  ~I8715d73b58270dfa33b903e9cfb50be8 + 1;
                end else begin
                    I8bbe1a2ace8f51aa22cca5d9fc66f136  <= I8715d73b58270dfa33b903e9cfb50be8 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib8c0317dafcfb91b3da5eb5afae1f2e2 != I5b7caaeb34c43e66e8d095a859e708fe[1] ) begin
                    If0a3b88a66a816b25f17ced5d0e8f775  <=  ~I7f60cb59895af6d314f5d0f401c80350 + 1;
                end else begin
                    If0a3b88a66a816b25f17ced5d0e8f775  <= I7f60cb59895af6d314f5d0f401c80350 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib8c0317dafcfb91b3da5eb5afae1f2e2 != I6330943c9295298c53e889d47c7904d9[2] ) begin
                    If7e146da4f3bd255b8457fd6902005f6  <=  ~I3e25e6e9de5ee9242a472ce957056762 + 1;
                end else begin
                    If7e146da4f3bd255b8457fd6902005f6  <= I3e25e6e9de5ee9242a472ce957056762 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib8c0317dafcfb91b3da5eb5afae1f2e2 != Ic2941d16ae6a5cbce70e8546a18ca4ff[1] ) begin
                    I89a3f8d5f760d1a650f85814cbfdc017  <=  ~I4c5f36517aaf872e7f05de2f7f76a6ce + 1;
                end else begin
                    I89a3f8d5f760d1a650f85814cbfdc017  <= I4c5f36517aaf872e7f05de2f7f76a6ce ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib8c0317dafcfb91b3da5eb5afae1f2e2 != I2fbf89398a148c47810456812dbee5a6[1] ) begin
                    I3e0e682047f7cc36142e668828cbff1e  <=  ~I0e993e6f98616632f17835a2994f45e3 + 1;
                end else begin
                    I3e0e682047f7cc36142e668828cbff1e  <= I0e993e6f98616632f17835a2994f45e3 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib8c0317dafcfb91b3da5eb5afae1f2e2 != If79ed5ee2b8710da0608c1e245d07d55[1] ) begin
                    I596ad7e132f272cb196b74faa8c75aa4  <=  ~I281f996740b16568b9d29ca41a3fa50d + 1;
                end else begin
                    I596ad7e132f272cb196b74faa8c75aa4  <= I281f996740b16568b9d29ca41a3fa50d ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib8c0317dafcfb91b3da5eb5afae1f2e2 != Ie9b2be4c32334220e134e041ca8dfc06[1] ) begin
                    I5267fa34449e6eebe891017fc32d0749  <=  ~I55bbb73d68871d9dbce4d590c029aeab + 1;
                end else begin
                    I5267fa34449e6eebe891017fc32d0749  <= I55bbb73d68871d9dbce4d590c029aeab ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib8c0317dafcfb91b3da5eb5afae1f2e2 != Iedd7d4ea8d082b40244c04946dfb14a0[0] ) begin
                    I2dc64c3b06588542b027f997437bee63  <=  ~Ida491561008f4984480d1b0f09d2fa77 + 1;
                end else begin
                    I2dc64c3b06588542b027f997437bee63  <= Ida491561008f4984480d1b0f09d2fa77 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I54e3f08f6f4cf784da57ac39f246b8fd != Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[2] ) begin
                    I753f92da60980736440aba814a156f1e  <=  ~I624e237f248d292c0417ff85056857b0 + 1;
                end else begin
                    I753f92da60980736440aba814a156f1e  <= I624e237f248d292c0417ff85056857b0 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I54e3f08f6f4cf784da57ac39f246b8fd != I61f0c04673dfb262ef6912eb2df39120[1] ) begin
                    I733605337bf6972630c089d32fd7f98f  <=  ~Ic7c1fd79ba76dbb254c6183017f40b3e + 1;
                end else begin
                    I733605337bf6972630c089d32fd7f98f  <= Ic7c1fd79ba76dbb254c6183017f40b3e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I54e3f08f6f4cf784da57ac39f246b8fd != I5686b595177e07dd5bf231a35ee41659[2] ) begin
                    Iba70e737d52e6812a67c159520e5192f  <=  ~I546d683af76dc209a5205c6274abe908 + 1;
                end else begin
                    Iba70e737d52e6812a67c159520e5192f  <= I546d683af76dc209a5205c6274abe908 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I54e3f08f6f4cf784da57ac39f246b8fd != I8e29ebe9ee25ea8ef3e52ff56fc29157[1] ) begin
                    I7d77ac9b64b2e8cae21c6e36947e3ca2  <=  ~I7b4bb785489c5bb22c84d9778192fe44 + 1;
                end else begin
                    I7d77ac9b64b2e8cae21c6e36947e3ca2  <= I7b4bb785489c5bb22c84d9778192fe44 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I54e3f08f6f4cf784da57ac39f246b8fd != Icac5a9001ee113e612e3457b4b49ee68[1] ) begin
                    Icd0622a90782b9c451950e7ab0399567  <=  ~Ifc6af7d7aeb7162d554b8604a44f3361 + 1;
                end else begin
                    Icd0622a90782b9c451950e7ab0399567  <= Ifc6af7d7aeb7162d554b8604a44f3361 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I54e3f08f6f4cf784da57ac39f246b8fd != I9497bbb4f746969a95cff948a3ee9ade[1] ) begin
                    I1487170cb1f3370ad45efc801cefc8ab  <=  ~I5b650c4c3291670b480a7f1095093dfb + 1;
                end else begin
                    I1487170cb1f3370ad45efc801cefc8ab  <= I5b650c4c3291670b480a7f1095093dfb ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I54e3f08f6f4cf784da57ac39f246b8fd != Id6f07dee3e47f39e3b43329c26f690f7[1] ) begin
                    Ic3ff7ce12c836bf0693252b9a7a7cfe8  <=  ~I2f5f88cb5e5e4723bd8a83c5fa80cc4c + 1;
                end else begin
                    Ic3ff7ce12c836bf0693252b9a7a7cfe8  <= I2f5f88cb5e5e4723bd8a83c5fa80cc4c ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I54e3f08f6f4cf784da57ac39f246b8fd != I56e1fe0c7a62589c123876f2b4e57a26[0] ) begin
                    Ib23d889edb5a6d9f27de977d3b1a2616  <=  ~Ic174b361182c98486e65b7f87b073274 + 1;
                end else begin
                    Ib23d889edb5a6d9f27de977d3b1a2616  <= Ic174b361182c98486e65b7f87b073274 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I16c7f1b874b0d05c6d120bbede254416 != Ib58043c04b5c4c86c1c67e57cc66dcf7[2] ) begin
                    I8f2986bc015fcc64ac5e5395ac6dd851  <=  ~I7ba2f7201745258dbf224de087a25233 + 1;
                end else begin
                    I8f2986bc015fcc64ac5e5395ac6dd851  <= I7ba2f7201745258dbf224de087a25233 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I16c7f1b874b0d05c6d120bbede254416 != Ibeb5edab51cd6aedad9c2ecedaded6f5[1] ) begin
                    I7d5041a6796c00188f74936d283defe6  <=  ~I131a4bd335fc23ee10f7ccb1881ab9cd + 1;
                end else begin
                    I7d5041a6796c00188f74936d283defe6  <= I131a4bd335fc23ee10f7ccb1881ab9cd ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I16c7f1b874b0d05c6d120bbede254416 != I9c0b88a0be66d62f8ab061aeaee7e60f[2] ) begin
                    I7a2e79d42779ad235bca6ce3757cf588  <=  ~I90cb3e06b42f25956b788a792eef371f + 1;
                end else begin
                    I7a2e79d42779ad235bca6ce3757cf588  <= I90cb3e06b42f25956b788a792eef371f ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I16c7f1b874b0d05c6d120bbede254416 != Ic3742290179b27b9865f9d1f88d66266[1] ) begin
                    Icd1da43a4d95230e79dbd35a7ae41066  <=  ~I56302770a8d56932e7bb5dcff56c71e2 + 1;
                end else begin
                    Icd1da43a4d95230e79dbd35a7ae41066  <= I56302770a8d56932e7bb5dcff56c71e2 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I16c7f1b874b0d05c6d120bbede254416 != I9461e92a5880cb9e04fcece2ef4674f0[1] ) begin
                    I5a0f27df5158309f32f0df31e8ae3ae3  <=  ~Id3b8c058b3838c388eb5ddcb31dfc799 + 1;
                end else begin
                    I5a0f27df5158309f32f0df31e8ae3ae3  <= Id3b8c058b3838c388eb5ddcb31dfc799 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I16c7f1b874b0d05c6d120bbede254416 != I651d700a00d7004d8728bc7356f30926[1] ) begin
                    I4255ac1af4367c321567c4e46b06ab25  <=  ~I7ca8ce63dfb821d10304958bada71737 + 1;
                end else begin
                    I4255ac1af4367c321567c4e46b06ab25  <= I7ca8ce63dfb821d10304958bada71737 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I16c7f1b874b0d05c6d120bbede254416 != Ic7f04c065f8ff82c2288f1de77d37189[1] ) begin
                    I72369dedfe36cb22269033cc305b730c  <=  ~I06ad44414b45d262f9542015d2dead8d + 1;
                end else begin
                    I72369dedfe36cb22269033cc305b730c  <= I06ad44414b45d262f9542015d2dead8d ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I16c7f1b874b0d05c6d120bbede254416 != Ia8a468877c9f96713c8141df9205f92a[0] ) begin
                    Ie65a0634454381e24bb3223a333e3ad0  <=  ~I833ef4acfed17e4699d65cbaa3e7dbd5 + 1;
                end else begin
                    Ie65a0634454381e24bb3223a333e3ad0  <= I833ef4acfed17e4699d65cbaa3e7dbd5 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I0c3cb2de514ecab0dd311e86a4dc3cdb != I61f0c04673dfb262ef6912eb2df39120[2] ) begin
                    Idcb1d8bbdeaed6768c2a418c3048e6ee  <=  ~Ia77e3db939408af719e0a8555dcb68ed + 1;
                end else begin
                    Idcb1d8bbdeaed6768c2a418c3048e6ee  <= Ia77e3db939408af719e0a8555dcb68ed ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I0c3cb2de514ecab0dd311e86a4dc3cdb != Ie1cd04c7668d3f450c387a6c1ad778c7[1] ) begin
                    If3e5161254eb9056914c46263b865c10  <=  ~I57ab4999187992eda55a82bf0f09b31f + 1;
                end else begin
                    If3e5161254eb9056914c46263b865c10  <= I57ab4999187992eda55a82bf0f09b31f ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I0c3cb2de514ecab0dd311e86a4dc3cdb != I8e29ebe9ee25ea8ef3e52ff56fc29157[2] ) begin
                    Ic1faed76fca5a9ceb7db26c2f43623d9  <=  ~I21f7b5402ae8e8954d99931bd5108250 + 1;
                end else begin
                    Ic1faed76fca5a9ceb7db26c2f43623d9  <= I21f7b5402ae8e8954d99931bd5108250 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I0c3cb2de514ecab0dd311e86a4dc3cdb != I04302edb2671c5bc0ca2673cd53935e1[1] ) begin
                    I1d1a7c5928982c278d068ebd262254da  <=  ~I3627708869b47d460182bc5040092f9a + 1;
                end else begin
                    I1d1a7c5928982c278d068ebd262254da  <= I3627708869b47d460182bc5040092f9a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I0c3cb2de514ecab0dd311e86a4dc3cdb != I33a6ffad80ddf99a4d316a049078244d[2] ) begin
                    I47b1695a74e4d27389b97543415dcc67  <=  ~Ifd88f0f0abd1c037434dc16e34550d2a + 1;
                end else begin
                    I47b1695a74e4d27389b97543415dcc67  <= Ifd88f0f0abd1c037434dc16e34550d2a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I0c3cb2de514ecab0dd311e86a4dc3cdb != I8e591d83170c8ba46d31c61935311b22[1] ) begin
                    I5c05da8a222ad5effb9815cbf3ec25f3  <=  ~I27eec53da48406e7e1202345a0810e08 + 1;
                end else begin
                    I5c05da8a222ad5effb9815cbf3ec25f3  <= I27eec53da48406e7e1202345a0810e08 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I0c3cb2de514ecab0dd311e86a4dc3cdb != Icac5a9001ee113e612e3457b4b49ee68[2] ) begin
                    I6493b3c087d4685a6b3f98c73dc2ff49  <=  ~I682d42afaaf103550ce4fbdba6192c88 + 1;
                end else begin
                    I6493b3c087d4685a6b3f98c73dc2ff49  <= I682d42afaaf103550ce4fbdba6192c88 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I0c3cb2de514ecab0dd311e86a4dc3cdb != I07930a807994815de45864af579902c4[2] ) begin
                    I2c72248cbe49ec0a0febac2437b8a6dc  <=  ~If225534847db8723768941c3819ed7c0 + 1;
                end else begin
                    I2c72248cbe49ec0a0febac2437b8a6dc  <= If225534847db8723768941c3819ed7c0 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I0c3cb2de514ecab0dd311e86a4dc3cdb != Ic2580cbeec8c11a19bd1e2ebc29d255e[2] ) begin
                    I6fd1b4395af175eff85b3bfeef4c329b  <=  ~I43a91b2232a47d1f6731bafc15ced5db + 1;
                end else begin
                    I6fd1b4395af175eff85b3bfeef4c329b  <= I43a91b2232a47d1f6731bafc15ced5db ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I0c3cb2de514ecab0dd311e86a4dc3cdb != I4267622319ca65909a3b40484dc74d3a[1] ) begin
                    I2508854bcbab37bd09c9465c377c06aa  <=  ~Ic54026604afd19b0c7c71ea1ac0f1c4e + 1;
                end else begin
                    I2508854bcbab37bd09c9465c377c06aa  <= Ic54026604afd19b0c7c71ea1ac0f1c4e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Icc5ba4554d7a44bc3b43377efbe3b5f8 != Ibeb5edab51cd6aedad9c2ecedaded6f5[2] ) begin
                    Iba7608ee0a01af103e022bcaf564bf6b  <=  ~I218bd69f079aa21f0dda241ae6e387ad + 1;
                end else begin
                    Iba7608ee0a01af103e022bcaf564bf6b  <= I218bd69f079aa21f0dda241ae6e387ad ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Icc5ba4554d7a44bc3b43377efbe3b5f8 != If511a6ea6aa5cda5353658d8e192791f[1] ) begin
                    Ia9642d79bb50567348083b4435c7d66d  <=  ~Iaaacca4d06ad0f202d839fd7674f1829 + 1;
                end else begin
                    Ia9642d79bb50567348083b4435c7d66d  <= Iaaacca4d06ad0f202d839fd7674f1829 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Icc5ba4554d7a44bc3b43377efbe3b5f8 != Ic3742290179b27b9865f9d1f88d66266[2] ) begin
                    Ice9079fb6e08d629f8c0c9ce332c8f11  <=  ~Iecddac410bb2121da0df2d73c2d23cb8 + 1;
                end else begin
                    Ice9079fb6e08d629f8c0c9ce332c8f11  <= Iecddac410bb2121da0df2d73c2d23cb8 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Icc5ba4554d7a44bc3b43377efbe3b5f8 != I480a0f6d6c3eb936de10a72749f6cd3f[1] ) begin
                    I39ff4663007dbc89b403f3b08a69bb6c  <=  ~I1aabc0c0b7b602297ad592ae48b23452 + 1;
                end else begin
                    I39ff4663007dbc89b403f3b08a69bb6c  <= I1aabc0c0b7b602297ad592ae48b23452 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Icc5ba4554d7a44bc3b43377efbe3b5f8 != I980165c1147ac5ff86619c841c6031dc[2] ) begin
                    Ib01cfd833a63500e03333f263805db3d  <=  ~Ida3aaf7237b1383cfe95eeccf3971a8e + 1;
                end else begin
                    Ib01cfd833a63500e03333f263805db3d  <= Ida3aaf7237b1383cfe95eeccf3971a8e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Icc5ba4554d7a44bc3b43377efbe3b5f8 != I02b62fafd371de339f299f8aefec6c43[1] ) begin
                    I0f034a8f077b0ab231727b6298e366d8  <=  ~Idd2a8ed39edf6697b0988ee4eb4f2d95 + 1;
                end else begin
                    I0f034a8f077b0ab231727b6298e366d8  <= Idd2a8ed39edf6697b0988ee4eb4f2d95 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Icc5ba4554d7a44bc3b43377efbe3b5f8 != I9461e92a5880cb9e04fcece2ef4674f0[2] ) begin
                    I17d9e19854cef197fd3267618617efc3  <=  ~I735c660d5232e03dd8fb129e2ca4b445 + 1;
                end else begin
                    I17d9e19854cef197fd3267618617efc3  <= I735c660d5232e03dd8fb129e2ca4b445 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Icc5ba4554d7a44bc3b43377efbe3b5f8 != I72a2f42b727a0503d43332c0f22d5ae3[2] ) begin
                    Iacf9640cbf486411d6ceb8fe1a2fd5c9  <=  ~Ia04d6065987df3f007658614406cbc28 + 1;
                end else begin
                    Iacf9640cbf486411d6ceb8fe1a2fd5c9  <= Ia04d6065987df3f007658614406cbc28 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Icc5ba4554d7a44bc3b43377efbe3b5f8 != If79ed5ee2b8710da0608c1e245d07d55[2] ) begin
                    Idc629414f6d0236ce0714cfaae23f065  <=  ~I7aeddde5b60828ac7f8b6c2addaf220b + 1;
                end else begin
                    Idc629414f6d0236ce0714cfaae23f065  <= I7aeddde5b60828ac7f8b6c2addaf220b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Icc5ba4554d7a44bc3b43377efbe3b5f8 != Iedd7d4ea8d082b40244c04946dfb14a0[1] ) begin
                    Id92a37c091100e9df08e24498ecb4022  <=  ~I150c28296847348d69cce123f20656c3 + 1;
                end else begin
                    Id92a37c091100e9df08e24498ecb4022  <= I150c28296847348d69cce123f20656c3 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I5e51f49adb6dce65a9f19ff736526c4b != Iceb64ab2ff8a2e0dfdb74803811d4cfe[2] ) begin
                    If6657f90c84ca5e2ba08ec705f34be03  <=  ~Ib94d38d19b3791fa2d1b42fdfde8435e + 1;
                end else begin
                    If6657f90c84ca5e2ba08ec705f34be03  <= Ib94d38d19b3791fa2d1b42fdfde8435e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I5e51f49adb6dce65a9f19ff736526c4b != Ib0bf69cc797f330fb2546eb46d2d6f76[1] ) begin
                    Ic51bb9184dfd103703cd0c6ad6edff4b  <=  ~I94865622898b2e481e86a244f7aa2759 + 1;
                end else begin
                    Ic51bb9184dfd103703cd0c6ad6edff4b  <= I94865622898b2e481e86a244f7aa2759 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I5e51f49adb6dce65a9f19ff736526c4b != I9ef21ef20099af28d9a8c794f70d45a5[2] ) begin
                    I4378d139db4b710e3587aa72df22b70d  <=  ~I1a4a432e735367f515ca747cef7d7d04 + 1;
                end else begin
                    I4378d139db4b710e3587aa72df22b70d  <= I1a4a432e735367f515ca747cef7d7d04 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I5e51f49adb6dce65a9f19ff736526c4b != I50976b0051e84b6a42fc1dbabd7d20ae[1] ) begin
                    Ie88285ce2b9c71de02ebd62e8f44ca72  <=  ~Ib3a2b744d8f38671a63da6f8f8f1a6a1 + 1;
                end else begin
                    Ie88285ce2b9c71de02ebd62e8f44ca72  <= Ib3a2b744d8f38671a63da6f8f8f1a6a1 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I5e51f49adb6dce65a9f19ff736526c4b != I19df055705f322292a3601fa63f0e5f9[2] ) begin
                    I88f1b5c12759a5efb2d2ded8483c9ed2  <=  ~I87716ad5a64592abb812ffe041ccc163 + 1;
                end else begin
                    I88f1b5c12759a5efb2d2ded8483c9ed2  <= I87716ad5a64592abb812ffe041ccc163 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I5e51f49adb6dce65a9f19ff736526c4b != I0e0b15868b02ca52b260f17f150d237e[1] ) begin
                    I6fc8044eb226a14ff1a786ddc96d2414  <=  ~I71b259faefbea7ce8f47e0ffb556a0be + 1;
                end else begin
                    I6fc8044eb226a14ff1a786ddc96d2414  <= I71b259faefbea7ce8f47e0ffb556a0be ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I5e51f49adb6dce65a9f19ff736526c4b != I6ebab438dc55ccf6c1600313891d9c38[2] ) begin
                    I14cf5d43fc9864820a8a25efcc5c6d86  <=  ~I2161b2ff3514dbdbb79d25da87eeec2b + 1;
                end else begin
                    I14cf5d43fc9864820a8a25efcc5c6d86  <= I2161b2ff3514dbdbb79d25da87eeec2b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I5e51f49adb6dce65a9f19ff736526c4b != I8b8b9c4777e6df3eb2b9313e69ef2c8c[2] ) begin
                    I1d9b9ff357667a362f0442f19986f451  <=  ~I860a3c9fca8d240c68ce3825192353b0 + 1;
                end else begin
                    I1d9b9ff357667a362f0442f19986f451  <= I860a3c9fca8d240c68ce3825192353b0 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I5e51f49adb6dce65a9f19ff736526c4b != I9497bbb4f746969a95cff948a3ee9ade[2] ) begin
                    Id88568dd34fbee42c9cb8cc15ac5c31d  <=  ~Ie4eb18c7e906c9a25c12e9980a9f61cb + 1;
                end else begin
                    Id88568dd34fbee42c9cb8cc15ac5c31d  <= Ie4eb18c7e906c9a25c12e9980a9f61cb ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I5e51f49adb6dce65a9f19ff736526c4b != I56e1fe0c7a62589c123876f2b4e57a26[1] ) begin
                    Ifaff9dd032cf96487be819c59b03000a  <=  ~I20a24846a74af76fa4470d6350546a9a + 1;
                end else begin
                    Ifaff9dd032cf96487be819c59b03000a  <= I20a24846a74af76fa4470d6350546a9a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Id57092394c7cda397f42374df4aa3fec != I5b7caaeb34c43e66e8d095a859e708fe[2] ) begin
                    I0374ada4fe50717f2158468b7ad205d4  <=  ~I90d40f6e9721a7d075512b8b81907453 + 1;
                end else begin
                    I0374ada4fe50717f2158468b7ad205d4  <= I90d40f6e9721a7d075512b8b81907453 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Id57092394c7cda397f42374df4aa3fec != Iec7404bc79c58d4d2538fcdf659e9134[1] ) begin
                    Iee6f2484a381bd42e441ff072ec582e4  <=  ~Ifc4525a25f38affb399004b057d1318c + 1;
                end else begin
                    Iee6f2484a381bd42e441ff072ec582e4  <= Ifc4525a25f38affb399004b057d1318c ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Id57092394c7cda397f42374df4aa3fec != Ic2941d16ae6a5cbce70e8546a18ca4ff[2] ) begin
                    Ifae345c79662c3df3dff0fe68ad68746  <=  ~Icc93649a2050b9ded1e625be936b411f + 1;
                end else begin
                    Ifae345c79662c3df3dff0fe68ad68746  <= Icc93649a2050b9ded1e625be936b411f ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Id57092394c7cda397f42374df4aa3fec != I82e0e091fba6f79cef97eacac4b43ecb[1] ) begin
                    I1eedecb1d8ff505c75be7787199afada  <=  ~Ibcc30c960ae0f29c4efb1266c9e490ac + 1;
                end else begin
                    I1eedecb1d8ff505c75be7787199afada  <= Ibcc30c960ae0f29c4efb1266c9e490ac ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Id57092394c7cda397f42374df4aa3fec != I3d50cfeaa4b69c09bb648b8873a6bc24[2] ) begin
                    Ie48be9e6b6fd63baa104d0a6a4561a1a  <=  ~I3b2ffa79fd2227a24c6468a89f2bd989 + 1;
                end else begin
                    Ie48be9e6b6fd63baa104d0a6a4561a1a  <= I3b2ffa79fd2227a24c6468a89f2bd989 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Id57092394c7cda397f42374df4aa3fec != I3c0b6f53f0a5cda5b6758b2ee2c83b92[1] ) begin
                    I8eef6ca0a61a21882ea28b3d63735228  <=  ~Ib489a11dfdd8a2b3ad561c965b3d7d2a + 1;
                end else begin
                    I8eef6ca0a61a21882ea28b3d63735228  <= Ib489a11dfdd8a2b3ad561c965b3d7d2a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Id57092394c7cda397f42374df4aa3fec != I2fbf89398a148c47810456812dbee5a6[2] ) begin
                    I99fb9030e8361e57818c07511479a9b8  <=  ~Ifa51cf9f9d3d1b91c72387f5daf05c79 + 1;
                end else begin
                    I99fb9030e8361e57818c07511479a9b8  <= Ifa51cf9f9d3d1b91c72387f5daf05c79 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Id57092394c7cda397f42374df4aa3fec != I4a16e8e7946d9a8220304fc1be3fb362[2] ) begin
                    Ief67e897e57b96e2ec200e82bbc7caeb  <=  ~Ifda20d77c574c8f13816620c56fff950 + 1;
                end else begin
                    Ief67e897e57b96e2ec200e82bbc7caeb  <= Ifda20d77c574c8f13816620c56fff950 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Id57092394c7cda397f42374df4aa3fec != I651d700a00d7004d8728bc7356f30926[2] ) begin
                    Ia445bdc7def7d8c1eec31ab892c25c41  <=  ~I03ce0915d3a170429959221b6c8cd16c + 1;
                end else begin
                    Ia445bdc7def7d8c1eec31ab892c25c41  <= I03ce0915d3a170429959221b6c8cd16c ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Id57092394c7cda397f42374df4aa3fec != Ia8a468877c9f96713c8141df9205f92a[1] ) begin
                    Iad166146f7df5e8068fc6efe4d3e4141  <=  ~I9c2da511df8277b7e61cf8611d04dd32 + 1;
                end else begin
                    Iad166146f7df5e8068fc6efe4d3e4141  <= I9c2da511df8277b7e61cf8611d04dd32 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Idd6a4f8ae94c431f2fa3312b4fd287ba != Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[3] ) begin
                    I4ac79b67a8904b95f7912d24af420585  <=  ~Ib8c628f3d97ffdf8a8b5db0fe90bbfa8 + 1;
                end else begin
                    I4ac79b67a8904b95f7912d24af420585  <= Ib8c628f3d97ffdf8a8b5db0fe90bbfa8 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Idd6a4f8ae94c431f2fa3312b4fd287ba != Iceb64ab2ff8a2e0dfdb74803811d4cfe[3] ) begin
                    I60ec7459bbe99fce295406bee1f2af46  <=  ~I42e0e42ae26723497a1da5e86e855499 + 1;
                end else begin
                    I60ec7459bbe99fce295406bee1f2af46  <= I42e0e42ae26723497a1da5e86e855499 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Idd6a4f8ae94c431f2fa3312b4fd287ba != I872f61d20baf011e867b44dc5539fc37[2] ) begin
                    I6fab46b1766878b26b53f352fee98223  <=  ~Id7e44a94fcaa2ca22ac9eb6756ecb830 + 1;
                end else begin
                    I6fab46b1766878b26b53f352fee98223  <= Id7e44a94fcaa2ca22ac9eb6756ecb830 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Idd6a4f8ae94c431f2fa3312b4fd287ba != Ida6059c6e0890f730536f97dfb83770b[0] ) begin
                    I36ca732e811d67cd742d24fd4cae887b  <=  ~Ie91db5e628b828dfaa8c1bd7d614d986 + 1;
                end else begin
                    I36ca732e811d67cd742d24fd4cae887b  <= Ie91db5e628b828dfaa8c1bd7d614d986 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9f1f8590dcf596097bc81001d51684b9 != Ib58043c04b5c4c86c1c67e57cc66dcf7[3] ) begin
                    I355725a804e0df68b4acf96ca98f2448  <=  ~I683ebfd7677d9e175d7a86479a5b42c6 + 1;
                end else begin
                    I355725a804e0df68b4acf96ca98f2448  <= I683ebfd7677d9e175d7a86479a5b42c6 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9f1f8590dcf596097bc81001d51684b9 != I5b7caaeb34c43e66e8d095a859e708fe[3] ) begin
                    I357137b41bb91e0659b1ac6ead9b5c12  <=  ~I11090ba16ce17a70438618b474837c33 + 1;
                end else begin
                    I357137b41bb91e0659b1ac6ead9b5c12  <= I11090ba16ce17a70438618b474837c33 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9f1f8590dcf596097bc81001d51684b9 != I6f5c991e5fdcf56d582c6f80eb6731df[2] ) begin
                    Ie3a336de822ac7baf8486b1618ef1126  <=  ~I845dd61995152e9d39cea7f0370b5a4d + 1;
                end else begin
                    Ie3a336de822ac7baf8486b1618ef1126  <= I845dd61995152e9d39cea7f0370b5a4d ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9f1f8590dcf596097bc81001d51684b9 != I1993c1ed200d7cdf838d23c72a0c1c0b[0] ) begin
                    I354fdd241d5d07f0d8380fe8924e0a8c  <=  ~Ia3e4dff8c98b38b6aebec9094ed26421 + 1;
                end else begin
                    I354fdd241d5d07f0d8380fe8924e0a8c  <= Ia3e4dff8c98b38b6aebec9094ed26421 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Icecd765baa87877675b0f3972d78c02f != Ibc0871b3c992fd278815fdbefcd2bac0[3] ) begin
                    I634484f00590216c0f74f975c9c83400  <=  ~Id69a54dc4854348a482f052c64a736ca + 1;
                end else begin
                    I634484f00590216c0f74f975c9c83400  <= Id69a54dc4854348a482f052c64a736ca ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Icecd765baa87877675b0f3972d78c02f != I61f0c04673dfb262ef6912eb2df39120[3] ) begin
                    Ia89da2f1890524ad3519ab403dd0686c  <=  ~I0f56c52253603ac01a22f3b942429262 + 1;
                end else begin
                    Ia89da2f1890524ad3519ab403dd0686c  <= I0f56c52253603ac01a22f3b942429262 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Icecd765baa87877675b0f3972d78c02f != Ia5cc3055ba3365e64cf59c4d4fd3f093[2] ) begin
                    Ib1357cb20f471f1670ac2448f964f8eb  <=  ~I718f82404f82fe0e822ee20d33ad20a2 + 1;
                end else begin
                    Ib1357cb20f471f1670ac2448f964f8eb  <= I718f82404f82fe0e822ee20d33ad20a2 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Icecd765baa87877675b0f3972d78c02f != I07e04e352df9aa1988ccf05d9cb2d1d7[0] ) begin
                    Id38b705f5d2863a020a475ffffc8afd6  <=  ~I6c86073aaa32b64a43d06eb1a2d9fba8 + 1;
                end else begin
                    Id38b705f5d2863a020a475ffffc8afd6  <= I6c86073aaa32b64a43d06eb1a2d9fba8 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I401a38ea1d71dcc71d17a4694ceb0988 != I8695e1e94cbfcbe4b9eae315b042529e[3] ) begin
                    I38c3e3e136acb79c8a0ff850bcc55f16  <=  ~Ie0c8e27167e6ba97a83dd238086f45e6 + 1;
                end else begin
                    I38c3e3e136acb79c8a0ff850bcc55f16  <= Ie0c8e27167e6ba97a83dd238086f45e6 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I401a38ea1d71dcc71d17a4694ceb0988 != Ibeb5edab51cd6aedad9c2ecedaded6f5[3] ) begin
                    Iedbe9d0e48bd36064f59faea51afddb9  <=  ~I6bb5e8ee16a2bc0c3b77c882cfb659e7 + 1;
                end else begin
                    Iedbe9d0e48bd36064f59faea51afddb9  <= I6bb5e8ee16a2bc0c3b77c882cfb659e7 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I401a38ea1d71dcc71d17a4694ceb0988 != Iea7da1f43ba202d753b0edb0be8b3fcf[2] ) begin
                    I6359856a1843d8c8b65dc478bccb3acd  <=  ~Ieef625ad664ddadc849be46d1c083748 + 1;
                end else begin
                    I6359856a1843d8c8b65dc478bccb3acd  <= Ieef625ad664ddadc849be46d1c083748 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I401a38ea1d71dcc71d17a4694ceb0988 != Ic4c0ebcc3711c9844a3aa3875483d2f7[0] ) begin
                    Id6e5d67e7bb7c4b999459374ea80459a  <=  ~Ice91b069200a91b2ad48fbf87bb2e766 + 1;
                end else begin
                    Id6e5d67e7bb7c4b999459374ea80459a  <= Ice91b069200a91b2ad48fbf87bb2e766 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I3db9b61e28a51e974e2d5e323ad53c1e != Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[4] ) begin
                    Iad44c932cfa5c249c5e59f8c706173a8  <=  ~I9d4c7c85b4da5f7003ff05ed3a240a2e + 1;
                end else begin
                    Iad44c932cfa5c249c5e59f8c706173a8  <= I9d4c7c85b4da5f7003ff05ed3a240a2e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I3db9b61e28a51e974e2d5e323ad53c1e != Ibeb5edab51cd6aedad9c2ecedaded6f5[4] ) begin
                    Ic3871325d57b310c95ca02fcaca529eb  <=  ~Ia8f1616f8a65025446a5ab4cc1624f9b + 1;
                end else begin
                    Ic3871325d57b310c95ca02fcaca529eb  <= Ia8f1616f8a65025446a5ab4cc1624f9b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I3db9b61e28a51e974e2d5e323ad53c1e != I50976b0051e84b6a42fc1dbabd7d20ae[2] ) begin
                    Ica1997c6c569c1d1f45224fbaa4e6b59  <=  ~I29848deb21ad480cdf155d849dc7bd48 + 1;
                end else begin
                    Ica1997c6c569c1d1f45224fbaa4e6b59  <= I29848deb21ad480cdf155d849dc7bd48 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I3db9b61e28a51e974e2d5e323ad53c1e != I02b62fafd371de339f299f8aefec6c43[2] ) begin
                    If9c12f8662333fb54a45cfa1bc5da487  <=  ~I1ae69988f89b200bd0e48f640211321c + 1;
                end else begin
                    If9c12f8662333fb54a45cfa1bc5da487  <= I1ae69988f89b200bd0e48f640211321c ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I3db9b61e28a51e974e2d5e323ad53c1e != I872f61d20baf011e867b44dc5539fc37[3] ) begin
                    Ieaf14683f40374c4531326d228cb43c3  <=  ~I7ddcc3c9f4d21aacc07d8eb285dee83e + 1;
                end else begin
                    Ieaf14683f40374c4531326d228cb43c3  <= I7ddcc3c9f4d21aacc07d8eb285dee83e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I3db9b61e28a51e974e2d5e323ad53c1e != I28e344560ba76bb3b76d01d8c53693a9[0] ) begin
                    I05341013abd4206eb66fcddfd63bfe26  <=  ~I28f7cf50ea7ac81667ff1353e0e121bd + 1;
                end else begin
                    I05341013abd4206eb66fcddfd63bfe26  <= I28f7cf50ea7ac81667ff1353e0e121bd ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I96d0a4387f9b959bc779ac13351182cc != Ib58043c04b5c4c86c1c67e57cc66dcf7[4] ) begin
                    I78212ae965ab2dcb2eed0b060d6b253f  <=  ~I09b7dd699ae0c4d34a7d1588efc90452 + 1;
                end else begin
                    I78212ae965ab2dcb2eed0b060d6b253f  <= I09b7dd699ae0c4d34a7d1588efc90452 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I96d0a4387f9b959bc779ac13351182cc != Iceb64ab2ff8a2e0dfdb74803811d4cfe[4] ) begin
                    I29ab844f80c105d247c5c15faa35863c  <=  ~Ic937101cc53e67403e56ac85011aa9ba + 1;
                end else begin
                    I29ab844f80c105d247c5c15faa35863c  <= Ic937101cc53e67403e56ac85011aa9ba ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I96d0a4387f9b959bc779ac13351182cc != I82e0e091fba6f79cef97eacac4b43ecb[2] ) begin
                    I7ef544597a185b1de63b4ffc4a1d44c2  <=  ~Ib42b03d2f76b8939ff3183008b17a969 + 1;
                end else begin
                    I7ef544597a185b1de63b4ffc4a1d44c2  <= Ib42b03d2f76b8939ff3183008b17a969 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I96d0a4387f9b959bc779ac13351182cc != I0e0b15868b02ca52b260f17f150d237e[2] ) begin
                    I27fd0073dbcdee599fbe85cf48806efc  <=  ~I4b99f00b1c2cdcee6bf4f1d2e8199ee4 + 1;
                end else begin
                    I27fd0073dbcdee599fbe85cf48806efc  <= I4b99f00b1c2cdcee6bf4f1d2e8199ee4 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I96d0a4387f9b959bc779ac13351182cc != I6f5c991e5fdcf56d582c6f80eb6731df[3] ) begin
                    I5fc3c26d6c5aa893dfd5caa0f677233a  <=  ~I01e153b020e1349eb66b47de581408df + 1;
                end else begin
                    I5fc3c26d6c5aa893dfd5caa0f677233a  <= I01e153b020e1349eb66b47de581408df ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I96d0a4387f9b959bc779ac13351182cc != I0600def6e6caada88ba6dedbb0d322ac[0] ) begin
                    I15da71a21f5842cb65b543d9bc3e267b  <=  ~I8ca1a48206ed8f1dc7ca57d77d0331a2 + 1;
                end else begin
                    I15da71a21f5842cb65b543d9bc3e267b  <= I8ca1a48206ed8f1dc7ca57d77d0331a2 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I64082bc75fdbeb69a52a4361ed2d5883 != Ibc0871b3c992fd278815fdbefcd2bac0[4] ) begin
                    Ib3b1db2d8b669988c887ed780e439b26  <=  ~I40e8430f50206db37e500c22f461b0c7 + 1;
                end else begin
                    Ib3b1db2d8b669988c887ed780e439b26  <= I40e8430f50206db37e500c22f461b0c7 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I64082bc75fdbeb69a52a4361ed2d5883 != I5b7caaeb34c43e66e8d095a859e708fe[4] ) begin
                    I5d70bc64cf7b3d3ef4180e082e533237  <=  ~I521128b7d945e025ded04037494c850a + 1;
                end else begin
                    I5d70bc64cf7b3d3ef4180e082e533237  <= I521128b7d945e025ded04037494c850a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I64082bc75fdbeb69a52a4361ed2d5883 != I04302edb2671c5bc0ca2673cd53935e1[2] ) begin
                    I6354a0e638340378124e4df7f3d145b8  <=  ~Ic24dbb1a30bb9a32c1992afcba90d4fb + 1;
                end else begin
                    I6354a0e638340378124e4df7f3d145b8  <= Ic24dbb1a30bb9a32c1992afcba90d4fb ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I64082bc75fdbeb69a52a4361ed2d5883 != I3c0b6f53f0a5cda5b6758b2ee2c83b92[2] ) begin
                    I438522d92cce6f7010246424746ca255  <=  ~I06cc903106b42e397fa7c4bc6c5edea4 + 1;
                end else begin
                    I438522d92cce6f7010246424746ca255  <= I06cc903106b42e397fa7c4bc6c5edea4 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I64082bc75fdbeb69a52a4361ed2d5883 != Ia5cc3055ba3365e64cf59c4d4fd3f093[3] ) begin
                    Iab953a8974a1eb619dc0f074c003b5f9  <=  ~I765dff22de01d419a6626919d23850f2 + 1;
                end else begin
                    Iab953a8974a1eb619dc0f074c003b5f9  <= I765dff22de01d419a6626919d23850f2 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I64082bc75fdbeb69a52a4361ed2d5883 != Iddbf50612c89b5b95a5c9efb5575cae3[0] ) begin
                    Iccf255fb3422c558465e45226068a16d  <=  ~Ie9538b63a057a50371de2d17898d3ad7 + 1;
                end else begin
                    Iccf255fb3422c558465e45226068a16d  <= Ie9538b63a057a50371de2d17898d3ad7 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I62929057b7c214bd38fd532e20ba5623 != I8695e1e94cbfcbe4b9eae315b042529e[4] ) begin
                    I35b2c7e9cdc53a98913e1c16a3a47b37  <=  ~If93a5596528db9017b8783fa0cf1dbc2 + 1;
                end else begin
                    I35b2c7e9cdc53a98913e1c16a3a47b37  <= If93a5596528db9017b8783fa0cf1dbc2 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I62929057b7c214bd38fd532e20ba5623 != I61f0c04673dfb262ef6912eb2df39120[4] ) begin
                    Ie33a780b0221084898c9fc5b237b244a  <=  ~I68016caaf170fbe2734c5b6aaf089894 + 1;
                end else begin
                    Ie33a780b0221084898c9fc5b237b244a  <= I68016caaf170fbe2734c5b6aaf089894 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I62929057b7c214bd38fd532e20ba5623 != I480a0f6d6c3eb936de10a72749f6cd3f[2] ) begin
                    I9590eb28a81c730b83b92ef7653e71a1  <=  ~I169b0fac6d01a713986b636bf8dfc3fb + 1;
                end else begin
                    I9590eb28a81c730b83b92ef7653e71a1  <= I169b0fac6d01a713986b636bf8dfc3fb ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I62929057b7c214bd38fd532e20ba5623 != I8e591d83170c8ba46d31c61935311b22[2] ) begin
                    Ib8bf21f32c0e8b9cfa42a53807bfe3a3  <=  ~Iddb14d68b464d04fe9e0b4e62789601a + 1;
                end else begin
                    Ib8bf21f32c0e8b9cfa42a53807bfe3a3  <= Iddb14d68b464d04fe9e0b4e62789601a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I62929057b7c214bd38fd532e20ba5623 != Iea7da1f43ba202d753b0edb0be8b3fcf[3] ) begin
                    If6f3d91c3c7a43622b9a522492cd83d3  <=  ~Ie5b71f77beb734a6ab7f7be6c6f9c252 + 1;
                end else begin
                    If6f3d91c3c7a43622b9a522492cd83d3  <= Ie5b71f77beb734a6ab7f7be6c6f9c252 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I62929057b7c214bd38fd532e20ba5623 != Iadc8f7f87b50bfff53d2d12d82489829[0] ) begin
                    I1c2674b2e6b269ed539827412c5199a5  <=  ~I59f9fa0b81ca88915c338ece1d1e08d5 + 1;
                end else begin
                    I1c2674b2e6b269ed539827412c5199a5  <= I59f9fa0b81ca88915c338ece1d1e08d5 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I641179f37fef63e7deec603b3291381c != Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[5] ) begin
                    I10f14b6433498e3b9e9bf021b60115e8  <=  ~I4f27922ccb21b65dcfe2dc0fcc97cdf3 + 1;
                end else begin
                    I10f14b6433498e3b9e9bf021b60115e8  <= I4f27922ccb21b65dcfe2dc0fcc97cdf3 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I641179f37fef63e7deec603b3291381c != I04302edb2671c5bc0ca2673cd53935e1[3] ) begin
                    I0236c912c6d684bf4862b725be9d5951  <=  ~Idd7ae55ba748fb36e49684037212936d + 1;
                end else begin
                    I0236c912c6d684bf4862b725be9d5951  <= Idd7ae55ba748fb36e49684037212936d ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I641179f37fef63e7deec603b3291381c != I3c0b6f53f0a5cda5b6758b2ee2c83b92[3] ) begin
                    I92496f68b44a94565af28a2c28d6fbae  <=  ~Ib8da505d1572487e814e7b0682e6dfa9 + 1;
                end else begin
                    I92496f68b44a94565af28a2c28d6fbae  <= Ib8da505d1572487e814e7b0682e6dfa9 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I641179f37fef63e7deec603b3291381c != I07930a807994815de45864af579902c4[3] ) begin
                    I964e17c41a134c080e9c43412a514f3f  <=  ~Idedb59a6fa2f6ad049f81ac652c645d8 + 1;
                end else begin
                    I964e17c41a134c080e9c43412a514f3f  <= Idedb59a6fa2f6ad049f81ac652c645d8 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I641179f37fef63e7deec603b3291381c != Iea7da1f43ba202d753b0edb0be8b3fcf[4] ) begin
                    Id023a6298e65da1f4da3831f5136afc2  <=  ~I7d50b49718ab2007accda67ac77a65d0 + 1;
                end else begin
                    Id023a6298e65da1f4da3831f5136afc2  <= I7d50b49718ab2007accda67ac77a65d0 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I641179f37fef63e7deec603b3291381c != I53a658b443200b9f11f1830547b5f42d[0] ) begin
                    I6a3f405bb4a0c4448d9b9d3dd95d036c  <=  ~I27e0600689451a7475a36143f0eb1079 + 1;
                end else begin
                    I6a3f405bb4a0c4448d9b9d3dd95d036c  <= I27e0600689451a7475a36143f0eb1079 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iff04b7ec87148f5bd408b4ec4b0590a5 != Ib58043c04b5c4c86c1c67e57cc66dcf7[5] ) begin
                    I0b56aa7a1b7549c91dddd3a06ecbaacf  <=  ~Iba6724b61ecb74552b9bb3cab96480c6 + 1;
                end else begin
                    I0b56aa7a1b7549c91dddd3a06ecbaacf  <= Iba6724b61ecb74552b9bb3cab96480c6 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iff04b7ec87148f5bd408b4ec4b0590a5 != I480a0f6d6c3eb936de10a72749f6cd3f[3] ) begin
                    I2ba1acca919bddcc22a41a28d43a4e3e  <=  ~I0abb44bd896fbc695e880fee67fb0c42 + 1;
                end else begin
                    I2ba1acca919bddcc22a41a28d43a4e3e  <= I0abb44bd896fbc695e880fee67fb0c42 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iff04b7ec87148f5bd408b4ec4b0590a5 != I8e591d83170c8ba46d31c61935311b22[3] ) begin
                    I7208256bb198bfce1be71390b01bc028  <=  ~Ifd714548110aa979e735cc6e13d3ef57 + 1;
                end else begin
                    I7208256bb198bfce1be71390b01bc028  <= Ifd714548110aa979e735cc6e13d3ef57 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iff04b7ec87148f5bd408b4ec4b0590a5 != I72a2f42b727a0503d43332c0f22d5ae3[3] ) begin
                    I9015033ab0caf3fa41dae4de43f24a82  <=  ~Ieeb6c7cdf1379ee3d2933d81bc812dbc + 1;
                end else begin
                    I9015033ab0caf3fa41dae4de43f24a82  <= Ieeb6c7cdf1379ee3d2933d81bc812dbc ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iff04b7ec87148f5bd408b4ec4b0590a5 != I872f61d20baf011e867b44dc5539fc37[4] ) begin
                    I5149125aaaad943d891df6a3c2be93a0  <=  ~Id682af5250edce8e3811d418ecf2dd10 + 1;
                end else begin
                    I5149125aaaad943d891df6a3c2be93a0  <= Id682af5250edce8e3811d418ecf2dd10 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iff04b7ec87148f5bd408b4ec4b0590a5 != I170f424df45651abe215ec74d649a9eb[0] ) begin
                    Ib528bb7a64cce4f694081d151fa6fa86  <=  ~I1d02127e28fb2e9aaf352815627960e7 + 1;
                end else begin
                    Ib528bb7a64cce4f694081d151fa6fa86  <= I1d02127e28fb2e9aaf352815627960e7 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I198bfb18d6f91c8f62777e6f592a88fa != Ibc0871b3c992fd278815fdbefcd2bac0[5] ) begin
                    I735db8b0ee0ec98e4cce0030b11508da  <=  ~Ibee34260749dc92b8523e83cd64d6a40 + 1;
                end else begin
                    I735db8b0ee0ec98e4cce0030b11508da  <= Ibee34260749dc92b8523e83cd64d6a40 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I198bfb18d6f91c8f62777e6f592a88fa != I50976b0051e84b6a42fc1dbabd7d20ae[3] ) begin
                    Iaf08bcaaeb15bb0c971432f7f8b16d0a  <=  ~Ie9a2a59c7b3571194198dca0c679c5f6 + 1;
                end else begin
                    Iaf08bcaaeb15bb0c971432f7f8b16d0a  <= Ie9a2a59c7b3571194198dca0c679c5f6 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I198bfb18d6f91c8f62777e6f592a88fa != I02b62fafd371de339f299f8aefec6c43[3] ) begin
                    Ie1681d905517daafcc7584725cd6014c  <=  ~Ie4b5a941feb385e88498a98e5f8ddc01 + 1;
                end else begin
                    Ie1681d905517daafcc7584725cd6014c  <= Ie4b5a941feb385e88498a98e5f8ddc01 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I198bfb18d6f91c8f62777e6f592a88fa != I8b8b9c4777e6df3eb2b9313e69ef2c8c[3] ) begin
                    Ice73589836da9028def6efb24a04dbbd  <=  ~I30b2b34a0cecfdbdeecba5f286befccd + 1;
                end else begin
                    Ice73589836da9028def6efb24a04dbbd  <= I30b2b34a0cecfdbdeecba5f286befccd ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I198bfb18d6f91c8f62777e6f592a88fa != I6f5c991e5fdcf56d582c6f80eb6731df[4] ) begin
                    Ie22b94121b58f17af14c75bfb27f96dd  <=  ~I8ce739ddc344cacb2de7f2c88a882170 + 1;
                end else begin
                    Ie22b94121b58f17af14c75bfb27f96dd  <= I8ce739ddc344cacb2de7f2c88a882170 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I198bfb18d6f91c8f62777e6f592a88fa != I3c897bfed190017a876c44fd73a7ecea[0] ) begin
                    Iaa40bd3abf668a21e0f87c7bda7b3f69  <=  ~I8b00260bb93e928e66e9d4aaeb0d9b55 + 1;
                end else begin
                    Iaa40bd3abf668a21e0f87c7bda7b3f69  <= I8b00260bb93e928e66e9d4aaeb0d9b55 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ia1562c88b4f56d8935c3a5d6ead0f816 != I8695e1e94cbfcbe4b9eae315b042529e[5] ) begin
                    Ib1a2b31d49ae476e2f1fb9acba2d5af0  <=  ~I9c1ca916654bad308af37d040b486cf8 + 1;
                end else begin
                    Ib1a2b31d49ae476e2f1fb9acba2d5af0  <= I9c1ca916654bad308af37d040b486cf8 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ia1562c88b4f56d8935c3a5d6ead0f816 != I82e0e091fba6f79cef97eacac4b43ecb[3] ) begin
                    Iadeedf3870f0b1eae98d0f7dbbeff04a  <=  ~I05749703a8a131453c563ed2264680a7 + 1;
                end else begin
                    Iadeedf3870f0b1eae98d0f7dbbeff04a  <= I05749703a8a131453c563ed2264680a7 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ia1562c88b4f56d8935c3a5d6ead0f816 != I0e0b15868b02ca52b260f17f150d237e[3] ) begin
                    Iaee6d725a8b2653eeac6d5acb91f8f36  <=  ~I4b76fe5f9863a41733b76decf9867d16 + 1;
                end else begin
                    Iaee6d725a8b2653eeac6d5acb91f8f36  <= I4b76fe5f9863a41733b76decf9867d16 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ia1562c88b4f56d8935c3a5d6ead0f816 != I4a16e8e7946d9a8220304fc1be3fb362[3] ) begin
                    Ide604e9bbe35cb55892a4602e18b2527  <=  ~I2805bb16fd574a64de548b39a532cd8a + 1;
                end else begin
                    Ide604e9bbe35cb55892a4602e18b2527  <= I2805bb16fd574a64de548b39a532cd8a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ia1562c88b4f56d8935c3a5d6ead0f816 != Ia5cc3055ba3365e64cf59c4d4fd3f093[4] ) begin
                    I6e37582849c2c98fd15ad92d22c222da  <=  ~Ide6a696c06f17f455d56bb28cad98bd0 + 1;
                end else begin
                    I6e37582849c2c98fd15ad92d22c222da  <= Ide6a696c06f17f455d56bb28cad98bd0 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ia1562c88b4f56d8935c3a5d6ead0f816 != Iaecbbae967be2c62cacf2fa7f9801899[0] ) begin
                    I919d36a7f6ad42c4bbc23222beb73106  <=  ~I39bce1f71ede4663c187ddfd6501eda1 + 1;
                end else begin
                    I919d36a7f6ad42c4bbc23222beb73106  <= I39bce1f71ede4663c187ddfd6501eda1 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iaccba3030d9d9f8a56f86d6e34ed6325 != Ibeb5edab51cd6aedad9c2ecedaded6f5[5] ) begin
                    I42f9b1f8ef24ad56c10086852678b456  <=  ~Id0e769bee61ae0a90c167fab061f5965 + 1;
                end else begin
                    I42f9b1f8ef24ad56c10086852678b456  <= Id0e769bee61ae0a90c167fab061f5965 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iaccba3030d9d9f8a56f86d6e34ed6325 != I82e0e091fba6f79cef97eacac4b43ecb[4] ) begin
                    I70ae07db9b44d530be220f06401d3d3d  <=  ~I83e03af8657a4a237641a9da7922e502 + 1;
                end else begin
                    I70ae07db9b44d530be220f06401d3d3d  <= I83e03af8657a4a237641a9da7922e502 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iaccba3030d9d9f8a56f86d6e34ed6325 != I0e0b15868b02ca52b260f17f150d237e[4] ) begin
                    I4afdeba4fc2a12a6cbe3567a519367fc  <=  ~I7565e071282ca6e77bb469afc522f1a2 + 1;
                end else begin
                    I4afdeba4fc2a12a6cbe3567a519367fc  <= I7565e071282ca6e77bb469afc522f1a2 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iaccba3030d9d9f8a56f86d6e34ed6325 != I872f61d20baf011e867b44dc5539fc37[5] ) begin
                    I770dff588ee1f52f58bea1921cb23383  <=  ~I5d0dc5d40385ab67bc7f540f212b6a97 + 1;
                end else begin
                    I770dff588ee1f52f58bea1921cb23383  <= I5d0dc5d40385ab67bc7f540f212b6a97 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iaccba3030d9d9f8a56f86d6e34ed6325 != I4267622319ca65909a3b40484dc74d3a[2] ) begin
                    I140078292f7209eccacd53a8bab18016  <=  ~I548cac395730b8386670cc4c7a64319a + 1;
                end else begin
                    I140078292f7209eccacd53a8bab18016  <= I548cac395730b8386670cc4c7a64319a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iaccba3030d9d9f8a56f86d6e34ed6325 != I52f867f1009f2e8d18b50a777942bde3[0] ) begin
                    I648d2a279dd1f587b1e45eeb35f2fa90  <=  ~Ic6d9bbbfb7890540edd10aa5758b0c4b + 1;
                end else begin
                    I648d2a279dd1f587b1e45eeb35f2fa90  <= Ic6d9bbbfb7890540edd10aa5758b0c4b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I953dfeeacee8c44c08d0a425fa549e49 != Iceb64ab2ff8a2e0dfdb74803811d4cfe[5] ) begin
                    I856fa68463aa5ef1ae53442699d38b33  <=  ~I7beb1f915a881a302f93c869d81417d1 + 1;
                end else begin
                    I856fa68463aa5ef1ae53442699d38b33  <= I7beb1f915a881a302f93c869d81417d1 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I953dfeeacee8c44c08d0a425fa549e49 != I04302edb2671c5bc0ca2673cd53935e1[4] ) begin
                    I6f3be51d69b2b64a04e55b8946d5dd56  <=  ~I5fc389bbc1ce31f7b326da719dc576d4 + 1;
                end else begin
                    I6f3be51d69b2b64a04e55b8946d5dd56  <= I5fc389bbc1ce31f7b326da719dc576d4 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I953dfeeacee8c44c08d0a425fa549e49 != I3c0b6f53f0a5cda5b6758b2ee2c83b92[4] ) begin
                    I66528f43f614f0edb715564eba3c77c1  <=  ~I922e6f05f7c6e0f6f0b1a5c9548df238 + 1;
                end else begin
                    I66528f43f614f0edb715564eba3c77c1  <= I922e6f05f7c6e0f6f0b1a5c9548df238 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I953dfeeacee8c44c08d0a425fa549e49 != I6f5c991e5fdcf56d582c6f80eb6731df[5] ) begin
                    I0d9f8c99194d9d6e187b4ad02fcce8b4  <=  ~I8c6bb234a1ca3deba637adf746672194 + 1;
                end else begin
                    I0d9f8c99194d9d6e187b4ad02fcce8b4  <= I8c6bb234a1ca3deba637adf746672194 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I953dfeeacee8c44c08d0a425fa549e49 != Iedd7d4ea8d082b40244c04946dfb14a0[2] ) begin
                    I74a4b9365391fd20c34588002ad40547  <=  ~Ide24ebd7423d4c4f43577b019f2e30e4 + 1;
                end else begin
                    I74a4b9365391fd20c34588002ad40547  <= Ide24ebd7423d4c4f43577b019f2e30e4 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I953dfeeacee8c44c08d0a425fa549e49 != I56a39a0c67b1de0a3cab6c61af3eebcf[0] ) begin
                    I194a64bef92ecf6714141eaa5d41c9d4  <=  ~Ifc412122eab7560c9021a17d7f8700c4 + 1;
                end else begin
                    I194a64bef92ecf6714141eaa5d41c9d4  <= Ifc412122eab7560c9021a17d7f8700c4 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I214a50bf9f879fe747904f4679fdd1f6 != I5b7caaeb34c43e66e8d095a859e708fe[5] ) begin
                    I7d9ad929660cd212387d893266b681da  <=  ~Ia5a56ed2c6b98e72002c6c5f946e7264 + 1;
                end else begin
                    I7d9ad929660cd212387d893266b681da  <= Ia5a56ed2c6b98e72002c6c5f946e7264 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I214a50bf9f879fe747904f4679fdd1f6 != I480a0f6d6c3eb936de10a72749f6cd3f[4] ) begin
                    I62d8efd4227cb3dc88aa08b6585fafc8  <=  ~Ia888ed8885f66084b777f66e25cef1e7 + 1;
                end else begin
                    I62d8efd4227cb3dc88aa08b6585fafc8  <= Ia888ed8885f66084b777f66e25cef1e7 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I214a50bf9f879fe747904f4679fdd1f6 != I8e591d83170c8ba46d31c61935311b22[4] ) begin
                    I49f2a06ceb3a59773c65b19f54ff362b  <=  ~I248229aecef00b87a70ce88920e407f5 + 1;
                end else begin
                    I49f2a06ceb3a59773c65b19f54ff362b  <= I248229aecef00b87a70ce88920e407f5 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I214a50bf9f879fe747904f4679fdd1f6 != Ia5cc3055ba3365e64cf59c4d4fd3f093[5] ) begin
                    If004de0cac6e5f7701a1fce48c6936d5  <=  ~I3d162a0ec918f220a7d5f4efdf89cb58 + 1;
                end else begin
                    If004de0cac6e5f7701a1fce48c6936d5  <= I3d162a0ec918f220a7d5f4efdf89cb58 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I214a50bf9f879fe747904f4679fdd1f6 != I56e1fe0c7a62589c123876f2b4e57a26[2] ) begin
                    I028ce03be0618b816e0ecdf43d4cd6e6  <=  ~I1ca0372f60e48f2f803778c9017023c0 + 1;
                end else begin
                    I028ce03be0618b816e0ecdf43d4cd6e6  <= I1ca0372f60e48f2f803778c9017023c0 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I214a50bf9f879fe747904f4679fdd1f6 != I490a65b3f7b30540906262ec5e12717b[0] ) begin
                    Id332e7f482524adeac7f7cdafcf5ca46  <=  ~Ieb9693d54f0808b0ba463fd3c316a80e + 1;
                end else begin
                    Id332e7f482524adeac7f7cdafcf5ca46  <= Ieb9693d54f0808b0ba463fd3c316a80e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ic88f2c344a8ad254fc7d7034cb594f6d != I61f0c04673dfb262ef6912eb2df39120[5] ) begin
                    Iabbd1668e0014df518ede5216232834c  <=  ~I63da03315d7e51fcacb0bc0298e506ed + 1;
                end else begin
                    Iabbd1668e0014df518ede5216232834c  <= I63da03315d7e51fcacb0bc0298e506ed ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ic88f2c344a8ad254fc7d7034cb594f6d != I50976b0051e84b6a42fc1dbabd7d20ae[4] ) begin
                    Idcb37cfc357cc088c775409fb9225b51  <=  ~I918f5a12e96bb96941f019940f27a5be + 1;
                end else begin
                    Idcb37cfc357cc088c775409fb9225b51  <= I918f5a12e96bb96941f019940f27a5be ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ic88f2c344a8ad254fc7d7034cb594f6d != I02b62fafd371de339f299f8aefec6c43[4] ) begin
                    I2ff3edcdb6158f1e3c9a555aeefc0850  <=  ~Ib4fb115f442ff544fa3d21b4e9d3f075 + 1;
                end else begin
                    I2ff3edcdb6158f1e3c9a555aeefc0850  <= Ib4fb115f442ff544fa3d21b4e9d3f075 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ic88f2c344a8ad254fc7d7034cb594f6d != Iea7da1f43ba202d753b0edb0be8b3fcf[5] ) begin
                    I6b24690f394792edb0d82b3b9e110851  <=  ~I387403482432a3196109484d1120d584 + 1;
                end else begin
                    I6b24690f394792edb0d82b3b9e110851  <= I387403482432a3196109484d1120d584 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ic88f2c344a8ad254fc7d7034cb594f6d != Ia8a468877c9f96713c8141df9205f92a[2] ) begin
                    I63e45abd4d27219bddcef06108b72021  <=  ~I619af17eaa4a56726d6ab322a74dd0a4 + 1;
                end else begin
                    I63e45abd4d27219bddcef06108b72021  <= I619af17eaa4a56726d6ab322a74dd0a4 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ic88f2c344a8ad254fc7d7034cb594f6d != Ib3c52fef8251d95e9abc8df0aad45d4e[0] ) begin
                    I226383d68f89db716cfd8d08b837865a  <=  ~I7a67ed3bb370520d0d25ce407ab8cd8b + 1;
                end else begin
                    I226383d68f89db716cfd8d08b837865a  <= I7a67ed3bb370520d0d25ce407ab8cd8b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (If299d1a4e044acbc70bc3b7bce9f86e9 != I8695e1e94cbfcbe4b9eae315b042529e[6] ) begin
                    Ic72f41f9bbf470aee3c9b9b8787b31c3  <=  ~I7629b35ca548190a81021a2c13d8919b + 1;
                end else begin
                    Ic72f41f9bbf470aee3c9b9b8787b31c3  <= I7629b35ca548190a81021a2c13d8919b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (If299d1a4e044acbc70bc3b7bce9f86e9 != Iceb64ab2ff8a2e0dfdb74803811d4cfe[6] ) begin
                    Ic3d00a27f15f8983a120395082854d6b  <=  ~I004851d3828f135ebe4d2e6ab83936bf + 1;
                end else begin
                    Ic3d00a27f15f8983a120395082854d6b  <= I004851d3828f135ebe4d2e6ab83936bf ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (If299d1a4e044acbc70bc3b7bce9f86e9 != Id6f07dee3e47f39e3b43329c26f690f7[2] ) begin
                    I19bba6a58ad3ef959b33701f82761984  <=  ~I0e2c382b2e62ed43b76697230e34b719 + 1;
                end else begin
                    I19bba6a58ad3ef959b33701f82761984  <= I0e2c382b2e62ed43b76697230e34b719 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (If299d1a4e044acbc70bc3b7bce9f86e9 != If75725e534dcb00364d73a42769539fb[0] ) begin
                    I2bdf5d319ba9089a4da34b108f5c5ae5  <=  ~I36dac27d10701db70fb2b5996a3f038f + 1;
                end else begin
                    I2bdf5d319ba9089a4da34b108f5c5ae5  <= I36dac27d10701db70fb2b5996a3f038f ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Idb373d2cf788f6a93a0e5df7f9179292 != Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[6] ) begin
                    I96008f47b9f134c9c4274cfcfb28e550  <=  ~I51d62ebd160eb0d073a7efb64d20079a + 1;
                end else begin
                    I96008f47b9f134c9c4274cfcfb28e550  <= I51d62ebd160eb0d073a7efb64d20079a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Idb373d2cf788f6a93a0e5df7f9179292 != I5b7caaeb34c43e66e8d095a859e708fe[6] ) begin
                    I34be4b353cf75603301372840c2f91c2  <=  ~Ib3545a88d68631af1c94ca2cb1f379af + 1;
                end else begin
                    I34be4b353cf75603301372840c2f91c2  <= Ib3545a88d68631af1c94ca2cb1f379af ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Idb373d2cf788f6a93a0e5df7f9179292 != Ic7f04c065f8ff82c2288f1de77d37189[2] ) begin
                    Iec71fe7fcebccf1ae0d10a5d187fcc44  <=  ~I81ad7b044118734f4dc32a1a4e8eba31 + 1;
                end else begin
                    Iec71fe7fcebccf1ae0d10a5d187fcc44  <= I81ad7b044118734f4dc32a1a4e8eba31 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Idb373d2cf788f6a93a0e5df7f9179292 != I9ddc427eef437ecc3ac4a2cf52aad4c3[0] ) begin
                    Ia91800792941ec7cc60415c3f844e4ed  <=  ~I5ad8c235d46349b6d310d0f175f84288 + 1;
                end else begin
                    Ia91800792941ec7cc60415c3f844e4ed  <= I5ad8c235d46349b6d310d0f175f84288 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ic73b8c8f76a985330d4ac1fa0cc28e7f != Ib58043c04b5c4c86c1c67e57cc66dcf7[6] ) begin
                    I71412803cc5229025487255aec62ec4f  <=  ~Ibc00920378e2427df2a63a47dc3eaded + 1;
                end else begin
                    I71412803cc5229025487255aec62ec4f  <= Ibc00920378e2427df2a63a47dc3eaded ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ic73b8c8f76a985330d4ac1fa0cc28e7f != I61f0c04673dfb262ef6912eb2df39120[6] ) begin
                    Ibd89458312687610aa166a9538968851  <=  ~Ic5195bbaa69d95059cca6e152dc9f705 + 1;
                end else begin
                    Ibd89458312687610aa166a9538968851  <= Ic5195bbaa69d95059cca6e152dc9f705 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ic73b8c8f76a985330d4ac1fa0cc28e7f != Ieb244944e7ee8236a207924f56fbc689[2] ) begin
                    I1c3c4ce44610e04c5eef2fcbc2ea5114  <=  ~Ia01f20e0bcf35c2ee4963e9c392c1004 + 1;
                end else begin
                    I1c3c4ce44610e04c5eef2fcbc2ea5114  <= Ia01f20e0bcf35c2ee4963e9c392c1004 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ic73b8c8f76a985330d4ac1fa0cc28e7f != I8999ca1f2fe9d4a30bd38fcb0daad2a4[0] ) begin
                    Id7c507d96098ee7a955af8a48ee5d72a  <=  ~I9f6f48fea88d1cd73ef2b24c7e819964 + 1;
                end else begin
                    Id7c507d96098ee7a955af8a48ee5d72a  <= I9f6f48fea88d1cd73ef2b24c7e819964 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I134dfb2c57d8cdffd2789e2f442c3247 != Ibc0871b3c992fd278815fdbefcd2bac0[6] ) begin
                    If1607e907e626902ee26d15020a64c21  <=  ~I847feea780cc8a06caea2d2ea79ad281 + 1;
                end else begin
                    If1607e907e626902ee26d15020a64c21  <= I847feea780cc8a06caea2d2ea79ad281 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I134dfb2c57d8cdffd2789e2f442c3247 != Ibeb5edab51cd6aedad9c2ecedaded6f5[6] ) begin
                    I3ed5d0fca86f35b3d4b4a89c6147d0cd  <=  ~I7ef6f4aeda7fd6775839c068c681f9bc + 1;
                end else begin
                    I3ed5d0fca86f35b3d4b4a89c6147d0cd  <= I7ef6f4aeda7fd6775839c068c681f9bc ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I134dfb2c57d8cdffd2789e2f442c3247 != Ie9b2be4c32334220e134e041ca8dfc06[2] ) begin
                    I599d01cfe6e54d8e45d64446c446818d  <=  ~I0645e741da20a4957747188273a655b1 + 1;
                end else begin
                    I599d01cfe6e54d8e45d64446c446818d  <= I0645e741da20a4957747188273a655b1 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I134dfb2c57d8cdffd2789e2f442c3247 != Ie11cf6677812bb739255b053a9c9cd56[0] ) begin
                    Ie15e4c1bcdb0e18085d4b320ac6a925c  <=  ~I71125dffdd2d37e44dbb46143c1e8d9a + 1;
                end else begin
                    Ie15e4c1bcdb0e18085d4b320ac6a925c  <= I71125dffdd2d37e44dbb46143c1e8d9a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I0c735e43be8030078ec10bdb6882e79c != I5b7caaeb34c43e66e8d095a859e708fe[7] ) begin
                    I14834fc8e6489775359bcecf5a37ff4d  <=  ~I50c166f958b22ce866cd40334918274c + 1;
                end else begin
                    I14834fc8e6489775359bcecf5a37ff4d  <= I50c166f958b22ce866cd40334918274c ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I0c735e43be8030078ec10bdb6882e79c != I2fbf89398a148c47810456812dbee5a6[3] ) begin
                    Ic87c3d7762a18772972552162e1d1a8c  <=  ~Icd225144fd331b870847044b4d02bed0 + 1;
                end else begin
                    Ic87c3d7762a18772972552162e1d1a8c  <= Icd225144fd331b870847044b4d02bed0 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I0c735e43be8030078ec10bdb6882e79c != If79ed5ee2b8710da0608c1e245d07d55[3] ) begin
                    I157fdf8775206858c08682db3039b084  <=  ~I5e876482090ce6007c2a2f2101c24654 + 1;
                end else begin
                    I157fdf8775206858c08682db3039b084  <= I5e876482090ce6007c2a2f2101c24654 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I0c735e43be8030078ec10bdb6882e79c != I872f61d20baf011e867b44dc5539fc37[6] ) begin
                    I8f0a90e761111a613d2488285534a500  <=  ~I026ded06f56d9ca93f47fd85aec4f7ad + 1;
                end else begin
                    I8f0a90e761111a613d2488285534a500  <= I026ded06f56d9ca93f47fd85aec4f7ad ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I0c735e43be8030078ec10bdb6882e79c != Iacc1d5a5c7811f0c9326ef80d1154fbb[0] ) begin
                    I5485d9edcafc6202f6e5f0969979802f  <=  ~Iec596e94ec168a564bccbbaa7df833c9 + 1;
                end else begin
                    I5485d9edcafc6202f6e5f0969979802f  <= Iec596e94ec168a564bccbbaa7df833c9 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie9951415c1d599570af1787767caa2dc != I61f0c04673dfb262ef6912eb2df39120[7] ) begin
                    Icbaf92a8e9875bcb19a1d074779a9ea5  <=  ~Ib514e01c261e43a725582a10596eed32 + 1;
                end else begin
                    Icbaf92a8e9875bcb19a1d074779a9ea5  <= Ib514e01c261e43a725582a10596eed32 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie9951415c1d599570af1787767caa2dc != Icac5a9001ee113e612e3457b4b49ee68[3] ) begin
                    I20c2057240417146df144b518b43d052  <=  ~Ic19a62cdecb2329370f7e11c48d3738d + 1;
                end else begin
                    I20c2057240417146df144b518b43d052  <= Ic19a62cdecb2329370f7e11c48d3738d ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie9951415c1d599570af1787767caa2dc != I9497bbb4f746969a95cff948a3ee9ade[3] ) begin
                    Ia30539545e66c4cfc16828140149180a  <=  ~Ib2f5691baa59adfbaad62f6ffc71fb05 + 1;
                end else begin
                    Ia30539545e66c4cfc16828140149180a  <= Ib2f5691baa59adfbaad62f6ffc71fb05 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie9951415c1d599570af1787767caa2dc != I6f5c991e5fdcf56d582c6f80eb6731df[6] ) begin
                    I71e101962e766a4d1484b3235359a4b5  <=  ~I9bdfaca6112385deb86e24ad7e45bbaa + 1;
                end else begin
                    I71e101962e766a4d1484b3235359a4b5  <= I9bdfaca6112385deb86e24ad7e45bbaa ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie9951415c1d599570af1787767caa2dc != I0efdadfd49c035a49d92243391395bca[0] ) begin
                    I7fe364f9f537cbef782e7007848a1c10  <=  ~I0e647bb8351cfe7828423e7099525585 + 1;
                end else begin
                    I7fe364f9f537cbef782e7007848a1c10  <= I0e647bb8351cfe7828423e7099525585 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I2630f187d63ba9b0af52c77093e6b760 != Ibeb5edab51cd6aedad9c2ecedaded6f5[7] ) begin
                    Ib0126fb335e32793c400a97c5a4a337c  <=  ~I185b758fb3e50bcfb1464fe2ab593cfe + 1;
                end else begin
                    Ib0126fb335e32793c400a97c5a4a337c  <= I185b758fb3e50bcfb1464fe2ab593cfe ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I2630f187d63ba9b0af52c77093e6b760 != I9461e92a5880cb9e04fcece2ef4674f0[3] ) begin
                    I2993acb61f1abe529f8a60c94a438550  <=  ~Ie25e944f9e3100c39b69bb38dffca177 + 1;
                end else begin
                    I2993acb61f1abe529f8a60c94a438550  <= Ie25e944f9e3100c39b69bb38dffca177 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I2630f187d63ba9b0af52c77093e6b760 != I651d700a00d7004d8728bc7356f30926[3] ) begin
                    Ic3b4752136ac08e343933ccc3a4ec47c  <=  ~I8e77032a54376578b3d16799e30c97f7 + 1;
                end else begin
                    Ic3b4752136ac08e343933ccc3a4ec47c  <= I8e77032a54376578b3d16799e30c97f7 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I2630f187d63ba9b0af52c77093e6b760 != Ia5cc3055ba3365e64cf59c4d4fd3f093[6] ) begin
                    Ic1efa395cc1fd2c5a1d1559fb169a5a0  <=  ~I4cd2a7f8f8ec378200b00d03e447ac92 + 1;
                end else begin
                    Ic1efa395cc1fd2c5a1d1559fb169a5a0  <= I4cd2a7f8f8ec378200b00d03e447ac92 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I2630f187d63ba9b0af52c77093e6b760 != Ie34d59bc77e06807937fe6f6860527e9[0] ) begin
                    I52dcf5bace9cadcf8a895aaa6a8c1da8  <=  ~I1b3c55aca0da232cf3f81d6d0914729f + 1;
                end else begin
                    I52dcf5bace9cadcf8a895aaa6a8c1da8  <= I1b3c55aca0da232cf3f81d6d0914729f ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I83db667ace2f04ef4950e2c186e0e6a4 != Iceb64ab2ff8a2e0dfdb74803811d4cfe[7] ) begin
                    I6b1d01c3cb8fb51e43cdb788b89816be  <=  ~I34c76f1a126120c4474e750e9b51e034 + 1;
                end else begin
                    I6b1d01c3cb8fb51e43cdb788b89816be  <= I34c76f1a126120c4474e750e9b51e034 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I83db667ace2f04ef4950e2c186e0e6a4 != I6ebab438dc55ccf6c1600313891d9c38[3] ) begin
                    I33b99994abbb5ecf8eed4de39033e4f8  <=  ~I0edb624c344787066a2267757052196b + 1;
                end else begin
                    I33b99994abbb5ecf8eed4de39033e4f8  <= I0edb624c344787066a2267757052196b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I83db667ace2f04ef4950e2c186e0e6a4 != Ic2580cbeec8c11a19bd1e2ebc29d255e[3] ) begin
                    I39e6d3fb468aa40ea73535e81556ea65  <=  ~Ia8443f199838742595ac114f35c00143 + 1;
                end else begin
                    I39e6d3fb468aa40ea73535e81556ea65  <= Ia8443f199838742595ac114f35c00143 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I83db667ace2f04ef4950e2c186e0e6a4 != Iea7da1f43ba202d753b0edb0be8b3fcf[6] ) begin
                    I5b55c285f7e3e78447fee68532ab9f7f  <=  ~Ib25b8a538c9d64880e114bf4a80ca42e + 1;
                end else begin
                    I5b55c285f7e3e78447fee68532ab9f7f  <= Ib25b8a538c9d64880e114bf4a80ca42e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I83db667ace2f04ef4950e2c186e0e6a4 != I9661cb126908d8550b585e2bad383bd6[0] ) begin
                    I13a9eec6175e695ab8bc4516cf57d6ec  <=  ~I25f6a3d7bb869082e4dbbd0ee8574c95 + 1;
                end else begin
                    I13a9eec6175e695ab8bc4516cf57d6ec  <= I25f6a3d7bb869082e4dbbd0ee8574c95 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie818c5ea3f3b879fded32e6cb06ca546 != Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[7] ) begin
                    Id0344146d1a53d418add6d2b185377dd  <=  ~If96057023747a1538d9f06966af48bc2 + 1;
                end else begin
                    Id0344146d1a53d418add6d2b185377dd  <= If96057023747a1538d9f06966af48bc2 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie818c5ea3f3b879fded32e6cb06ca546 != Ibeb5edab51cd6aedad9c2ecedaded6f5[8] ) begin
                    I20590d8fb97ec0b2164ffe17826136a7  <=  ~I199e995390462e06853b1f5cdbd46e0a + 1;
                end else begin
                    I20590d8fb97ec0b2164ffe17826136a7  <= I199e995390462e06853b1f5cdbd46e0a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie818c5ea3f3b879fded32e6cb06ca546 != I3d50cfeaa4b69c09bb648b8873a6bc24[3] ) begin
                    I05370777439b01811fe7f750d2f724f4  <=  ~Iec6325d585ddd0a9f86bb5cd0229960d + 1;
                end else begin
                    I05370777439b01811fe7f750d2f724f4  <= Iec6325d585ddd0a9f86bb5cd0229960d ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie818c5ea3f3b879fded32e6cb06ca546 != I3c0b6f53f0a5cda5b6758b2ee2c83b92[5] ) begin
                    I8cab9fba615b94fd4bb6934325be8ab8  <=  ~I4be1ccfec148a522fbf5b8375245cbb3 + 1;
                end else begin
                    I8cab9fba615b94fd4bb6934325be8ab8  <= I4be1ccfec148a522fbf5b8375245cbb3 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie818c5ea3f3b879fded32e6cb06ca546 != Ic0b832fbcbdb57745fefcc1ac1438808[0] ) begin
                    Iee73a7c685a4cee03f33d3ef379b1c8a  <=  ~I074386ff6a3d8d644f4b2501c69f26c7 + 1;
                end else begin
                    Iee73a7c685a4cee03f33d3ef379b1c8a  <= I074386ff6a3d8d644f4b2501c69f26c7 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I3a67a175863091a52844aae6ad277da0 != Ib58043c04b5c4c86c1c67e57cc66dcf7[7] ) begin
                    I32fcb28a27356bc6f403528836ea4c1f  <=  ~I83b378e5534c553b57beb22c5178a3ce + 1;
                end else begin
                    I32fcb28a27356bc6f403528836ea4c1f  <= I83b378e5534c553b57beb22c5178a3ce ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I3a67a175863091a52844aae6ad277da0 != Iceb64ab2ff8a2e0dfdb74803811d4cfe[8] ) begin
                    Ib74a56900c1f8b159ad381f61acee801  <=  ~I14f79d67f75af6a495d6eb2986210cda + 1;
                end else begin
                    Ib74a56900c1f8b159ad381f61acee801  <= I14f79d67f75af6a495d6eb2986210cda ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I3a67a175863091a52844aae6ad277da0 != I33a6ffad80ddf99a4d316a049078244d[3] ) begin
                    Ieb38fa62119a5a77c060d6634e051298  <=  ~Iacd805413ec1eb001b3083554f187554 + 1;
                end else begin
                    Ieb38fa62119a5a77c060d6634e051298  <= Iacd805413ec1eb001b3083554f187554 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I3a67a175863091a52844aae6ad277da0 != I8e591d83170c8ba46d31c61935311b22[5] ) begin
                    I86e495dc894d2aace15c1aff89798bf7  <=  ~I3e61e09fcc81a0011a79f5c5ce77bc46 + 1;
                end else begin
                    I86e495dc894d2aace15c1aff89798bf7  <= I3e61e09fcc81a0011a79f5c5ce77bc46 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I3a67a175863091a52844aae6ad277da0 != I2afd96714b26f30483c3935c2a68e64f[0] ) begin
                    I740dc91716e3906ad078e2c7cc3c925a  <=  ~I6e6cbb7dba8eb3c02b5b4e4469e23cea + 1;
                end else begin
                    I740dc91716e3906ad078e2c7cc3c925a  <= I6e6cbb7dba8eb3c02b5b4e4469e23cea ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ia3aba80aead67feab12e4800fef82322 != Ibc0871b3c992fd278815fdbefcd2bac0[7] ) begin
                    I081b38dbb37d4c14a6a9fd3fefa13daa  <=  ~I8b25822c33f7d506ef69216af3fdab44 + 1;
                end else begin
                    I081b38dbb37d4c14a6a9fd3fefa13daa  <= I8b25822c33f7d506ef69216af3fdab44 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ia3aba80aead67feab12e4800fef82322 != I5b7caaeb34c43e66e8d095a859e708fe[8] ) begin
                    I633a74e4dfa841c9fd13dbb6564c8493  <=  ~I06fd642cbc8aa2f65197801d7459cfa2 + 1;
                end else begin
                    I633a74e4dfa841c9fd13dbb6564c8493  <= I06fd642cbc8aa2f65197801d7459cfa2 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ia3aba80aead67feab12e4800fef82322 != I980165c1147ac5ff86619c841c6031dc[3] ) begin
                    I0b7b4c0a8503c751229edfe0237cc903  <=  ~I22202e6c3de9b06c04ce9514af28933e + 1;
                end else begin
                    I0b7b4c0a8503c751229edfe0237cc903  <= I22202e6c3de9b06c04ce9514af28933e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ia3aba80aead67feab12e4800fef82322 != I02b62fafd371de339f299f8aefec6c43[5] ) begin
                    I43b380be6df7df0d354223d0a0d6d6b6  <=  ~Ib991cdbb91133cb82e154c575e00a174 + 1;
                end else begin
                    I43b380be6df7df0d354223d0a0d6d6b6  <= Ib991cdbb91133cb82e154c575e00a174 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ia3aba80aead67feab12e4800fef82322 != Id6d4165b752630a1ce7ceb77fdcee477[0] ) begin
                    I514d2dc697e9b39ba027c418a6df6cb9  <=  ~I5590364df6874420e169aa444ab520b9 + 1;
                end else begin
                    I514d2dc697e9b39ba027c418a6df6cb9  <= I5590364df6874420e169aa444ab520b9 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I1181d42b560fca7bb5c924a81a5db1fc != I8695e1e94cbfcbe4b9eae315b042529e[7] ) begin
                    I3ea4c33a9419820ed54460eb64134dff  <=  ~I43a9e393037fb4aa84741dca22648459 + 1;
                end else begin
                    I3ea4c33a9419820ed54460eb64134dff  <= I43a9e393037fb4aa84741dca22648459 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I1181d42b560fca7bb5c924a81a5db1fc != I61f0c04673dfb262ef6912eb2df39120[8] ) begin
                    I80f3c8559da8e97bc5397bb8b621a0bd  <=  ~Ibb4d8301d90c66fdfac92b3fbc53c019 + 1;
                end else begin
                    I80f3c8559da8e97bc5397bb8b621a0bd  <= Ibb4d8301d90c66fdfac92b3fbc53c019 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I1181d42b560fca7bb5c924a81a5db1fc != I19df055705f322292a3601fa63f0e5f9[3] ) begin
                    Iaf4ae293c576af16f5f43a8b86c1aa3d  <=  ~Ibae217fa4b808e4accbeb8f4a9a976ab + 1;
                end else begin
                    Iaf4ae293c576af16f5f43a8b86c1aa3d  <= Ibae217fa4b808e4accbeb8f4a9a976ab ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I1181d42b560fca7bb5c924a81a5db1fc != I0e0b15868b02ca52b260f17f150d237e[5] ) begin
                    Ib42816335dd8475dcc78662c4c0786c1  <=  ~Ia8bd7a3594f7084a57e64da023bf784c + 1;
                end else begin
                    Ib42816335dd8475dcc78662c4c0786c1  <= Ia8bd7a3594f7084a57e64da023bf784c ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I1181d42b560fca7bb5c924a81a5db1fc != I59baaf1ad22721cde9064b8aad65ac76[0] ) begin
                    I782726e317a2aada9e755bcbc4b0d3fa  <=  ~I3ce4b9d41f5472bf60ed2802a2ab10eb + 1;
                end else begin
                    I782726e317a2aada9e755bcbc4b0d3fa  <= I3ce4b9d41f5472bf60ed2802a2ab10eb ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie4e5f3d7c5d2df30653f5666d14567bf != Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[8] ) begin
                    I1eede74f12d37331b399eb7136bc621f  <=  ~I93ec9bc6fbd056e7e52496546493e727 + 1;
                end else begin
                    I1eede74f12d37331b399eb7136bc621f  <= I93ec9bc6fbd056e7e52496546493e727 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie4e5f3d7c5d2df30653f5666d14567bf != I0e0b15868b02ca52b260f17f150d237e[6] ) begin
                    I343c9efe71164c01e9c7d599e032864a  <=  ~I2374b90dde1cf481baa40af31e1a43e3 + 1;
                end else begin
                    I343c9efe71164c01e9c7d599e032864a  <= I2374b90dde1cf481baa40af31e1a43e3 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie4e5f3d7c5d2df30653f5666d14567bf != I8b8b9c4777e6df3eb2b9313e69ef2c8c[4] ) begin
                    Idb72c046c5996fbbd80b706666ffbd92  <=  ~I0cee595f488a909ade8a3b4c90dbb0c7 + 1;
                end else begin
                    Idb72c046c5996fbbd80b706666ffbd92  <= I0cee595f488a909ade8a3b4c90dbb0c7 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie4e5f3d7c5d2df30653f5666d14567bf != I4267622319ca65909a3b40484dc74d3a[3] ) begin
                    I141fb1cbe09f9abe282cffd4de815d25  <=  ~Iba4c3d91d492b000ab1de7add9f171a9 + 1;
                end else begin
                    I141fb1cbe09f9abe282cffd4de815d25  <= Iba4c3d91d492b000ab1de7add9f171a9 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie4e5f3d7c5d2df30653f5666d14567bf != I9094f4e9c5b60add3acee212118a1dfa[0] ) begin
                    I11eb26cf0f0b3a334e8f7317bf8d9eb0  <=  ~I2b4152aa4c51cc1c1ffabac78cea267c + 1;
                end else begin
                    I11eb26cf0f0b3a334e8f7317bf8d9eb0  <= I2b4152aa4c51cc1c1ffabac78cea267c ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ifd9345cf219c58291c0b437aac093d78 != Ib58043c04b5c4c86c1c67e57cc66dcf7[8] ) begin
                    Iad354d876cb9fc72fc0143e6f7da9357  <=  ~Ie4c3dd5c191aff00a6d62006223c2b76 + 1;
                end else begin
                    Iad354d876cb9fc72fc0143e6f7da9357  <= Ie4c3dd5c191aff00a6d62006223c2b76 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ifd9345cf219c58291c0b437aac093d78 != I3c0b6f53f0a5cda5b6758b2ee2c83b92[6] ) begin
                    I92d9fec22d36b1baac8bd78abfc1bbd5  <=  ~Ie4c0ba9510f9b924999bb5f432137271 + 1;
                end else begin
                    I92d9fec22d36b1baac8bd78abfc1bbd5  <= Ie4c0ba9510f9b924999bb5f432137271 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ifd9345cf219c58291c0b437aac093d78 != I4a16e8e7946d9a8220304fc1be3fb362[4] ) begin
                    I262f2390e77ec486ccd3a6ed05816e2d  <=  ~I5bad544a17b384973d5672acbe0ac0d5 + 1;
                end else begin
                    I262f2390e77ec486ccd3a6ed05816e2d  <= I5bad544a17b384973d5672acbe0ac0d5 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ifd9345cf219c58291c0b437aac093d78 != Iedd7d4ea8d082b40244c04946dfb14a0[3] ) begin
                    I461195b7ae78743e09ee50486ad6ebe5  <=  ~I231bfb8e19e1d9c4bbd29a0bd75c1ed3 + 1;
                end else begin
                    I461195b7ae78743e09ee50486ad6ebe5  <= I231bfb8e19e1d9c4bbd29a0bd75c1ed3 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ifd9345cf219c58291c0b437aac093d78 != I13168bab2231ed22a3509142f990e408[0] ) begin
                    I26cb63ba20245b2c332b09e25c4409aa  <=  ~I1ecf87e33de04d02db9e64590bcaffde + 1;
                end else begin
                    I26cb63ba20245b2c332b09e25c4409aa  <= I1ecf87e33de04d02db9e64590bcaffde ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I4f2d7bb48918ce51efe6b3b12f9f8e65 != Ibc0871b3c992fd278815fdbefcd2bac0[8] ) begin
                    Ibac5e7b6d4bf5cd6926358318f0c418f  <=  ~I60c97bf58193f004e3fcfdbd6a03ce6e + 1;
                end else begin
                    Ibac5e7b6d4bf5cd6926358318f0c418f  <= I60c97bf58193f004e3fcfdbd6a03ce6e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I4f2d7bb48918ce51efe6b3b12f9f8e65 != I8e591d83170c8ba46d31c61935311b22[6] ) begin
                    I0d53bb5344cabe5fa5ce3ecf7122a260  <=  ~Ib71065a3fe70d3ab5f05b0c393278631 + 1;
                end else begin
                    I0d53bb5344cabe5fa5ce3ecf7122a260  <= Ib71065a3fe70d3ab5f05b0c393278631 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I4f2d7bb48918ce51efe6b3b12f9f8e65 != I07930a807994815de45864af579902c4[4] ) begin
                    I94f1724740defe5bb7e40041d0e266a0  <=  ~I984074a5c77445ad266463e20d77899e + 1;
                end else begin
                    I94f1724740defe5bb7e40041d0e266a0  <= I984074a5c77445ad266463e20d77899e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I4f2d7bb48918ce51efe6b3b12f9f8e65 != I56e1fe0c7a62589c123876f2b4e57a26[3] ) begin
                    I6ae2523095237282533e0b5f1c26b488  <=  ~I50bb40691aa09c42e0b64a076b50a971 + 1;
                end else begin
                    I6ae2523095237282533e0b5f1c26b488  <= I50bb40691aa09c42e0b64a076b50a971 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I4f2d7bb48918ce51efe6b3b12f9f8e65 != I280145f996e5e249788cacca7caf0095[0] ) begin
                    Idd7691d31f8d0c09ee988116d574ec59  <=  ~I753bff437b6c563f5fddf19685405504 + 1;
                end else begin
                    Idd7691d31f8d0c09ee988116d574ec59  <= I753bff437b6c563f5fddf19685405504 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ifa612e6208151c616c3a0319182a96f1 != I8695e1e94cbfcbe4b9eae315b042529e[8] ) begin
                    Ia0d940e16c8cbd4f7544f5a5cd7d83b2  <=  ~I21f2ec69bcc507756e2a5f85d3ead3e8 + 1;
                end else begin
                    Ia0d940e16c8cbd4f7544f5a5cd7d83b2  <= I21f2ec69bcc507756e2a5f85d3ead3e8 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ifa612e6208151c616c3a0319182a96f1 != I02b62fafd371de339f299f8aefec6c43[6] ) begin
                    I23eb1dc4d1c992f804dd04a2d823c778  <=  ~Iddec4486996054e475499d370016a685 + 1;
                end else begin
                    I23eb1dc4d1c992f804dd04a2d823c778  <= Iddec4486996054e475499d370016a685 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ifa612e6208151c616c3a0319182a96f1 != I72a2f42b727a0503d43332c0f22d5ae3[4] ) begin
                    Ia630e59cbce82a570ae3890a6c0221e5  <=  ~I3d3edd06f8907f4369b825062348da87 + 1;
                end else begin
                    Ia630e59cbce82a570ae3890a6c0221e5  <= I3d3edd06f8907f4369b825062348da87 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ifa612e6208151c616c3a0319182a96f1 != Ia8a468877c9f96713c8141df9205f92a[3] ) begin
                    Id1bacd13718f7c29c26b63c239d04dd8  <=  ~I72467ef10ecced8395a6870a39525787 + 1;
                end else begin
                    Id1bacd13718f7c29c26b63c239d04dd8  <= I72467ef10ecced8395a6870a39525787 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ifa612e6208151c616c3a0319182a96f1 != Ia9db6d176e9b9579a1aa5f257cd1a9f6[0] ) begin
                    Iecc02842a2d2b9b9e8187f2d39e62e05  <=  ~I9b74b672f55e7bf7560ba4dd2d0c79fd + 1;
                end else begin
                    Iecc02842a2d2b9b9e8187f2d39e62e05  <= I9b74b672f55e7bf7560ba4dd2d0c79fd ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9cb28a0cc6358610854c8f8d1dd3c707 != I5b7caaeb34c43e66e8d095a859e708fe[9] ) begin
                    I157bd468200e63385583b9045758d81e  <=  ~I285b012d2fb5e2279a79cf8edca24ac8 + 1;
                end else begin
                    I157bd468200e63385583b9045758d81e  <= I285b012d2fb5e2279a79cf8edca24ac8 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9cb28a0cc6358610854c8f8d1dd3c707 != I9c0b88a0be66d62f8ab061aeaee7e60f[3] ) begin
                    I09e9a3cd4c12d204f760758e873a177b  <=  ~I8faf911a7d1ea8b0abe54f6688068ca0 + 1;
                end else begin
                    I09e9a3cd4c12d204f760758e873a177b  <= I8faf911a7d1ea8b0abe54f6688068ca0 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9cb28a0cc6358610854c8f8d1dd3c707 != Iea7da1f43ba202d753b0edb0be8b3fcf[7] ) begin
                    I32701d9e4b96853c53f0ab651a6a4ba2  <=  ~I3dca974bf2d5631a47ebf8b945efab20 + 1;
                end else begin
                    I32701d9e4b96853c53f0ab651a6a4ba2  <= I3dca974bf2d5631a47ebf8b945efab20 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9cb28a0cc6358610854c8f8d1dd3c707 != I0ed43cf9eec83545457c57cfb6181d3c[0] ) begin
                    I5551342f1751fc64f32744a46b9649be  <=  ~I12141c45d147b058a9e392f3b7d7d06e + 1;
                end else begin
                    I5551342f1751fc64f32744a46b9649be  <= I12141c45d147b058a9e392f3b7d7d06e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I40bcc924f5cf1f7d587aa35267022261 != I61f0c04673dfb262ef6912eb2df39120[9] ) begin
                    I7a0eada108891aba06cecab5071232c9  <=  ~Ia527c96e30b782f837bc6206961400e4 + 1;
                end else begin
                    I7a0eada108891aba06cecab5071232c9  <= Ia527c96e30b782f837bc6206961400e4 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I40bcc924f5cf1f7d587aa35267022261 != Id88b9265ff08e0730e6a41abe1f80a32[3] ) begin
                    I4df3d4dac24877b14e6d361bafc1a800  <=  ~I6adbdb64422a08be9bf9e538db97463b + 1;
                end else begin
                    I4df3d4dac24877b14e6d361bafc1a800  <= I6adbdb64422a08be9bf9e538db97463b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I40bcc924f5cf1f7d587aa35267022261 != I872f61d20baf011e867b44dc5539fc37[7] ) begin
                    I765a8825e42180a6c63f7b33703bb483  <=  ~I958cdf5367c7b0bd58b70b763d3af8aa + 1;
                end else begin
                    I765a8825e42180a6c63f7b33703bb483  <= I958cdf5367c7b0bd58b70b763d3af8aa ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I40bcc924f5cf1f7d587aa35267022261 != I5b74f5fc705a0406ff2376cb8ac11db4[0] ) begin
                    Iff7c29299f005c1cd5a16b64601e727e  <=  ~I91b7b8e8887b5dd9853297463c55b78d + 1;
                end else begin
                    Iff7c29299f005c1cd5a16b64601e727e  <= I91b7b8e8887b5dd9853297463c55b78d ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I5238f7273b05b8b9f376314acdc6cc42 != Ibeb5edab51cd6aedad9c2ecedaded6f5[9] ) begin
                    I3c128efc9f80c9b8334bf7b61de71b43  <=  ~I6162978f0c57958ad0403246fb0530dd + 1;
                end else begin
                    I3c128efc9f80c9b8334bf7b61de71b43  <= I6162978f0c57958ad0403246fb0530dd ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I5238f7273b05b8b9f376314acdc6cc42 != I6330943c9295298c53e889d47c7904d9[3] ) begin
                    Ied00d87af99ae55144fdde41ebfc1357  <=  ~I508142e70fd04513977130556aa574ef + 1;
                end else begin
                    Ied00d87af99ae55144fdde41ebfc1357  <= I508142e70fd04513977130556aa574ef ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I5238f7273b05b8b9f376314acdc6cc42 != I6f5c991e5fdcf56d582c6f80eb6731df[7] ) begin
                    If2539da6722562bbf31786fd0036666a  <=  ~I2afab673e4b803ffd888f187de47fa49 + 1;
                end else begin
                    If2539da6722562bbf31786fd0036666a  <= I2afab673e4b803ffd888f187de47fa49 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I5238f7273b05b8b9f376314acdc6cc42 != I14f0d3ad4fec9ca492d6b36eb29a5dea[0] ) begin
                    I17a5446e942bcc1dc2c96930e0a87a70  <=  ~I7a56f81596920126a9ea2c9fb3a19285 + 1;
                end else begin
                    I17a5446e942bcc1dc2c96930e0a87a70  <= I7a56f81596920126a9ea2c9fb3a19285 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I7137f56eeb4c4ae08bbc238db4cd3441 != Iceb64ab2ff8a2e0dfdb74803811d4cfe[9] ) begin
                    Ia5eba52d169755c507b9e0094e467fab  <=  ~Ic6252de2c819f2243476ddf82e22d137 + 1;
                end else begin
                    Ia5eba52d169755c507b9e0094e467fab  <= Ic6252de2c819f2243476ddf82e22d137 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I7137f56eeb4c4ae08bbc238db4cd3441 != I5686b595177e07dd5bf231a35ee41659[3] ) begin
                    Ib9ceb8315f0cd848f861bab677c2c694  <=  ~Ieea8672b2f23711c6ba893de5c5d8bc2 + 1;
                end else begin
                    Ib9ceb8315f0cd848f861bab677c2c694  <= Ieea8672b2f23711c6ba893de5c5d8bc2 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I7137f56eeb4c4ae08bbc238db4cd3441 != Ia5cc3055ba3365e64cf59c4d4fd3f093[7] ) begin
                    I8e96c69e7d872be23229353808c34953  <=  ~I3a4dbdf517b8f9c93b567f91870e6160 + 1;
                end else begin
                    I8e96c69e7d872be23229353808c34953  <= I3a4dbdf517b8f9c93b567f91870e6160 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I7137f56eeb4c4ae08bbc238db4cd3441 != I3a25c80d9bf7655f4ce70cf29843db43[0] ) begin
                    I719b67f84e07e90dfd29a8cd5d94cf39  <=  ~I4731ee7a0e08c69e2bd2a8bcea0838c2 + 1;
                end else begin
                    I719b67f84e07e90dfd29a8cd5d94cf39  <= I4731ee7a0e08c69e2bd2a8bcea0838c2 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I02335be013799e2560a98b6a82a0c528 != Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[9] ) begin
                    I3e4754acc31d99bc71525789bdee0c1a  <=  ~I1b6cbbcf01a65cd1c2f1e241f849c904 + 1;
                end else begin
                    I3e4754acc31d99bc71525789bdee0c1a  <= I1b6cbbcf01a65cd1c2f1e241f849c904 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I02335be013799e2560a98b6a82a0c528 != Iceb64ab2ff8a2e0dfdb74803811d4cfe[10] ) begin
                    I0899e8fec1a7209cd94757c0b2f87c9a  <=  ~I663aee79f824c854f57c19e87207529b + 1;
                end else begin
                    I0899e8fec1a7209cd94757c0b2f87c9a  <= I663aee79f824c854f57c19e87207529b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I02335be013799e2560a98b6a82a0c528 != Icac5a9001ee113e612e3457b4b49ee68[4] ) begin
                    Ied029d0bdea3bf134744c99426fa72dc  <=  ~I34ff7299c9d83affa4512b7da302c199 + 1;
                end else begin
                    Ied029d0bdea3bf134744c99426fa72dc  <= I34ff7299c9d83affa4512b7da302c199 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I02335be013799e2560a98b6a82a0c528 != I56e1fe0c7a62589c123876f2b4e57a26[4] ) begin
                    I5aba6218461e8d571be03a3ef041ebaa  <=  ~I70ca6c9d0a5c99e0036479f7b5dd760a + 1;
                end else begin
                    I5aba6218461e8d571be03a3ef041ebaa  <= I70ca6c9d0a5c99e0036479f7b5dd760a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I02335be013799e2560a98b6a82a0c528 != I260dc9154b3a9fe38b0948e807bdb42d[0] ) begin
                    I2c835dfb3596b8bf057a7cc21122c81f  <=  ~I835bb7345787eaadc41816858e0a71a1 + 1;
                end else begin
                    I2c835dfb3596b8bf057a7cc21122c81f  <= I835bb7345787eaadc41816858e0a71a1 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Id327bb65156c8307901dfcb4184bb65f != Ib58043c04b5c4c86c1c67e57cc66dcf7[9] ) begin
                    If6e745bb85abba7282dae1f6f701225e  <=  ~I3c7f6fdd0e9cc7426df76027912d1ccb + 1;
                end else begin
                    If6e745bb85abba7282dae1f6f701225e  <= I3c7f6fdd0e9cc7426df76027912d1ccb ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Id327bb65156c8307901dfcb4184bb65f != I5b7caaeb34c43e66e8d095a859e708fe[10] ) begin
                    I918c46173eebc5b2a95e041cfd91d958  <=  ~I9ff512085174a7720705d0fb37c4ec34 + 1;
                end else begin
                    I918c46173eebc5b2a95e041cfd91d958  <= I9ff512085174a7720705d0fb37c4ec34 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Id327bb65156c8307901dfcb4184bb65f != I9461e92a5880cb9e04fcece2ef4674f0[4] ) begin
                    Ic8be2c94235fb40f78da33179ce4873a  <=  ~I6a69cdf2bae1ea68c9be56dcc4e76a59 + 1;
                end else begin
                    Ic8be2c94235fb40f78da33179ce4873a  <= I6a69cdf2bae1ea68c9be56dcc4e76a59 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Id327bb65156c8307901dfcb4184bb65f != Ia8a468877c9f96713c8141df9205f92a[4] ) begin
                    Ia3104c69fb4f7abfb5efa3874169a7ad  <=  ~I855ddead34ac131137ba644afbfea2b7 + 1;
                end else begin
                    Ia3104c69fb4f7abfb5efa3874169a7ad  <= I855ddead34ac131137ba644afbfea2b7 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Id327bb65156c8307901dfcb4184bb65f != Ic49b2c150e2face8c362e33f2d87f9c4[0] ) begin
                    Ib71b3d357c98dcdfae5c777ca3082275  <=  ~Ib1a463388daf270eb0ce698d7b5ded4b + 1;
                end else begin
                    Ib71b3d357c98dcdfae5c777ca3082275  <= Ib1a463388daf270eb0ce698d7b5ded4b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I56331cb7b310613016958553732cdf40 != Ibc0871b3c992fd278815fdbefcd2bac0[9] ) begin
                    Iadfc60386481092ae85cc148a2c40abb  <=  ~I74e4bb7530c02073f9b15a6389659d4b + 1;
                end else begin
                    Iadfc60386481092ae85cc148a2c40abb  <= I74e4bb7530c02073f9b15a6389659d4b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I56331cb7b310613016958553732cdf40 != I61f0c04673dfb262ef6912eb2df39120[10] ) begin
                    Ie21a2c9b22e7bf8425fb5c0f33e5f4f7  <=  ~I6721b13abeddc76139bdc7380434cc2a + 1;
                end else begin
                    Ie21a2c9b22e7bf8425fb5c0f33e5f4f7  <= I6721b13abeddc76139bdc7380434cc2a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I56331cb7b310613016958553732cdf40 != I6ebab438dc55ccf6c1600313891d9c38[4] ) begin
                    I7c3291f0250d13ca94802b0b071a95c6  <=  ~I84fba239c5705bcd92096e204cc9438c + 1;
                end else begin
                    I7c3291f0250d13ca94802b0b071a95c6  <= I84fba239c5705bcd92096e204cc9438c ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I56331cb7b310613016958553732cdf40 != I4267622319ca65909a3b40484dc74d3a[4] ) begin
                    If79d1d378f7c6fd29fc3335ec5f5c51d  <=  ~I4d46e4d50176768fda897949545e2125 + 1;
                end else begin
                    If79d1d378f7c6fd29fc3335ec5f5c51d  <= I4d46e4d50176768fda897949545e2125 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I56331cb7b310613016958553732cdf40 != I714350b3b56a3249aad06d5f59fbb291[0] ) begin
                    I086bf19f620c8a8f6888e775cb1ed7f4  <=  ~I57086cfab3b163c3911c3cf7bfb3141a + 1;
                end else begin
                    I086bf19f620c8a8f6888e775cb1ed7f4  <= I57086cfab3b163c3911c3cf7bfb3141a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie3b00960f8af88a5aba7a2104dfca9a7 != I8695e1e94cbfcbe4b9eae315b042529e[9] ) begin
                    I4a8abfa0896ce414d9b98093ef84455f  <=  ~Ice174debd5dc911fdf5d5756cff8d731 + 1;
                end else begin
                    I4a8abfa0896ce414d9b98093ef84455f  <= Ice174debd5dc911fdf5d5756cff8d731 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie3b00960f8af88a5aba7a2104dfca9a7 != Ibeb5edab51cd6aedad9c2ecedaded6f5[10] ) begin
                    Ic7147944f8835e26b9838fdbdc18ca41  <=  ~Ie369670edc5b602d305904f3a4a4381f + 1;
                end else begin
                    Ic7147944f8835e26b9838fdbdc18ca41  <= Ie369670edc5b602d305904f3a4a4381f ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie3b00960f8af88a5aba7a2104dfca9a7 != I2fbf89398a148c47810456812dbee5a6[4] ) begin
                    I7e393e6c1d1bc44daaab120d55f5dd59  <=  ~I41f66f79339962ef42fab3b88e571170 + 1;
                end else begin
                    I7e393e6c1d1bc44daaab120d55f5dd59  <= I41f66f79339962ef42fab3b88e571170 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie3b00960f8af88a5aba7a2104dfca9a7 != Iedd7d4ea8d082b40244c04946dfb14a0[4] ) begin
                    I356d747600182675699a2d2634d4c5ce  <=  ~I5cbd2fad4d90bd77ba3d2448a37ac60f + 1;
                end else begin
                    I356d747600182675699a2d2634d4c5ce  <= I5cbd2fad4d90bd77ba3d2448a37ac60f ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie3b00960f8af88a5aba7a2104dfca9a7 != Ia318eb500b8bd71048bde375c1db65a6[0] ) begin
                    I802c554d5b04af6b949677819a4966ed  <=  ~Id86a2869148e2885633d9e277f7041c3 + 1;
                end else begin
                    I802c554d5b04af6b949677819a4966ed  <= Id86a2869148e2885633d9e277f7041c3 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I7d1ef47f35b7a4c3ea2e4383732de398 != I5b7caaeb34c43e66e8d095a859e708fe[11] ) begin
                    I4f8792c18bd07b23e82bbc44b4ca947f  <=  ~Ifb7b585189db23efabfb522c9b45bede + 1;
                end else begin
                    I4f8792c18bd07b23e82bbc44b4ca947f  <= Ifb7b585189db23efabfb522c9b45bede ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I7d1ef47f35b7a4c3ea2e4383732de398 != I33a6ffad80ddf99a4d316a049078244d[4] ) begin
                    I3459d98131faef5a5040a03847890b55  <=  ~I7763f0d28d8065d8c94ef8df96b2ab06 + 1;
                end else begin
                    I3459d98131faef5a5040a03847890b55  <= I7763f0d28d8065d8c94ef8df96b2ab06 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I7d1ef47f35b7a4c3ea2e4383732de398 != I872f61d20baf011e867b44dc5539fc37[8] ) begin
                    I512cc8f6519aa08aee18225b56d47c9f  <=  ~I115ba88588187c7115977e95bd26ee5a + 1;
                end else begin
                    I512cc8f6519aa08aee18225b56d47c9f  <= I115ba88588187c7115977e95bd26ee5a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I7d1ef47f35b7a4c3ea2e4383732de398 != I4267622319ca65909a3b40484dc74d3a[5] ) begin
                    I4a41999cea9357a85c73a0af509eeac9  <=  ~I6e7f2bdd0c8231a3689893ef4877fdba + 1;
                end else begin
                    I4a41999cea9357a85c73a0af509eeac9  <= I6e7f2bdd0c8231a3689893ef4877fdba ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I7d1ef47f35b7a4c3ea2e4383732de398 != Ia2c4192b1e4f180402550aebcf1dcd1f[0] ) begin
                    Iceefb06cb3715e1b41e6f7d89420e5ba  <=  ~I546c513d5357ac1a6fe669888dfaf717 + 1;
                end else begin
                    Iceefb06cb3715e1b41e6f7d89420e5ba  <= I546c513d5357ac1a6fe669888dfaf717 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ibb013f036fc42687a04bdcbe2d0bbd8a != I61f0c04673dfb262ef6912eb2df39120[11] ) begin
                    Iaa5b2807e5cc2403c5787eeb3d10ca6b  <=  ~Ib3e12c614471912d0b276cb9f0382b1b + 1;
                end else begin
                    Iaa5b2807e5cc2403c5787eeb3d10ca6b  <= Ib3e12c614471912d0b276cb9f0382b1b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ibb013f036fc42687a04bdcbe2d0bbd8a != I980165c1147ac5ff86619c841c6031dc[4] ) begin
                    Iace01234164c8a9f7c98eeb83268745b  <=  ~I7187a2499e3319da90b6d6fc64411b46 + 1;
                end else begin
                    Iace01234164c8a9f7c98eeb83268745b  <= I7187a2499e3319da90b6d6fc64411b46 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ibb013f036fc42687a04bdcbe2d0bbd8a != I6f5c991e5fdcf56d582c6f80eb6731df[8] ) begin
                    I22c8ccd4a9018ad1c129aa058bf579d8  <=  ~I9b46582473bb4dd5541a35ac708486f4 + 1;
                end else begin
                    I22c8ccd4a9018ad1c129aa058bf579d8  <= I9b46582473bb4dd5541a35ac708486f4 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ibb013f036fc42687a04bdcbe2d0bbd8a != Iedd7d4ea8d082b40244c04946dfb14a0[5] ) begin
                    I87d6a5d30c3e4202cf51f33c7a770c51  <=  ~I929796fe327ee9c8a05e6bb683ae5d7c + 1;
                end else begin
                    I87d6a5d30c3e4202cf51f33c7a770c51  <= I929796fe327ee9c8a05e6bb683ae5d7c ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ibb013f036fc42687a04bdcbe2d0bbd8a != I1686a95674ecad0c4e234b8aa6e22dd9[0] ) begin
                    I56948bc48c0220893d68004615a6ebaa  <=  ~Ib6638da8b69373c2026d3f5305825cde + 1;
                end else begin
                    I56948bc48c0220893d68004615a6ebaa  <= Ib6638da8b69373c2026d3f5305825cde ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I77eae49d321f1d1e39dd7c75829aaedc != Ibeb5edab51cd6aedad9c2ecedaded6f5[11] ) begin
                    I698b1dbc9d8664d1c86c7a763d97b3b7  <=  ~I28c26bf4cf9693d1807818b2ca7883ac + 1;
                end else begin
                    I698b1dbc9d8664d1c86c7a763d97b3b7  <= I28c26bf4cf9693d1807818b2ca7883ac ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I77eae49d321f1d1e39dd7c75829aaedc != I19df055705f322292a3601fa63f0e5f9[4] ) begin
                    I68b575fcbc5321d4d26a22bcdbb506f6  <=  ~I291fc4eef4b80d1020c96488b869727e + 1;
                end else begin
                    I68b575fcbc5321d4d26a22bcdbb506f6  <= I291fc4eef4b80d1020c96488b869727e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I77eae49d321f1d1e39dd7c75829aaedc != Ia5cc3055ba3365e64cf59c4d4fd3f093[8] ) begin
                    Ib6aded6c73a8cc3cb964b0ae895b859e  <=  ~I53006ed50f6211439681aa7659647e35 + 1;
                end else begin
                    Ib6aded6c73a8cc3cb964b0ae895b859e  <= I53006ed50f6211439681aa7659647e35 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I77eae49d321f1d1e39dd7c75829aaedc != I56e1fe0c7a62589c123876f2b4e57a26[5] ) begin
                    I6ca8a1fa2c72b1c61d11dc7d1ba5f37b  <=  ~I47fe32973727237ae0cd4c306c7efbfb + 1;
                end else begin
                    I6ca8a1fa2c72b1c61d11dc7d1ba5f37b  <= I47fe32973727237ae0cd4c306c7efbfb ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I77eae49d321f1d1e39dd7c75829aaedc != I5ee21680396395f8338477fa2bb314ec[0] ) begin
                    Iec1368f034655d61354ab5b5e94d7d89  <=  ~Ic3e0c7d71f13a56a9a63e158c7f2cfa8 + 1;
                end else begin
                    Iec1368f034655d61354ab5b5e94d7d89  <= Ic3e0c7d71f13a56a9a63e158c7f2cfa8 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I420a4d69a077dc1996ddb4b715d63e15 != Iceb64ab2ff8a2e0dfdb74803811d4cfe[11] ) begin
                    I08ece7cd684e593e02321612b7a88cee  <=  ~If383f241447cbea4e18f4f79fcdbf144 + 1;
                end else begin
                    I08ece7cd684e593e02321612b7a88cee  <= If383f241447cbea4e18f4f79fcdbf144 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I420a4d69a077dc1996ddb4b715d63e15 != I3d50cfeaa4b69c09bb648b8873a6bc24[4] ) begin
                    Icdcd83341f6b5c404f91ec7e97d0550c  <=  ~Ia05354d3b4f61299d5897832639df2c2 + 1;
                end else begin
                    Icdcd83341f6b5c404f91ec7e97d0550c  <= Ia05354d3b4f61299d5897832639df2c2 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I420a4d69a077dc1996ddb4b715d63e15 != Iea7da1f43ba202d753b0edb0be8b3fcf[8] ) begin
                    I82f266e5792cdb6e7ebd264e246161f5  <=  ~I9faec40665477e8b3237773d606af2f0 + 1;
                end else begin
                    I82f266e5792cdb6e7ebd264e246161f5  <= I9faec40665477e8b3237773d606af2f0 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I420a4d69a077dc1996ddb4b715d63e15 != Ia8a468877c9f96713c8141df9205f92a[5] ) begin
                    Ie1b7257c99831ec5864f65958ecf14fb  <=  ~Id231ab3133d4bed02aad7e5f560ee5f0 + 1;
                end else begin
                    Ie1b7257c99831ec5864f65958ecf14fb  <= Id231ab3133d4bed02aad7e5f560ee5f0 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I420a4d69a077dc1996ddb4b715d63e15 != I005e89f0a9a9a52aec92752813a70f81[0] ) begin
                    I1e43c0aeeb8a2461d208eba24967af30  <=  ~I13616c8c7be221cf4d2c13ae87c38bed + 1;
                end else begin
                    I1e43c0aeeb8a2461d208eba24967af30  <= I13616c8c7be221cf4d2c13ae87c38bed ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I652202a4dc8f102d29334b4811f5628d != Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[10] ) begin
                    I11c1fc94a3bd6dffa17e1571cc6ae97c  <=  ~I8793bc728a4d423fb96a88c83bb9746f + 1;
                end else begin
                    I11c1fc94a3bd6dffa17e1571cc6ae97c  <= I8793bc728a4d423fb96a88c83bb9746f ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I652202a4dc8f102d29334b4811f5628d != I651d700a00d7004d8728bc7356f30926[4] ) begin
                    Ica6707efd6d44ba6bbb87c0593a3d828  <=  ~I2fb6af0f152232550a3cadd55656df20 + 1;
                end else begin
                    Ica6707efd6d44ba6bbb87c0593a3d828  <= I2fb6af0f152232550a3cadd55656df20 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I652202a4dc8f102d29334b4811f5628d != Ia5cc3055ba3365e64cf59c4d4fd3f093[9] ) begin
                    I939368b76d98b43826c68c7f468a5632  <=  ~I5144918fcd4ce1a061644240730fc52a + 1;
                end else begin
                    I939368b76d98b43826c68c7f468a5632  <= I5144918fcd4ce1a061644240730fc52a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I652202a4dc8f102d29334b4811f5628d != I0daca3ad02a67285295cd9fc330d8027[0] ) begin
                    Ia6eb85b127cf9c1a437611556296b967  <=  ~I1821eb21cdf8208ff6c2f28d963f7bd6 + 1;
                end else begin
                    Ia6eb85b127cf9c1a437611556296b967  <= I1821eb21cdf8208ff6c2f28d963f7bd6 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I0e33e0cdf39fc4cc99f6696e9f2784de != Ib58043c04b5c4c86c1c67e57cc66dcf7[10] ) begin
                    I93bb43c1b89d4c70a57bdc019d64fd22  <=  ~I80471575b1d4b69ef073056f798394ea + 1;
                end else begin
                    I93bb43c1b89d4c70a57bdc019d64fd22  <= I80471575b1d4b69ef073056f798394ea ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I0e33e0cdf39fc4cc99f6696e9f2784de != Ic2580cbeec8c11a19bd1e2ebc29d255e[4] ) begin
                    Iae449b74e50e0907feae9e60f2329426  <=  ~I890bf9b72cc3c71351547178d72796e5 + 1;
                end else begin
                    Iae449b74e50e0907feae9e60f2329426  <= I890bf9b72cc3c71351547178d72796e5 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I0e33e0cdf39fc4cc99f6696e9f2784de != Iea7da1f43ba202d753b0edb0be8b3fcf[9] ) begin
                    Ibfacfe5b83819afe7fbd4bffa2d6d4e2  <=  ~Icc9d28b84fa91028ae96cc9b8bae7555 + 1;
                end else begin
                    Ibfacfe5b83819afe7fbd4bffa2d6d4e2  <= Icc9d28b84fa91028ae96cc9b8bae7555 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I0e33e0cdf39fc4cc99f6696e9f2784de != I0d2ddde9edfef483482e6c177a084f6e[0] ) begin
                    Ieba89aa901e61218074af53a2484a74b  <=  ~I0b0d167c415f8c14594bd61907d46d80 + 1;
                end else begin
                    Ieba89aa901e61218074af53a2484a74b  <= I0b0d167c415f8c14594bd61907d46d80 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib9479328689dec62f900946e56ba0eb4 != Ibc0871b3c992fd278815fdbefcd2bac0[10] ) begin
                    Ie0ee5445c56a5f9b41640b57422206de  <=  ~I9577d49a74520355e53a1818f479db0e + 1;
                end else begin
                    Ie0ee5445c56a5f9b41640b57422206de  <= I9577d49a74520355e53a1818f479db0e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib9479328689dec62f900946e56ba0eb4 != If79ed5ee2b8710da0608c1e245d07d55[4] ) begin
                    Iacbb4daf5ce5c7eb1a2afe30d0cb5382  <=  ~Ie6e888d582ba9e600e91b119e2804642 + 1;
                end else begin
                    Iacbb4daf5ce5c7eb1a2afe30d0cb5382  <= Ie6e888d582ba9e600e91b119e2804642 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib9479328689dec62f900946e56ba0eb4 != I872f61d20baf011e867b44dc5539fc37[9] ) begin
                    If08370fd0e8af818c6db20f43e74034d  <=  ~Iccfac3d489b4b110d6b6e005a5ba45d8 + 1;
                end else begin
                    If08370fd0e8af818c6db20f43e74034d  <= Iccfac3d489b4b110d6b6e005a5ba45d8 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib9479328689dec62f900946e56ba0eb4 != I932ad562b582e2c9795f241c82901188[0] ) begin
                    I8b3b875c6c07bd97ba598a5139156fa4  <=  ~I69a67481ca8fd01dc5400dbe887b4f83 + 1;
                end else begin
                    I8b3b875c6c07bd97ba598a5139156fa4  <= I69a67481ca8fd01dc5400dbe887b4f83 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I2728682c0f749d1a9e8afeacdf44bfb7 != I8695e1e94cbfcbe4b9eae315b042529e[10] ) begin
                    I680be647bf2a62e0ee9b5d379dc87b4f  <=  ~I1f36f045becec7f0528f4a935d3da2ff + 1;
                end else begin
                    I680be647bf2a62e0ee9b5d379dc87b4f  <= I1f36f045becec7f0528f4a935d3da2ff ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I2728682c0f749d1a9e8afeacdf44bfb7 != I9497bbb4f746969a95cff948a3ee9ade[4] ) begin
                    Icbfbb37bad6344005dd233b3605a784f  <=  ~I530fe7720e3bcda35e940aa4973a7da4 + 1;
                end else begin
                    Icbfbb37bad6344005dd233b3605a784f  <= I530fe7720e3bcda35e940aa4973a7da4 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I2728682c0f749d1a9e8afeacdf44bfb7 != I6f5c991e5fdcf56d582c6f80eb6731df[9] ) begin
                    I83330fef69470d2f5def8e6d7d9c50d2  <=  ~I03069dda9fa863172d8747408800eeba + 1;
                end else begin
                    I83330fef69470d2f5def8e6d7d9c50d2  <= I03069dda9fa863172d8747408800eeba ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I2728682c0f749d1a9e8afeacdf44bfb7 != Ifee4aa12e36833c935c54ef27b1917da[0] ) begin
                    I7b33ddad346077928620344542b9481e  <=  ~Ie7f36ee89f2b092555fbf8031d2347d9 + 1;
                end else begin
                    I7b33ddad346077928620344542b9481e  <= Ie7f36ee89f2b092555fbf8031d2347d9 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I07da3bb5f943db6271fe1867a358df35 != I5b7caaeb34c43e66e8d095a859e708fe[12] ) begin
                    I8d0a1ae4c47edf1f2b99d1175aaa7197  <=  ~I18af7980562b28c537be3bea8dc5252b + 1;
                end else begin
                    I8d0a1ae4c47edf1f2b99d1175aaa7197  <= I18af7980562b28c537be3bea8dc5252b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I07da3bb5f943db6271fe1867a358df35 != I8b8b9c4777e6df3eb2b9313e69ef2c8c[5] ) begin
                    Ie5757e7b1647ab7d43cdbcf98cbb77fc  <=  ~I22ec20f9396d28ed39c5fc4bf060c44a + 1;
                end else begin
                    Ie5757e7b1647ab7d43cdbcf98cbb77fc  <= I22ec20f9396d28ed39c5fc4bf060c44a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I07da3bb5f943db6271fe1867a358df35 != I6f5c991e5fdcf56d582c6f80eb6731df[10] ) begin
                    I0539d598bbe3d50940329a282c801328  <=  ~I105eac4e38f4661c7c7ca32161e42baa + 1;
                end else begin
                    I0539d598bbe3d50940329a282c801328  <= I105eac4e38f4661c7c7ca32161e42baa ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I07da3bb5f943db6271fe1867a358df35 != Id6f07dee3e47f39e3b43329c26f690f7[3] ) begin
                    I8acc93b34974c1e708b0e1591f7b2d3d  <=  ~I5030734bfa54065cbef20c1350cd647d + 1;
                end else begin
                    I8acc93b34974c1e708b0e1591f7b2d3d  <= I5030734bfa54065cbef20c1350cd647d ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I07da3bb5f943db6271fe1867a358df35 != I51e5b79f738795719ac21c6a88711a01[0] ) begin
                    I11d967a5c5d14c88b5587d4cfed1d05f  <=  ~Ieccf25e3abd6bae7dcf08baf815f3439 + 1;
                end else begin
                    I11d967a5c5d14c88b5587d4cfed1d05f  <= Ieccf25e3abd6bae7dcf08baf815f3439 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I61fc44808c85a75909b9d9fd4035f147 != I61f0c04673dfb262ef6912eb2df39120[12] ) begin
                    I6da2b3a481ee71b85f3087b36b399288  <=  ~I600c21fca7901299f8e95e8fa0ea0eb0 + 1;
                end else begin
                    I6da2b3a481ee71b85f3087b36b399288  <= I600c21fca7901299f8e95e8fa0ea0eb0 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I61fc44808c85a75909b9d9fd4035f147 != I4a16e8e7946d9a8220304fc1be3fb362[5] ) begin
                    I280e20c20c0b4f26278b3de9b2ff84e4  <=  ~Ic4363dfd133124dd45ec2211499d0788 + 1;
                end else begin
                    I280e20c20c0b4f26278b3de9b2ff84e4  <= Ic4363dfd133124dd45ec2211499d0788 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I61fc44808c85a75909b9d9fd4035f147 != Ia5cc3055ba3365e64cf59c4d4fd3f093[10] ) begin
                    I544f6263f16cd5e0b7cf28c511a8f6e3  <=  ~I7c0bc779c09847e3beb0a139e8826511 + 1;
                end else begin
                    I544f6263f16cd5e0b7cf28c511a8f6e3  <= I7c0bc779c09847e3beb0a139e8826511 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I61fc44808c85a75909b9d9fd4035f147 != Ic7f04c065f8ff82c2288f1de77d37189[3] ) begin
                    Ie11da10808c4ca84f399535df6261307  <=  ~If64db4386bf8f7d07292f14e3b313520 + 1;
                end else begin
                    Ie11da10808c4ca84f399535df6261307  <= If64db4386bf8f7d07292f14e3b313520 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I61fc44808c85a75909b9d9fd4035f147 != I4e41e628a8af629421544cb4c6f45265[0] ) begin
                    I27458d76b3ac6520fb379405c6b2956f  <=  ~Ibf51e537b992c4b4c0539dda9948f45c + 1;
                end else begin
                    I27458d76b3ac6520fb379405c6b2956f  <= Ibf51e537b992c4b4c0539dda9948f45c ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ic5075ee0ad355c20dd45ed594f2a8c3f != Ibeb5edab51cd6aedad9c2ecedaded6f5[12] ) begin
                    I508bbade361787127e1a2e8687ec884c  <=  ~I9f83063bdc3c352024f702cb9dc71ce8 + 1;
                end else begin
                    I508bbade361787127e1a2e8687ec884c  <= I9f83063bdc3c352024f702cb9dc71ce8 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ic5075ee0ad355c20dd45ed594f2a8c3f != I07930a807994815de45864af579902c4[5] ) begin
                    Ic19486b6ab0373b9c0ad8f7597782d8f  <=  ~I72127f6d422ec68dcd47126b87b3d3b1 + 1;
                end else begin
                    Ic19486b6ab0373b9c0ad8f7597782d8f  <= I72127f6d422ec68dcd47126b87b3d3b1 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ic5075ee0ad355c20dd45ed594f2a8c3f != Iea7da1f43ba202d753b0edb0be8b3fcf[10] ) begin
                    Ib8e68a77ad8b9e7cf415bee17645c3f9  <=  ~I0b4a1b48d110b820d8d87f6e94d32988 + 1;
                end else begin
                    Ib8e68a77ad8b9e7cf415bee17645c3f9  <= I0b4a1b48d110b820d8d87f6e94d32988 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ic5075ee0ad355c20dd45ed594f2a8c3f != Ieb244944e7ee8236a207924f56fbc689[3] ) begin
                    Ie84be0ae8311d906eff08f7f5b214943  <=  ~I2e3aeede695007fabe0d6247a93ed403 + 1;
                end else begin
                    Ie84be0ae8311d906eff08f7f5b214943  <= I2e3aeede695007fabe0d6247a93ed403 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ic5075ee0ad355c20dd45ed594f2a8c3f != I9b2ec7db66661f7c9d85cfb1bc41893b[0] ) begin
                    I2525111a2fb5f10d64bbd16e148653b8  <=  ~I8c5ea3dc59fdcdea1c5f503dde1e815f + 1;
                end else begin
                    I2525111a2fb5f10d64bbd16e148653b8  <= I8c5ea3dc59fdcdea1c5f503dde1e815f ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ic0a651f45a502ead495cf14f97d65bfc != Iceb64ab2ff8a2e0dfdb74803811d4cfe[12] ) begin
                    I691c84d81c60a462e28e2b2bae3ea845  <=  ~I873c4dbe95220e40d7388870520261bd + 1;
                end else begin
                    I691c84d81c60a462e28e2b2bae3ea845  <= I873c4dbe95220e40d7388870520261bd ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ic0a651f45a502ead495cf14f97d65bfc != I72a2f42b727a0503d43332c0f22d5ae3[5] ) begin
                    I4904ab14b19fa1b6befc218bc7be3842  <=  ~I561fa67a9bfbedffcb04e7a4d6b76a64 + 1;
                end else begin
                    I4904ab14b19fa1b6befc218bc7be3842  <= I561fa67a9bfbedffcb04e7a4d6b76a64 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ic0a651f45a502ead495cf14f97d65bfc != I872f61d20baf011e867b44dc5539fc37[10] ) begin
                    I0ff382edfc8051459657ffa3899f5f73  <=  ~Ia55752d6c4f20378ff570a661ab31d9a + 1;
                end else begin
                    I0ff382edfc8051459657ffa3899f5f73  <= Ia55752d6c4f20378ff570a661ab31d9a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ic0a651f45a502ead495cf14f97d65bfc != Ie9b2be4c32334220e134e041ca8dfc06[3] ) begin
                    I8f94dbafaac589ac9f14b56d4556ff96  <=  ~Ia13307be43e9155ed0333df62ccc8bf2 + 1;
                end else begin
                    I8f94dbafaac589ac9f14b56d4556ff96  <= Ia13307be43e9155ed0333df62ccc8bf2 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ic0a651f45a502ead495cf14f97d65bfc != I0a594a36728c7ac6244c504b8ea9c9af[0] ) begin
                    I7b7cbcd1c6d2a2eeaaff474536a69eed  <=  ~I07b3d1451487a55fbbedda48b0cb6c73 + 1;
                end else begin
                    I7b7cbcd1c6d2a2eeaaff474536a69eed  <= I07b3d1451487a55fbbedda48b0cb6c73 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ic1c05ea22f708f620f626cc8c5ca309c != Iceb64ab2ff8a2e0dfdb74803811d4cfe[13] ) begin
                    I58dc9cce6384160c0a85c6efb3319cdb  <=  ~I9f8cf1a6cd0182fba35a49bd232f062a + 1;
                end else begin
                    I58dc9cce6384160c0a85c6efb3319cdb  <= I9f8cf1a6cd0182fba35a49bd232f062a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ic1c05ea22f708f620f626cc8c5ca309c != I04302edb2671c5bc0ca2673cd53935e1[5] ) begin
                    Icde3e6dbcf985682041f30903ad95572  <=  ~Ie2e488a8589559deeec8598cf6726f1f + 1;
                end else begin
                    Icde3e6dbcf985682041f30903ad95572  <= Ie2e488a8589559deeec8598cf6726f1f ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ic1c05ea22f708f620f626cc8c5ca309c != Iea7da1f43ba202d753b0edb0be8b3fcf[11] ) begin
                    I644ee0055a55f54ab3544bb532e39c61  <=  ~I9118ee5ff8c9ba9b125e5baa07bf52e0 + 1;
                end else begin
                    I644ee0055a55f54ab3544bb532e39c61  <= I9118ee5ff8c9ba9b125e5baa07bf52e0 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ic1c05ea22f708f620f626cc8c5ca309c != Ieb244944e7ee8236a207924f56fbc689[4] ) begin
                    Ic90b98708faa8c8b75d4bd9a52c292f7  <=  ~I13b894057e2deae2c00787385de252a8 + 1;
                end else begin
                    Ic90b98708faa8c8b75d4bd9a52c292f7  <= I13b894057e2deae2c00787385de252a8 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ic1c05ea22f708f620f626cc8c5ca309c != Ibd943ebf64fe56a1818d2bb8b9f9f8bd[0] ) begin
                    Id2a7f0781d18dccc7c4e0b383b7cddfa  <=  ~I7797a3ea5b97b514a797243cf9fe890a + 1;
                end else begin
                    Id2a7f0781d18dccc7c4e0b383b7cddfa  <= I7797a3ea5b97b514a797243cf9fe890a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I61a18378aadae4556da501ce997321b4 != I5b7caaeb34c43e66e8d095a859e708fe[13] ) begin
                    I734e601f5f9d568a44a48834559e04db  <=  ~I3af78697aacc410108d0be7fd13c686b + 1;
                end else begin
                    I734e601f5f9d568a44a48834559e04db  <= I3af78697aacc410108d0be7fd13c686b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I61a18378aadae4556da501ce997321b4 != I480a0f6d6c3eb936de10a72749f6cd3f[5] ) begin
                    I749e987266a20840bb8a4b1a2a2fc5b0  <=  ~I871cb63247618a543b444aa3f888fffe + 1;
                end else begin
                    I749e987266a20840bb8a4b1a2a2fc5b0  <= I871cb63247618a543b444aa3f888fffe ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I61a18378aadae4556da501ce997321b4 != I872f61d20baf011e867b44dc5539fc37[11] ) begin
                    I9d2864024148337277523ef7fa2e1600  <=  ~I124404013f8fc6b302661900b9ad8ed8 + 1;
                end else begin
                    I9d2864024148337277523ef7fa2e1600  <= I124404013f8fc6b302661900b9ad8ed8 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I61a18378aadae4556da501ce997321b4 != Ie9b2be4c32334220e134e041ca8dfc06[4] ) begin
                    I754563caea429d3d0e22df5d193b84eb  <=  ~I8e413271c9d13748a1aa2d1a018ff28f + 1;
                end else begin
                    I754563caea429d3d0e22df5d193b84eb  <= I8e413271c9d13748a1aa2d1a018ff28f ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I61a18378aadae4556da501ce997321b4 != I8c3ba90c84f9375001e727b711dead8d[0] ) begin
                    If8bc141d98ebe1be7fa81cde5c65868e  <=  ~I4d799e93b4dfcabd69977ddb25634a69 + 1;
                end else begin
                    If8bc141d98ebe1be7fa81cde5c65868e  <= I4d799e93b4dfcabd69977ddb25634a69 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib1fc521709a1ce2198fd8df5b41d0177 != I61f0c04673dfb262ef6912eb2df39120[13] ) begin
                    I11094e852295755925c3c61f1df81643  <=  ~I1487f0027b7d16f4bc85bb00e537cbaf + 1;
                end else begin
                    I11094e852295755925c3c61f1df81643  <= I1487f0027b7d16f4bc85bb00e537cbaf ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib1fc521709a1ce2198fd8df5b41d0177 != I50976b0051e84b6a42fc1dbabd7d20ae[5] ) begin
                    Ic419255414995e7168afb97b051fa64f  <=  ~I1a5cdaa10022adf0ffbbc0f58b3e690a + 1;
                end else begin
                    Ic419255414995e7168afb97b051fa64f  <= I1a5cdaa10022adf0ffbbc0f58b3e690a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib1fc521709a1ce2198fd8df5b41d0177 != I6f5c991e5fdcf56d582c6f80eb6731df[11] ) begin
                    I202f88fdc946494d55fc8831c2e8a34c  <=  ~I98246759d003e9bc6676ceb2d093a06b + 1;
                end else begin
                    I202f88fdc946494d55fc8831c2e8a34c  <= I98246759d003e9bc6676ceb2d093a06b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib1fc521709a1ce2198fd8df5b41d0177 != Id6f07dee3e47f39e3b43329c26f690f7[4] ) begin
                    Ib60d4ac0fcadcdfce5a14fb92f58423f  <=  ~Ia3c2dfb3c4a45091be7cfecfad11f3ec + 1;
                end else begin
                    Ib60d4ac0fcadcdfce5a14fb92f58423f  <= Ia3c2dfb3c4a45091be7cfecfad11f3ec ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib1fc521709a1ce2198fd8df5b41d0177 != I387ca23d0e2183522ab041ec48bffef4[0] ) begin
                    I8645e1326c66f5efef4b9c923599d1a3  <=  ~I74cda651bcb24472a7697ba017f831a4 + 1;
                end else begin
                    I8645e1326c66f5efef4b9c923599d1a3  <= I74cda651bcb24472a7697ba017f831a4 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I1bb5511c9cda1a595c45ecde48e9ebc7 != Ibeb5edab51cd6aedad9c2ecedaded6f5[13] ) begin
                    I2afeb2a7b199c0c6738938f156ae4274  <=  ~Id7ba55b14ac0f471142011dc2d57cc4b + 1;
                end else begin
                    I2afeb2a7b199c0c6738938f156ae4274  <= Id7ba55b14ac0f471142011dc2d57cc4b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I1bb5511c9cda1a595c45ecde48e9ebc7 != I82e0e091fba6f79cef97eacac4b43ecb[5] ) begin
                    I7992ea31927b4f0e268462a3b0f18c5d  <=  ~I5890643c88c4255a0e5efd45f8af3ee2 + 1;
                end else begin
                    I7992ea31927b4f0e268462a3b0f18c5d  <= I5890643c88c4255a0e5efd45f8af3ee2 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I1bb5511c9cda1a595c45ecde48e9ebc7 != Ia5cc3055ba3365e64cf59c4d4fd3f093[11] ) begin
                    I484545c4d2c869d79eb17f51e11070a3  <=  ~I4f53e4955e9e506a7169ae810da5dde6 + 1;
                end else begin
                    I484545c4d2c869d79eb17f51e11070a3  <= I4f53e4955e9e506a7169ae810da5dde6 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I1bb5511c9cda1a595c45ecde48e9ebc7 != Ic7f04c065f8ff82c2288f1de77d37189[4] ) begin
                    I280fa9d114e227cd649bf0e55e845651  <=  ~Ifc7c1ea337b122fb720767f1890f1a6a + 1;
                end else begin
                    I280fa9d114e227cd649bf0e55e845651  <= Ifc7c1ea337b122fb720767f1890f1a6a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I1bb5511c9cda1a595c45ecde48e9ebc7 != Ib933575f5224d414f87bc71fa7498534[0] ) begin
                    I0426ef66185128dd1ef4dbb68dcda585  <=  ~Id40d6f3a8dd09678b25b3e579dd5fb68 + 1;
                end else begin
                    I0426ef66185128dd1ef4dbb68dcda585  <= Id40d6f3a8dd09678b25b3e579dd5fb68 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I4a29c37ed36b6e12f1f8e263c92bdbc1 != Ib58043c04b5c4c86c1c67e57cc66dcf7[11] ) begin
                    I7a2e554d07bbea291f2cfc18694fca3a  <=  ~I7002830b0a5f40ba2a2fe7a00c7b6d58 + 1;
                end else begin
                    I7a2e554d07bbea291f2cfc18694fca3a  <= I7002830b0a5f40ba2a2fe7a00c7b6d58 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I4a29c37ed36b6e12f1f8e263c92bdbc1 != I980165c1147ac5ff86619c841c6031dc[5] ) begin
                    Iace8b3b3a4c16763132b5aaa6b24212d  <=  ~I3f377e8994959ef8182a08538e393d9a + 1;
                end else begin
                    Iace8b3b3a4c16763132b5aaa6b24212d  <= I3f377e8994959ef8182a08538e393d9a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I4a29c37ed36b6e12f1f8e263c92bdbc1 != I8e591d83170c8ba46d31c61935311b22[7] ) begin
                    Ib2f5f5fc77ea8b529f2471c54388f2d1  <=  ~I71bf29f3519e3238cec112ef97ce0579 + 1;
                end else begin
                    Ib2f5f5fc77ea8b529f2471c54388f2d1  <= I71bf29f3519e3238cec112ef97ce0579 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I4a29c37ed36b6e12f1f8e263c92bdbc1 != Ibfe1bddf32fa63ea87c68de7a3af1815[0] ) begin
                    Iddd954df5bae9b4240e0512f746669a9  <=  ~Iaa4bc2f51984f383479b597e6cd4c873 + 1;
                end else begin
                    Iddd954df5bae9b4240e0512f746669a9  <= Iaa4bc2f51984f383479b597e6cd4c873 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I4bf02a07719402890405fb2e7b679ed9 != Ibc0871b3c992fd278815fdbefcd2bac0[11] ) begin
                    Ie5f8620371236cb11c9e88c16b509ee8  <=  ~I9066a5cf776f80ebf89bdac1f2edb4ac + 1;
                end else begin
                    Ie5f8620371236cb11c9e88c16b509ee8  <= I9066a5cf776f80ebf89bdac1f2edb4ac ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I4bf02a07719402890405fb2e7b679ed9 != I19df055705f322292a3601fa63f0e5f9[5] ) begin
                    Idf600b93ee1018ecf969ed7944b6bc7b  <=  ~I7319203d7231bebb6d6e52422cce5ed2 + 1;
                end else begin
                    Idf600b93ee1018ecf969ed7944b6bc7b  <= I7319203d7231bebb6d6e52422cce5ed2 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I4bf02a07719402890405fb2e7b679ed9 != I02b62fafd371de339f299f8aefec6c43[7] ) begin
                    I7f90f96c0260560ad5e6dc7448b2670a  <=  ~I4e8309976fd6011d78728cef935dc3c1 + 1;
                end else begin
                    I7f90f96c0260560ad5e6dc7448b2670a  <= I4e8309976fd6011d78728cef935dc3c1 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I4bf02a07719402890405fb2e7b679ed9 != I719c50f9bbc66decebe794fe6ea017dd[0] ) begin
                    I29e940970d87e8e09b26ab1b0b8f2286  <=  ~I5ed502118c175d5bdb4607973554a3a3 + 1;
                end else begin
                    I29e940970d87e8e09b26ab1b0b8f2286  <= I5ed502118c175d5bdb4607973554a3a3 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I75bd82990cb60b6d7ccd7aa2982da7aa != I8695e1e94cbfcbe4b9eae315b042529e[11] ) begin
                    If4d75f83299a21802b6fbe136913489f  <=  ~If457f80b3d29b60b840f886fa928297c + 1;
                end else begin
                    If4d75f83299a21802b6fbe136913489f  <= If457f80b3d29b60b840f886fa928297c ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I75bd82990cb60b6d7ccd7aa2982da7aa != I3d50cfeaa4b69c09bb648b8873a6bc24[5] ) begin
                    Ibba4e82d1510ddc16eb4ef64893cec02  <=  ~I7e0f785ec7554540c9a4a413a3afa75f + 1;
                end else begin
                    Ibba4e82d1510ddc16eb4ef64893cec02  <= I7e0f785ec7554540c9a4a413a3afa75f ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I75bd82990cb60b6d7ccd7aa2982da7aa != I0e0b15868b02ca52b260f17f150d237e[7] ) begin
                    I108c269ceec4adcff9afeda01101b838  <=  ~Id3662bbe1b5191995d1656045fe6b6a6 + 1;
                end else begin
                    I108c269ceec4adcff9afeda01101b838  <= Id3662bbe1b5191995d1656045fe6b6a6 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I75bd82990cb60b6d7ccd7aa2982da7aa != I833b0433a33dac70cb215bc8cc9f4863[0] ) begin
                    I488f6d9676aa85a55d030bf12e8997a7  <=  ~Idf922fab93bc2357ac1f66f73f3ead0b + 1;
                end else begin
                    I488f6d9676aa85a55d030bf12e8997a7  <= Idf922fab93bc2357ac1f66f73f3ead0b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ia6d3e38249f8a1208540b68f54c46769 != Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[11] ) begin
                    I5395ee57418c31e11cf847f0f514ec19  <=  ~I780371393ef898aa144c5bc36e74c654 + 1;
                end else begin
                    I5395ee57418c31e11cf847f0f514ec19  <= I780371393ef898aa144c5bc36e74c654 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ia6d3e38249f8a1208540b68f54c46769 != I33a6ffad80ddf99a4d316a049078244d[5] ) begin
                    Ie9b9221b2122087cd5f309570b6d31ca  <=  ~I79696cd10cffa4c0181a2089da6b3262 + 1;
                end else begin
                    Ie9b9221b2122087cd5f309570b6d31ca  <= I79696cd10cffa4c0181a2089da6b3262 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ia6d3e38249f8a1208540b68f54c46769 != I3c0b6f53f0a5cda5b6758b2ee2c83b92[7] ) begin
                    I4eadce87f47df6d8f0e4acd057de5a09  <=  ~I073155ab0359a13b77f730653dcfc08d + 1;
                end else begin
                    I4eadce87f47df6d8f0e4acd057de5a09  <= I073155ab0359a13b77f730653dcfc08d ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ia6d3e38249f8a1208540b68f54c46769 != I9769761eb863e3273f9253ace4c69585[0] ) begin
                    I99d761b75ade1fb2e8afbb1a77752609  <=  ~I1b44f781d81438654f69bb7fbdb94011 + 1;
                end else begin
                    I99d761b75ade1fb2e8afbb1a77752609  <= I1b44f781d81438654f69bb7fbdb94011 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Idf548b72357ab28fd956791e84e5d65c != Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[12] ) begin
                    Iff125392fa39afebae1637a19c4e23ec  <=  ~Id68f1a0ec8ff80da3190fe517bd935e3 + 1;
                end else begin
                    Iff125392fa39afebae1637a19c4e23ec  <= Id68f1a0ec8ff80da3190fe517bd935e3 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Idf548b72357ab28fd956791e84e5d65c != I61f0c04673dfb262ef6912eb2df39120[14] ) begin
                    I9c633aa620cca127b0ff8cf882178e76  <=  ~I3704464d41956032b779eebe27511815 + 1;
                end else begin
                    I9c633aa620cca127b0ff8cf882178e76  <= I3704464d41956032b779eebe27511815 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Idf548b72357ab28fd956791e84e5d65c != If79ed5ee2b8710da0608c1e245d07d55[5] ) begin
                    I4e08021c0235fafb60200aab97827a8f  <=  ~Ie6756ee9631791940ffc6fddb223b4d0 + 1;
                end else begin
                    I4e08021c0235fafb60200aab97827a8f  <= Ie6756ee9631791940ffc6fddb223b4d0 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Idf548b72357ab28fd956791e84e5d65c != I1fc63f388d047207a9375842c85e87f7[0] ) begin
                    Iac4e3d20178049f9c59abf374752dccc  <=  ~I085151dfc2e773a7a485f5ef1b7cd6bd + 1;
                end else begin
                    Iac4e3d20178049f9c59abf374752dccc  <= I085151dfc2e773a7a485f5ef1b7cd6bd ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I50b6f2e0ef2831535ac8c18cd7ca9379 != Ib58043c04b5c4c86c1c67e57cc66dcf7[12] ) begin
                    I3e59b2419c7dd1553b792d536208514e  <=  ~I2654e83fff153df7760c341f59a23396 + 1;
                end else begin
                    I3e59b2419c7dd1553b792d536208514e  <= I2654e83fff153df7760c341f59a23396 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I50b6f2e0ef2831535ac8c18cd7ca9379 != Ibeb5edab51cd6aedad9c2ecedaded6f5[14] ) begin
                    I86255756ddd1f88b74e070b19f8c3bfa  <=  ~Iee3eec7a9d7a3a5c22281545ec143e50 + 1;
                end else begin
                    I86255756ddd1f88b74e070b19f8c3bfa  <= Iee3eec7a9d7a3a5c22281545ec143e50 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I50b6f2e0ef2831535ac8c18cd7ca9379 != I9497bbb4f746969a95cff948a3ee9ade[5] ) begin
                    I91a6408a11fab36a8ba3dbd3f895a803  <=  ~Ied2b9ca07a6d498abada30fb0726df24 + 1;
                end else begin
                    I91a6408a11fab36a8ba3dbd3f895a803  <= Ied2b9ca07a6d498abada30fb0726df24 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I50b6f2e0ef2831535ac8c18cd7ca9379 != I414c4d389ecc00197f2138eff0b6454e[0] ) begin
                    I618d33f26badabfa578908903a613bce  <=  ~If95315702519e7a08386a870e599aab0 + 1;
                end else begin
                    I618d33f26badabfa578908903a613bce  <= If95315702519e7a08386a870e599aab0 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I4003a2515229ca8eb6fefa2bef289ca6 != Ibc0871b3c992fd278815fdbefcd2bac0[12] ) begin
                    I8d7c1fe2e33bbd45379b0325a3c5e989  <=  ~I1091064aef7d915ba8fb6cbded069102 + 1;
                end else begin
                    I8d7c1fe2e33bbd45379b0325a3c5e989  <= I1091064aef7d915ba8fb6cbded069102 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I4003a2515229ca8eb6fefa2bef289ca6 != Iceb64ab2ff8a2e0dfdb74803811d4cfe[14] ) begin
                    I56bf74b5890ec67090f499afdc0a9c88  <=  ~I40685c7d2c8be12698f734ec6213b5b4 + 1;
                end else begin
                    I56bf74b5890ec67090f499afdc0a9c88  <= I40685c7d2c8be12698f734ec6213b5b4 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I4003a2515229ca8eb6fefa2bef289ca6 != I651d700a00d7004d8728bc7356f30926[5] ) begin
                    I739267bcc50c54b8a685cb3c6afc5cc1  <=  ~Icc7775fe34c162006b93662530fd4944 + 1;
                end else begin
                    I739267bcc50c54b8a685cb3c6afc5cc1  <= Icc7775fe34c162006b93662530fd4944 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I4003a2515229ca8eb6fefa2bef289ca6 != Ibe387e8fe6f35588e028ba29cda5b912[0] ) begin
                    I822d7973afe090b2764335f1b72dfd0e  <=  ~I2e6f1a5695ad23b8ca282b344832ee8e + 1;
                end else begin
                    I822d7973afe090b2764335f1b72dfd0e  <= I2e6f1a5695ad23b8ca282b344832ee8e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I48672f8b83eef8c406694676746469e7 != I8695e1e94cbfcbe4b9eae315b042529e[12] ) begin
                    Ibddfda6413e3dd2f483c3174ea836b6a  <=  ~I016ce894bebdaa7e56af9deb1ccfb3f5 + 1;
                end else begin
                    Ibddfda6413e3dd2f483c3174ea836b6a  <= I016ce894bebdaa7e56af9deb1ccfb3f5 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I48672f8b83eef8c406694676746469e7 != I5b7caaeb34c43e66e8d095a859e708fe[14] ) begin
                    Ie421da1dc5aaea57c50d0c7d9c5a2717  <=  ~Iad2dd0815c1107160992e5070632f76c + 1;
                end else begin
                    Ie421da1dc5aaea57c50d0c7d9c5a2717  <= Iad2dd0815c1107160992e5070632f76c ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I48672f8b83eef8c406694676746469e7 != Ic2580cbeec8c11a19bd1e2ebc29d255e[5] ) begin
                    Iebf769a6bdaf214c1006c55c608d4eda  <=  ~Iefaba2acd282081b9a0a98ed057ca85e + 1;
                end else begin
                    Iebf769a6bdaf214c1006c55c608d4eda  <= Iefaba2acd282081b9a0a98ed057ca85e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I48672f8b83eef8c406694676746469e7 != I98191a7e6c56aae1b56e3d623004ed75[0] ) begin
                    I12c1035353e553b3b6a13bb174ce6020  <=  ~Id4ef94eb8d5db8810bca4c9d669f0b7f + 1;
                end else begin
                    I12c1035353e553b3b6a13bb174ce6020  <= Id4ef94eb8d5db8810bca4c9d669f0b7f ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ia14a60c9497c0faf3f1f448ff2abe553 != Iceb64ab2ff8a2e0dfdb74803811d4cfe[15] ) begin
                    Ibaf2f1f8bda2f6b932dc30f8369c0e1f  <=  ~I04e845e6a5ed71978b636593dd749b12 + 1;
                end else begin
                    Ibaf2f1f8bda2f6b932dc30f8369c0e1f  <= I04e845e6a5ed71978b636593dd749b12 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ia14a60c9497c0faf3f1f448ff2abe553 != Ic2941d16ae6a5cbce70e8546a18ca4ff[3] ) begin
                    I88a61cf72347d695489909d0819332ab  <=  ~I0b2760b437be2cb79382f8d6a7b8969e + 1;
                end else begin
                    I88a61cf72347d695489909d0819332ab  <= I0b2760b437be2cb79382f8d6a7b8969e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ia14a60c9497c0faf3f1f448ff2abe553 != Ia5cc3055ba3365e64cf59c4d4fd3f093[12] ) begin
                    I39289e6385a9bc378a9b8dd440249a7f  <=  ~I1b0fdaeebe5fee6fbb2e13aac5e233a1 + 1;
                end else begin
                    I39289e6385a9bc378a9b8dd440249a7f  <= I1b0fdaeebe5fee6fbb2e13aac5e233a1 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ia14a60c9497c0faf3f1f448ff2abe553 != Icd0f5c370462670cd18d30dfc0c81c02[0] ) begin
                    Ia6d61947d36fc128c689808c82db80f6  <=  ~Iee872d17e4a28075be0ad7086c3acc91 + 1;
                end else begin
                    Ia6d61947d36fc128c689808c82db80f6  <= Iee872d17e4a28075be0ad7086c3acc91 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I0ef3962dd323e8ec64c4a881bd4b3044 != I5b7caaeb34c43e66e8d095a859e708fe[15] ) begin
                    Ief5cbddfbfb98fce4812a676849b9a98  <=  ~I87656ddd4ef8f1ae36c7566d5e7892d8 + 1;
                end else begin
                    Ief5cbddfbfb98fce4812a676849b9a98  <= I87656ddd4ef8f1ae36c7566d5e7892d8 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I0ef3962dd323e8ec64c4a881bd4b3044 != I8e29ebe9ee25ea8ef3e52ff56fc29157[3] ) begin
                    I3ca2b9b77ed8d78a10aff42a07a53b07  <=  ~I865cd0535644db7f17db1180c85f1744 + 1;
                end else begin
                    I3ca2b9b77ed8d78a10aff42a07a53b07  <= I865cd0535644db7f17db1180c85f1744 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I0ef3962dd323e8ec64c4a881bd4b3044 != Iea7da1f43ba202d753b0edb0be8b3fcf[12] ) begin
                    Ic5467e42aa377c6ffd8f70673808774f  <=  ~I71d46741fa94df65e1bdf6abff53d2ba + 1;
                end else begin
                    Ic5467e42aa377c6ffd8f70673808774f  <= I71d46741fa94df65e1bdf6abff53d2ba ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I0ef3962dd323e8ec64c4a881bd4b3044 != I15c59dc8eba10ff8eadfa6078678773b[0] ) begin
                    Ie9b042f686381739b9ff219041f1e0ce  <=  ~Ic223d7941250d739ce9bb0ae5013646e + 1;
                end else begin
                    Ie9b042f686381739b9ff219041f1e0ce  <= Ic223d7941250d739ce9bb0ae5013646e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie9b64c34e31dab63c03b3de4528d53fe != I61f0c04673dfb262ef6912eb2df39120[15] ) begin
                    I694d471fd353eb54aae08a2afa7b645a  <=  ~I1ef9b548b943a1f2012b91c7e0b445f2 + 1;
                end else begin
                    I694d471fd353eb54aae08a2afa7b645a  <= I1ef9b548b943a1f2012b91c7e0b445f2 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie9b64c34e31dab63c03b3de4528d53fe != Ic3742290179b27b9865f9d1f88d66266[3] ) begin
                    I15fafe2baba4d2f28037023a81ce0a81  <=  ~I88b6d7894d82ff394e89c7471c80dd5b + 1;
                end else begin
                    I15fafe2baba4d2f28037023a81ce0a81  <= I88b6d7894d82ff394e89c7471c80dd5b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie9b64c34e31dab63c03b3de4528d53fe != I872f61d20baf011e867b44dc5539fc37[12] ) begin
                    I1c85a2d1df6749a194072eb731506bfe  <=  ~Ia5fc7e1f991f30042b848888a546534b + 1;
                end else begin
                    I1c85a2d1df6749a194072eb731506bfe  <= Ia5fc7e1f991f30042b848888a546534b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie9b64c34e31dab63c03b3de4528d53fe != I3870d672343c002ad9c83c816fd40567[0] ) begin
                    I0c4268c01aed70ce4fc71531bf4bb862  <=  ~If699df4c8261ebce5c5d1aebe062cd61 + 1;
                end else begin
                    I0c4268c01aed70ce4fc71531bf4bb862  <= If699df4c8261ebce5c5d1aebe062cd61 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I5941476ded9f6dc25d7394f5d133955b != Ibeb5edab51cd6aedad9c2ecedaded6f5[15] ) begin
                    I7d4924388dc5373ad7936dca76797473  <=  ~I19338369553e96bb2476d80fe84dec3e + 1;
                end else begin
                    I7d4924388dc5373ad7936dca76797473  <= I19338369553e96bb2476d80fe84dec3e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I5941476ded9f6dc25d7394f5d133955b != I9ef21ef20099af28d9a8c794f70d45a5[3] ) begin
                    Ifa43d74fa91b7b9884969f575ef9ca8e  <=  ~I9844ff02042cbc04dd5f4179908bbb2d + 1;
                end else begin
                    Ifa43d74fa91b7b9884969f575ef9ca8e  <= I9844ff02042cbc04dd5f4179908bbb2d ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I5941476ded9f6dc25d7394f5d133955b != I6f5c991e5fdcf56d582c6f80eb6731df[12] ) begin
                    I3ee10f6a7785a236db317515fdd23a2d  <=  ~I89cc6a060b714985b24f724adc782e7b + 1;
                end else begin
                    I3ee10f6a7785a236db317515fdd23a2d  <= I89cc6a060b714985b24f724adc782e7b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I5941476ded9f6dc25d7394f5d133955b != Ic341b9d947f2d3ac57aa41f408214434[0] ) begin
                    Ia34e42f8de91fa4861b0c6cac5dcfc29  <=  ~I39d94ce7fbe37a74404e0043060441ed + 1;
                end else begin
                    Ia34e42f8de91fa4861b0c6cac5dcfc29  <= I39d94ce7fbe37a74404e0043060441ed ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib46c78ff661ee6fb69c704d39235ffe1 != Ib58043c04b5c4c86c1c67e57cc66dcf7[13] ) begin
                    I46894c6526983bf1ce4b503159131b41  <=  ~I0a1c9a8d59dbcffd6847f3a65107c407 + 1;
                end else begin
                    I46894c6526983bf1ce4b503159131b41  <= I0a1c9a8d59dbcffd6847f3a65107c407 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib46c78ff661ee6fb69c704d39235ffe1 != Icac5a9001ee113e612e3457b4b49ee68[5] ) begin
                    Icb82c9ff4cb58159a1c3115c6fdd5f8c  <=  ~I2328556c467a9e639f2b6ba1d0cb99b7 + 1;
                end else begin
                    Icb82c9ff4cb58159a1c3115c6fdd5f8c  <= I2328556c467a9e639f2b6ba1d0cb99b7 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib46c78ff661ee6fb69c704d39235ffe1 != I56e1fe0c7a62589c123876f2b4e57a26[6] ) begin
                    I3ec5819176ad4b0895a9118d90ab22b5  <=  ~I5c9d75d6431d69db1abe412e591000a7 + 1;
                end else begin
                    I3ec5819176ad4b0895a9118d90ab22b5  <= I5c9d75d6431d69db1abe412e591000a7 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib46c78ff661ee6fb69c704d39235ffe1 != Ied40f6b7847158bd08cbd932254dd6ba[0] ) begin
                    Ib7c5850b4f7cc77be2048d114a2128d9  <=  ~I8dc3dcdefc85b6ff8ecfa09cfc7e69fa + 1;
                end else begin
                    Ib7c5850b4f7cc77be2048d114a2128d9  <= I8dc3dcdefc85b6ff8ecfa09cfc7e69fa ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iadabc5abc7dfbc1dd747179ad7e37850 != Ibc0871b3c992fd278815fdbefcd2bac0[13] ) begin
                    I4fbdc4ee57a3be42b62d9bd43078d6ef  <=  ~I69f6c909ea6b207c200b154e00e13a05 + 1;
                end else begin
                    I4fbdc4ee57a3be42b62d9bd43078d6ef  <= I69f6c909ea6b207c200b154e00e13a05 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iadabc5abc7dfbc1dd747179ad7e37850 != I9461e92a5880cb9e04fcece2ef4674f0[5] ) begin
                    Ib3367565e4456da15e7c2315dccdb5e4  <=  ~Id365c9f8f7f97c777bd5da0ce9490511 + 1;
                end else begin
                    Ib3367565e4456da15e7c2315dccdb5e4  <= Id365c9f8f7f97c777bd5da0ce9490511 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iadabc5abc7dfbc1dd747179ad7e37850 != Ia8a468877c9f96713c8141df9205f92a[6] ) begin
                    I4accbad1b451ed2b622e15ef9ae16d13  <=  ~Idf0206d2ad2bdef7db1d30a2d715cc6a + 1;
                end else begin
                    I4accbad1b451ed2b622e15ef9ae16d13  <= Idf0206d2ad2bdef7db1d30a2d715cc6a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iadabc5abc7dfbc1dd747179ad7e37850 != I6ab04d323306b7290cc89ed66dbd93bf[0] ) begin
                    I32bb50faa2b246b2d3b462a79be597c5  <=  ~I07d1c54431eed887554a136f15f86d22 + 1;
                end else begin
                    I32bb50faa2b246b2d3b462a79be597c5  <= I07d1c54431eed887554a136f15f86d22 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I97a6b5f0976feceee3a5b5890d4d76a0 != I8695e1e94cbfcbe4b9eae315b042529e[13] ) begin
                    I33bddb0adcc2af7b12a83bf843036385  <=  ~Ic16809a3c82787ed88819fc9e9613f85 + 1;
                end else begin
                    I33bddb0adcc2af7b12a83bf843036385  <= Ic16809a3c82787ed88819fc9e9613f85 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I97a6b5f0976feceee3a5b5890d4d76a0 != I6ebab438dc55ccf6c1600313891d9c38[5] ) begin
                    I2c926fd9d306e9ae13364e07c4b0395b  <=  ~I1613ae89442495e703a52e65b8a0bf9f + 1;
                end else begin
                    I2c926fd9d306e9ae13364e07c4b0395b  <= I1613ae89442495e703a52e65b8a0bf9f ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I97a6b5f0976feceee3a5b5890d4d76a0 != I4267622319ca65909a3b40484dc74d3a[6] ) begin
                    I8e517c401d62dbb10dcc96ab536f6afb  <=  ~I6089da825af433e847c0b1bb9ff7d373 + 1;
                end else begin
                    I8e517c401d62dbb10dcc96ab536f6afb  <= I6089da825af433e847c0b1bb9ff7d373 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I97a6b5f0976feceee3a5b5890d4d76a0 != Iac4a5fdede87b021e6a8150d3bf34b66[0] ) begin
                    Idc6d40a49f05c5422758cee50f787eb1  <=  ~I6aa7fccf4e225fa70063fd24dab74e6b + 1;
                end else begin
                    Idc6d40a49f05c5422758cee50f787eb1  <= I6aa7fccf4e225fa70063fd24dab74e6b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I7217d4790fec9797a1eb8cab1ebce71b != Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[13] ) begin
                    Ia6308e16fae5428f4ab6560f5b21479a  <=  ~Ibe2a5f680405f233256b6fd806b72ae5 + 1;
                end else begin
                    Ia6308e16fae5428f4ab6560f5b21479a  <= Ibe2a5f680405f233256b6fd806b72ae5 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I7217d4790fec9797a1eb8cab1ebce71b != I2fbf89398a148c47810456812dbee5a6[5] ) begin
                    I448f126fd3932d5065abbe7bb2d92c56  <=  ~I662d408ffd8fb9f249e531a167161429 + 1;
                end else begin
                    I448f126fd3932d5065abbe7bb2d92c56  <= I662d408ffd8fb9f249e531a167161429 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I7217d4790fec9797a1eb8cab1ebce71b != Iedd7d4ea8d082b40244c04946dfb14a0[6] ) begin
                    I960768a84aec9d5b8bc7c1c523024a25  <=  ~Ie95b8a5c2da6c0877d49c646c194f5b7 + 1;
                end else begin
                    I960768a84aec9d5b8bc7c1c523024a25  <= Ie95b8a5c2da6c0877d49c646c194f5b7 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I7217d4790fec9797a1eb8cab1ebce71b != Id92b1676e19c5818fa813d06dc9a01f3[0] ) begin
                    Ide1d7dc22a4b271ef764df14ac22366a  <=  ~If940f33461f5e297e158db54f6aad610 + 1;
                end else begin
                    Ide1d7dc22a4b271ef764df14ac22366a  <= If940f33461f5e297e158db54f6aad610 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I3dd024db4130c105a6817e8a4935de0d != Iceb64ab2ff8a2e0dfdb74803811d4cfe[16] ) begin
                    Id9364a29fd79b52d0442e18dc0227854  <=  ~I54aa9d4c6333d94970eae97aeb3603fa + 1;
                end else begin
                    Id9364a29fd79b52d0442e18dc0227854  <= I54aa9d4c6333d94970eae97aeb3603fa ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I3dd024db4130c105a6817e8a4935de0d != If511a6ea6aa5cda5353658d8e192791f[2] ) begin
                    I2b2bd845428c49346ef8e94e95b618f8  <=  ~Ib82fc62720e6346e1c05cc33d596447e + 1;
                end else begin
                    I2b2bd845428c49346ef8e94e95b618f8  <= Ib82fc62720e6346e1c05cc33d596447e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I3dd024db4130c105a6817e8a4935de0d != I93da1192f27c33e21e03b9a2748774ea[0] ) begin
                    I7ace6778ac86b3e05939a3fcc716136f  <=  ~I24873624848b61f313865e10e77e35c6 + 1;
                end else begin
                    I7ace6778ac86b3e05939a3fcc716136f  <= I24873624848b61f313865e10e77e35c6 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iae502e5a5ae518fb7b817afff28b7932 != I5b7caaeb34c43e66e8d095a859e708fe[16] ) begin
                    Id113cab2dd1949d32e3c1c15273185c8  <=  ~Icc3915d8325c22fc172f731553798fef + 1;
                end else begin
                    Id113cab2dd1949d32e3c1c15273185c8  <= Icc3915d8325c22fc172f731553798fef ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iae502e5a5ae518fb7b817afff28b7932 != Ib0bf69cc797f330fb2546eb46d2d6f76[2] ) begin
                    I103f1449c78c47396d6a54dc1c810934  <=  ~I93b9837e63103431a0fdaf319a465c90 + 1;
                end else begin
                    I103f1449c78c47396d6a54dc1c810934  <= I93b9837e63103431a0fdaf319a465c90 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iae502e5a5ae518fb7b817afff28b7932 != I69a0c79d41af6b6340430b8b337fb0ca[0] ) begin
                    I044e01e8d2df46e03f00a0af2beb0bf5  <=  ~I91237af3aa2af551dbbc626bb701215e + 1;
                end else begin
                    I044e01e8d2df46e03f00a0af2beb0bf5  <= I91237af3aa2af551dbbc626bb701215e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib8b2b1d90204af5b100379ecad20fc0f != I61f0c04673dfb262ef6912eb2df39120[16] ) begin
                    I816704585ad393f685731104ad3ec64f  <=  ~Ib254d9701567f642d3586641edf85128 + 1;
                end else begin
                    I816704585ad393f685731104ad3ec64f  <= Ib254d9701567f642d3586641edf85128 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib8b2b1d90204af5b100379ecad20fc0f != Iec7404bc79c58d4d2538fcdf659e9134[2] ) begin
                    I53121a39de0bcba91a4d0438be2ae958  <=  ~I25c50067a62d2b3599d15f12f89d384e + 1;
                end else begin
                    I53121a39de0bcba91a4d0438be2ae958  <= I25c50067a62d2b3599d15f12f89d384e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib8b2b1d90204af5b100379ecad20fc0f != Ibd47f48d306ec44d94865a0a81e4f9dc[0] ) begin
                    I45a7ddcda2662e36b7617dfe64514346  <=  ~I238be7f0e4a209a6b4201a024c8aed82 + 1;
                end else begin
                    I45a7ddcda2662e36b7617dfe64514346  <= I238be7f0e4a209a6b4201a024c8aed82 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Idf0e651d0b13e167df3c0cc40d149c29 != Ibeb5edab51cd6aedad9c2ecedaded6f5[16] ) begin
                    Ie317e5ea2ca4ba2060d0f491290af96f  <=  ~I233f5ddadd45c0df2108ea6c1d634f3c + 1;
                end else begin
                    Ie317e5ea2ca4ba2060d0f491290af96f  <= I233f5ddadd45c0df2108ea6c1d634f3c ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Idf0e651d0b13e167df3c0cc40d149c29 != Ie1cd04c7668d3f450c387a6c1ad778c7[2] ) begin
                    I58703e8b6d04f8c69ac38f5fcfdc4efc  <=  ~I87a320ddaa1478146ff6e519dc65c40a + 1;
                end else begin
                    I58703e8b6d04f8c69ac38f5fcfdc4efc  <= I87a320ddaa1478146ff6e519dc65c40a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Idf0e651d0b13e167df3c0cc40d149c29 != Ia5707d1275138a5145b2a42190d95183[0] ) begin
                    Idada779a1ac7b844867571d77054b657  <=  ~Ibf03d6940c0a38bef038a28b6a7b625d + 1;
                end else begin
                    Idada779a1ac7b844867571d77054b657  <= Ibf03d6940c0a38bef038a28b6a7b625d ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I89daaca029498d05ca62c095db439eb5 != Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[14] ) begin
                    I5ea02b5349cd4d99ccbcb6b26f0cfdd7  <=  ~I90942470e2057e50ce4f5745ed68b81c + 1;
                end else begin
                    I5ea02b5349cd4d99ccbcb6b26f0cfdd7  <= I90942470e2057e50ce4f5745ed68b81c ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I89daaca029498d05ca62c095db439eb5 != I9c0b88a0be66d62f8ab061aeaee7e60f[4] ) begin
                    I30b0b1d54912c1a41a02a25ab238bb54  <=  ~I77fbc3f3b65962b610e39f4b085ecb7e + 1;
                end else begin
                    I30b0b1d54912c1a41a02a25ab238bb54  <= I77fbc3f3b65962b610e39f4b085ecb7e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I89daaca029498d05ca62c095db439eb5 != I50976b0051e84b6a42fc1dbabd7d20ae[6] ) begin
                    Iee6da3120d73373627b25ab7c0dedd28  <=  ~I701845efaf1b02aefa381d4f6b45c401 + 1;
                end else begin
                    Iee6da3120d73373627b25ab7c0dedd28  <= I701845efaf1b02aefa381d4f6b45c401 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I89daaca029498d05ca62c095db439eb5 != I33bc2f42d997a2963b063326eb210d1c[0] ) begin
                    Ieeba01b18a244ab8c0ac263c138fabcc  <=  ~Id446ddfd713c6e1592c562cfb123ea8b + 1;
                end else begin
                    Ieeba01b18a244ab8c0ac263c138fabcc  <= Id446ddfd713c6e1592c562cfb123ea8b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I0fe5a34ceda936d0924efdd07fad11e5 != Ib58043c04b5c4c86c1c67e57cc66dcf7[14] ) begin
                    I6404d0df952b5bf8292c753e4c6f35d8  <=  ~If4f752779d27392e7536565d425bce25 + 1;
                end else begin
                    I6404d0df952b5bf8292c753e4c6f35d8  <= If4f752779d27392e7536565d425bce25 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I0fe5a34ceda936d0924efdd07fad11e5 != Id88b9265ff08e0730e6a41abe1f80a32[4] ) begin
                    I913d818403024510c55b65b56a38dd89  <=  ~If112169057d6293326a56443ac3cf517 + 1;
                end else begin
                    I913d818403024510c55b65b56a38dd89  <= If112169057d6293326a56443ac3cf517 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I0fe5a34ceda936d0924efdd07fad11e5 != I82e0e091fba6f79cef97eacac4b43ecb[6] ) begin
                    Iadf927d18644a232ad1f1eba7db82934  <=  ~I78f727f8d85b5d7f0ffa57f02538f939 + 1;
                end else begin
                    Iadf927d18644a232ad1f1eba7db82934  <= I78f727f8d85b5d7f0ffa57f02538f939 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I0fe5a34ceda936d0924efdd07fad11e5 != Ib22e39b701614cd9986061c32adfbc66[0] ) begin
                    Ie4c9797a955778694dd8615219cb51e7  <=  ~I01ec629f60c17c2251f977205234cd44 + 1;
                end else begin
                    Ie4c9797a955778694dd8615219cb51e7  <= I01ec629f60c17c2251f977205234cd44 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I7876cbb2b5d8aba3652ec8b218080dff != Ibc0871b3c992fd278815fdbefcd2bac0[14] ) begin
                    I5510b88bfd65811b3200adf4ef975b48  <=  ~I23f774adb64807c0edaa9941c75651b6 + 1;
                end else begin
                    I5510b88bfd65811b3200adf4ef975b48  <= I23f774adb64807c0edaa9941c75651b6 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I7876cbb2b5d8aba3652ec8b218080dff != I6330943c9295298c53e889d47c7904d9[4] ) begin
                    I7774313f1ae5a2de98855aad572b3676  <=  ~I2361ef4fd70e4c05b25289d0845564c4 + 1;
                end else begin
                    I7774313f1ae5a2de98855aad572b3676  <= I2361ef4fd70e4c05b25289d0845564c4 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I7876cbb2b5d8aba3652ec8b218080dff != I04302edb2671c5bc0ca2673cd53935e1[6] ) begin
                    I46ee30b46020d91707689f3468f00e26  <=  ~Ic3067b434ca17be7bad595e1f9b822c5 + 1;
                end else begin
                    I46ee30b46020d91707689f3468f00e26  <= Ic3067b434ca17be7bad595e1f9b822c5 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I7876cbb2b5d8aba3652ec8b218080dff != I9b08176fde1cd08c9d7686a659213580[0] ) begin
                    I28a5ed4c239e64c76bb6e566b50cfd23  <=  ~I3546ddbae9c9db4517802db56cee35f0 + 1;
                end else begin
                    I28a5ed4c239e64c76bb6e566b50cfd23  <= I3546ddbae9c9db4517802db56cee35f0 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (If692ff56ce90d22d7af881599c54df75 != I8695e1e94cbfcbe4b9eae315b042529e[14] ) begin
                    I529f92b82248efe2cf64f7da0ec8283c  <=  ~I35e91092ed503831ed818f36a1ce1537 + 1;
                end else begin
                    I529f92b82248efe2cf64f7da0ec8283c  <= I35e91092ed503831ed818f36a1ce1537 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (If692ff56ce90d22d7af881599c54df75 != I5686b595177e07dd5bf231a35ee41659[4] ) begin
                    I7846bc2cc11e08d05f7c853c4920d555  <=  ~I973f185cf29e13193abf0108d4faa9d1 + 1;
                end else begin
                    I7846bc2cc11e08d05f7c853c4920d555  <= I973f185cf29e13193abf0108d4faa9d1 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (If692ff56ce90d22d7af881599c54df75 != I480a0f6d6c3eb936de10a72749f6cd3f[6] ) begin
                    I7607af5d98e8070e3d15cee23cdf877e  <=  ~Iee58b0442a6cccf0990ebb551b47fa92 + 1;
                end else begin
                    I7607af5d98e8070e3d15cee23cdf877e  <= Iee58b0442a6cccf0990ebb551b47fa92 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (If692ff56ce90d22d7af881599c54df75 != I1b4e65357a818998d08b83d21584e18c[0] ) begin
                    I79a705ee1e414fe4a5fb14e9b3ce9597  <=  ~I2cb3207a5c1b25386ac7eb532955f260 + 1;
                end else begin
                    I79a705ee1e414fe4a5fb14e9b3ce9597  <= I2cb3207a5c1b25386ac7eb532955f260 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I18a7a4fe8931c79df3a69223af46c440 != Iceb64ab2ff8a2e0dfdb74803811d4cfe[17] ) begin
                    Ica3a41ace27f7d94377981079952f4f7  <=  ~Icd4f07bc30c66f7f5b431ed97e7ac7b6 + 1;
                end else begin
                    Ica3a41ace27f7d94377981079952f4f7  <= Icd4f07bc30c66f7f5b431ed97e7ac7b6 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I18a7a4fe8931c79df3a69223af46c440 != If511a6ea6aa5cda5353658d8e192791f[3] ) begin
                    Ib730fdb59198f23d1e590f6d6039e96a  <=  ~Ifec6f3a1e10144acb320d5d502ed1ea3 + 1;
                end else begin
                    Ib730fdb59198f23d1e590f6d6039e96a  <= Ifec6f3a1e10144acb320d5d502ed1ea3 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I18a7a4fe8931c79df3a69223af46c440 != I07930a807994815de45864af579902c4[6] ) begin
                    I31243de90dc2a1656ca9d5e03bdd78da  <=  ~Ic87bff64a597e6d02583041b552328ee + 1;
                end else begin
                    I31243de90dc2a1656ca9d5e03bdd78da  <= Ic87bff64a597e6d02583041b552328ee ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I18a7a4fe8931c79df3a69223af46c440 != Ibb865ea5891db706b7b54e5c6fa383d0[0] ) begin
                    I04f90a907f10a7fa1ae3591b48094d5c  <=  ~I489f21ef8243ef8caa1c29f034c3e2ac + 1;
                end else begin
                    I04f90a907f10a7fa1ae3591b48094d5c  <= I489f21ef8243ef8caa1c29f034c3e2ac ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I8eec3538b8cc9c046954b6804cc656b0 != I5b7caaeb34c43e66e8d095a859e708fe[17] ) begin
                    Icfe1a689e33b2b9aa9dba692d6d610b9  <=  ~I773901563077961acada85962209d68a + 1;
                end else begin
                    Icfe1a689e33b2b9aa9dba692d6d610b9  <= I773901563077961acada85962209d68a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I8eec3538b8cc9c046954b6804cc656b0 != Ib0bf69cc797f330fb2546eb46d2d6f76[3] ) begin
                    I56b3a97dc3037f0bb2eed93a9482c813  <=  ~Ifbd176fe3e78bc2dc2e0e77ba3ccd2d0 + 1;
                end else begin
                    I56b3a97dc3037f0bb2eed93a9482c813  <= Ifbd176fe3e78bc2dc2e0e77ba3ccd2d0 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I8eec3538b8cc9c046954b6804cc656b0 != I72a2f42b727a0503d43332c0f22d5ae3[6] ) begin
                    I282d2eb4e74e034694e33273b9cb19d5  <=  ~I53f68a4cb81c71ee7bd6f61171b7478d + 1;
                end else begin
                    I282d2eb4e74e034694e33273b9cb19d5  <= I53f68a4cb81c71ee7bd6f61171b7478d ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I8eec3538b8cc9c046954b6804cc656b0 != I32d42cfd2d516af2e68fc2db4d5dce03[0] ) begin
                    I31d25b1b49e65216e90b39aa27acd6be  <=  ~I7568ec59f1359bedce86dbc6af50df71 + 1;
                end else begin
                    I31d25b1b49e65216e90b39aa27acd6be  <= I7568ec59f1359bedce86dbc6af50df71 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I653767e659590c1676edf6c25fc0e253 != I61f0c04673dfb262ef6912eb2df39120[17] ) begin
                    I85d95015a9ce27a18ccbf73bbbcdbd70  <=  ~Id2bf82d6bf0a201f80a58357038a0992 + 1;
                end else begin
                    I85d95015a9ce27a18ccbf73bbbcdbd70  <= Id2bf82d6bf0a201f80a58357038a0992 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I653767e659590c1676edf6c25fc0e253 != Iec7404bc79c58d4d2538fcdf659e9134[3] ) begin
                    Iff7950f24f0a6b0073942c37fff49d37  <=  ~I22442354ca2b77306f25839ce6124699 + 1;
                end else begin
                    Iff7950f24f0a6b0073942c37fff49d37  <= I22442354ca2b77306f25839ce6124699 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I653767e659590c1676edf6c25fc0e253 != I8b8b9c4777e6df3eb2b9313e69ef2c8c[6] ) begin
                    I6072331f838d82329a07a4ffa340c7b6  <=  ~I71a5c2876a07d8edd001ef2d108e59c1 + 1;
                end else begin
                    I6072331f838d82329a07a4ffa340c7b6  <= I71a5c2876a07d8edd001ef2d108e59c1 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I653767e659590c1676edf6c25fc0e253 != I4d0e8d475a5d2a7da24daca60f23f3d6[0] ) begin
                    I1f6540c5f037d861dee2c0091cba01ec  <=  ~Iaf333aa6b135927cf1ad1f76298ccd63 + 1;
                end else begin
                    I1f6540c5f037d861dee2c0091cba01ec  <= Iaf333aa6b135927cf1ad1f76298ccd63 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I5ff863be142b92dff89f7916d0d088c1 != Ibeb5edab51cd6aedad9c2ecedaded6f5[17] ) begin
                    I56ea52c50a188ec47e48740839a031c9  <=  ~Ia71cfd8cf9bea4e600ea204e41271c7d + 1;
                end else begin
                    I56ea52c50a188ec47e48740839a031c9  <= Ia71cfd8cf9bea4e600ea204e41271c7d ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I5ff863be142b92dff89f7916d0d088c1 != Ie1cd04c7668d3f450c387a6c1ad778c7[3] ) begin
                    Ie1f41720e296ced1b74cb325b666d88f  <=  ~I164b032929ac2b8cf1a6672859639a30 + 1;
                end else begin
                    Ie1f41720e296ced1b74cb325b666d88f  <= I164b032929ac2b8cf1a6672859639a30 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I5ff863be142b92dff89f7916d0d088c1 != I4a16e8e7946d9a8220304fc1be3fb362[6] ) begin
                    Ib3a0307176d424a4733720416d71069d  <=  ~I2ef0447f5c64fd5c65e23c16069a62ef + 1;
                end else begin
                    Ib3a0307176d424a4733720416d71069d  <= I2ef0447f5c64fd5c65e23c16069a62ef ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I5ff863be142b92dff89f7916d0d088c1 != Ie3850345b207e59aaaa5c944dab40b90[0] ) begin
                    I9632bb500b7faaaaeb649d74c21cbe8c  <=  ~Ide7008ee7f1fba156dc6145b3505e553 + 1;
                end else begin
                    I9632bb500b7faaaaeb649d74c21cbe8c  <= Ide7008ee7f1fba156dc6145b3505e553 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I49f9fd0e0719be527f2a54814dab83ea != Ib58043c04b5c4c86c1c67e57cc66dcf7[15] ) begin
                    I8522c402e654d007abffcb0e904af5e6  <=  ~I129a7ced6bc6f48f20fa552e2519925c + 1;
                end else begin
                    I8522c402e654d007abffcb0e904af5e6  <= I129a7ced6bc6f48f20fa552e2519925c ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I49f9fd0e0719be527f2a54814dab83ea != I04302edb2671c5bc0ca2673cd53935e1[7] ) begin
                    I2605f078c1a9006c93855a9a2b0cf6b9  <=  ~I67123cf825352e52cf0158060ad69a13 + 1;
                end else begin
                    I2605f078c1a9006c93855a9a2b0cf6b9  <= I67123cf825352e52cf0158060ad69a13 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I49f9fd0e0719be527f2a54814dab83ea != I4a9a1c932db30dcf04cb105a8d7384f9[0] ) begin
                    Idd0217a35c3adc8abc7bb581a5df7a2d  <=  ~I09923d784a9f9625a37221f639537941 + 1;
                end else begin
                    Idd0217a35c3adc8abc7bb581a5df7a2d  <= I09923d784a9f9625a37221f639537941 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I945f2476eb599844cbee0cd89038e392 != Ibc0871b3c992fd278815fdbefcd2bac0[15] ) begin
                    Ib57ef2f577cca54713c16717cbbd1ce9  <=  ~I5947be93fdb18bf0ad341fb826c9e6d7 + 1;
                end else begin
                    Ib57ef2f577cca54713c16717cbbd1ce9  <= I5947be93fdb18bf0ad341fb826c9e6d7 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I945f2476eb599844cbee0cd89038e392 != I480a0f6d6c3eb936de10a72749f6cd3f[7] ) begin
                    I2e11a697d7f17ac30302eadb500de72d  <=  ~I08621ee033cd49702ad08af4d31eb999 + 1;
                end else begin
                    I2e11a697d7f17ac30302eadb500de72d  <= I08621ee033cd49702ad08af4d31eb999 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I945f2476eb599844cbee0cd89038e392 != I0ef689822226332f5feaf79fcf8f6674[0] ) begin
                    Ic05b46168884322644db4e331d37d759  <=  ~Id5eca60b22d3835119571fe4b1a03479 + 1;
                end else begin
                    Ic05b46168884322644db4e331d37d759  <= Id5eca60b22d3835119571fe4b1a03479 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ied0c5f8a9243cd9d93672ad6cc907d21 != I8695e1e94cbfcbe4b9eae315b042529e[15] ) begin
                    I2f34af0036985cd94ade9cc905bec065  <=  ~I7267ba2b9cb511a48a3a7044e854f7da + 1;
                end else begin
                    I2f34af0036985cd94ade9cc905bec065  <= I7267ba2b9cb511a48a3a7044e854f7da ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ied0c5f8a9243cd9d93672ad6cc907d21 != I50976b0051e84b6a42fc1dbabd7d20ae[7] ) begin
                    I56fc99a22960232b305d6e683c66fcc7  <=  ~I5893fa21ec8bbdcea9677cc12fc4057a + 1;
                end else begin
                    I56fc99a22960232b305d6e683c66fcc7  <= I5893fa21ec8bbdcea9677cc12fc4057a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ied0c5f8a9243cd9d93672ad6cc907d21 != Ib5744c2130bb5a9d0ccdd975fdf2ff9c[0] ) begin
                    I53c88dc237bb2cd02d50fd7f0a168a48  <=  ~I564896fe01ec799a0fbe790473753559 + 1;
                end else begin
                    I53c88dc237bb2cd02d50fd7f0a168a48  <= I564896fe01ec799a0fbe790473753559 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9134c7f579723c7615af60b4344efe76 != Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[15] ) begin
                    I21de4f6194dec9e3c401934db92c25e7  <=  ~If279ab7c515c4039c8272b913c2fa107 + 1;
                end else begin
                    I21de4f6194dec9e3c401934db92c25e7  <= If279ab7c515c4039c8272b913c2fa107 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9134c7f579723c7615af60b4344efe76 != I82e0e091fba6f79cef97eacac4b43ecb[7] ) begin
                    I2a9c673cdd7ded79e09ada38c0f47e6f  <=  ~Ib61705ff5820f531eb17c40ed05f6ec3 + 1;
                end else begin
                    I2a9c673cdd7ded79e09ada38c0f47e6f  <= Ib61705ff5820f531eb17c40ed05f6ec3 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9134c7f579723c7615af60b4344efe76 != I039a7ddcb25972501d80c45c938cf683[0] ) begin
                    I7450d4ab3ef0227e93a02bfd620d047b  <=  ~I50149e5de41ca2998c4e8cc4b19e166b + 1;
                end else begin
                    I7450d4ab3ef0227e93a02bfd620d047b  <= I50149e5de41ca2998c4e8cc4b19e166b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie92388a9d1e71d73c07ed86e9bf6c887 != Iec7404bc79c58d4d2538fcdf659e9134[4] ) begin
                    Ide86f019e9573706c25bd8b4552396a8  <=  ~Id40cac3272643f3f91b73c6aa1740f3b + 1;
                end else begin
                    Ide86f019e9573706c25bd8b4552396a8  <= Id40cac3272643f3f91b73c6aa1740f3b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie92388a9d1e71d73c07ed86e9bf6c887 != I02b62fafd371de339f299f8aefec6c43[8] ) begin
                    I07b417cdcc99eaea3413f563e26ddc73  <=  ~Ic63eee2d700493c41ee2d186ff7111b9 + 1;
                end else begin
                    I07b417cdcc99eaea3413f563e26ddc73  <= Ic63eee2d700493c41ee2d186ff7111b9 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie92388a9d1e71d73c07ed86e9bf6c887 != Ieb244944e7ee8236a207924f56fbc689[5] ) begin
                    I8eba6f14f42701d22859fbea94bd1871  <=  ~I51de42598e0df4a76cf7b02c61ae9550 + 1;
                end else begin
                    I8eba6f14f42701d22859fbea94bd1871  <= I51de42598e0df4a76cf7b02c61ae9550 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie92388a9d1e71d73c07ed86e9bf6c887 != I56e1fe0c7a62589c123876f2b4e57a26[7] ) begin
                    I49b64469d298012dbb131d879bff38d6  <=  ~Ia89a1a58f6327ee3c105cae860942171 + 1;
                end else begin
                    I49b64469d298012dbb131d879bff38d6  <= Ia89a1a58f6327ee3c105cae860942171 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie92388a9d1e71d73c07ed86e9bf6c887 != Ic5f36c15ebad061dfbd5301e02ce2ffe[0] ) begin
                    I2b16e5b4e279bb29c3c675b72083e5fe  <=  ~Ib149a5872e31cd5df77b66298b4aad12 + 1;
                end else begin
                    I2b16e5b4e279bb29c3c675b72083e5fe  <= Ib149a5872e31cd5df77b66298b4aad12 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I6804fecdf59233c6cf14409bf2f1e430 != Ie1cd04c7668d3f450c387a6c1ad778c7[4] ) begin
                    I5d5701435c96f1078e741921b56e3c65  <=  ~Iaa16c14572ad0442eb3c58a97bef5ada + 1;
                end else begin
                    I5d5701435c96f1078e741921b56e3c65  <= Iaa16c14572ad0442eb3c58a97bef5ada ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I6804fecdf59233c6cf14409bf2f1e430 != I0e0b15868b02ca52b260f17f150d237e[8] ) begin
                    I761983331fb6e3c6c437b3f1660f0b6b  <=  ~I88d5d48e05b1c9a6d8060f58917e3834 + 1;
                end else begin
                    I761983331fb6e3c6c437b3f1660f0b6b  <= I88d5d48e05b1c9a6d8060f58917e3834 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I6804fecdf59233c6cf14409bf2f1e430 != Ie9b2be4c32334220e134e041ca8dfc06[5] ) begin
                    If7f373506cac70f8ba1222db135c27e8  <=  ~I4269e18c2df4d39c683ffb7d01a08322 + 1;
                end else begin
                    If7f373506cac70f8ba1222db135c27e8  <= I4269e18c2df4d39c683ffb7d01a08322 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I6804fecdf59233c6cf14409bf2f1e430 != Ia8a468877c9f96713c8141df9205f92a[7] ) begin
                    I5ce8b2f633011e89356243a1a71edeb6  <=  ~Ia29017fa9327fdaa7c10b2797f8aa6ec + 1;
                end else begin
                    I5ce8b2f633011e89356243a1a71edeb6  <= Ia29017fa9327fdaa7c10b2797f8aa6ec ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I6804fecdf59233c6cf14409bf2f1e430 != Idf0d9dac06522293f8d7e00a93b6bbb5[0] ) begin
                    I70c92e8ada46476d15ef4b3c620d2601  <=  ~Ia142ac799256541fe33f898a6a31dd71 + 1;
                end else begin
                    I70c92e8ada46476d15ef4b3c620d2601  <= Ia142ac799256541fe33f898a6a31dd71 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9e777a342bf53eaba0280737ae404bc1 != If511a6ea6aa5cda5353658d8e192791f[4] ) begin
                    I644e83f0a7d432fba38ffb2d99088eca  <=  ~I4c039794243933a9bb7ad6db7eda6a87 + 1;
                end else begin
                    I644e83f0a7d432fba38ffb2d99088eca  <= I4c039794243933a9bb7ad6db7eda6a87 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9e777a342bf53eaba0280737ae404bc1 != I3c0b6f53f0a5cda5b6758b2ee2c83b92[8] ) begin
                    I73203143fe37933c16fff873c1abf512  <=  ~I0debb3ed4f9540c162cd525588e0ae3f + 1;
                end else begin
                    I73203143fe37933c16fff873c1abf512  <= I0debb3ed4f9540c162cd525588e0ae3f ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9e777a342bf53eaba0280737ae404bc1 != Id6f07dee3e47f39e3b43329c26f690f7[5] ) begin
                    I039f05d5be891a37e04556f1eae674d2  <=  ~I681eed68ee814fb18fd794207d9266e1 + 1;
                end else begin
                    I039f05d5be891a37e04556f1eae674d2  <= I681eed68ee814fb18fd794207d9266e1 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9e777a342bf53eaba0280737ae404bc1 != I4267622319ca65909a3b40484dc74d3a[7] ) begin
                    I8ad3627f171eadcc960a688ac0afcbc0  <=  ~Ic260784b8910f5a0483afee9b68efb31 + 1;
                end else begin
                    I8ad3627f171eadcc960a688ac0afcbc0  <= Ic260784b8910f5a0483afee9b68efb31 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9e777a342bf53eaba0280737ae404bc1 != Id557db735a70dbb14504bc3088e8798e[0] ) begin
                    Ib193b07804d6d5f111b06bda487bfa5f  <=  ~I22cd2d30a7684002cacca4deae4c95a0 + 1;
                end else begin
                    Ib193b07804d6d5f111b06bda487bfa5f  <= I22cd2d30a7684002cacca4deae4c95a0 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ied53820aab06b5c3423b1d878c71948f != Ib0bf69cc797f330fb2546eb46d2d6f76[4] ) begin
                    I51e98035b35a35fdc52f5bab8f19c152  <=  ~I136b4136d582f9fad21f90297cfafea3 + 1;
                end else begin
                    I51e98035b35a35fdc52f5bab8f19c152  <= I136b4136d582f9fad21f90297cfafea3 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ied53820aab06b5c3423b1d878c71948f != I8e591d83170c8ba46d31c61935311b22[8] ) begin
                    Idcada1bfb3c0d1f2a09aab58a2071a57  <=  ~Id8d6be9677d3b0ceca26b3b671757c2c + 1;
                end else begin
                    Idcada1bfb3c0d1f2a09aab58a2071a57  <= Id8d6be9677d3b0ceca26b3b671757c2c ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ied53820aab06b5c3423b1d878c71948f != Ic7f04c065f8ff82c2288f1de77d37189[5] ) begin
                    I94c4e11670b4233fa072517a8f19c901  <=  ~I6a93f928c104ea211dcc8a461506327d + 1;
                end else begin
                    I94c4e11670b4233fa072517a8f19c901  <= I6a93f928c104ea211dcc8a461506327d ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ied53820aab06b5c3423b1d878c71948f != Iedd7d4ea8d082b40244c04946dfb14a0[7] ) begin
                    I09b5273bb15d48a7fd78559930fa6d1c  <=  ~I240da147648bec33195a5f5c273fc6f4 + 1;
                end else begin
                    I09b5273bb15d48a7fd78559930fa6d1c  <= I240da147648bec33195a5f5c273fc6f4 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ied53820aab06b5c3423b1d878c71948f != I150d31ef31093fdfc5f145d84bb35156[0] ) begin
                    I885433b0ab16c6d87abe45af13c9e529  <=  ~I55494d0e8454e3cbb4158559e0d29984 + 1;
                end else begin
                    I885433b0ab16c6d87abe45af13c9e529  <= I55494d0e8454e3cbb4158559e0d29984 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I24cceded372d782c67b33f3a78b16045 != Ib58043c04b5c4c86c1c67e57cc66dcf7[16] ) begin
                    I5ed85845c39337c37791f16e718069b4  <=  ~Ied3cc579b3cf126081acf8e1117007cf + 1;
                end else begin
                    I5ed85845c39337c37791f16e718069b4  <= Ied3cc579b3cf126081acf8e1117007cf ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I24cceded372d782c67b33f3a78b16045 != I19df055705f322292a3601fa63f0e5f9[6] ) begin
                    I1cd93172cf5996bc870063aa642188a2  <=  ~I76140bdc374dd6031097575fd231b468 + 1;
                end else begin
                    I1cd93172cf5996bc870063aa642188a2  <= I76140bdc374dd6031097575fd231b468 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I24cceded372d782c67b33f3a78b16045 != I7e40e6f9d82d9b9fc546672e8e8621bb[0] ) begin
                    I198c055930cb89d0390c336eda8fed4f  <=  ~I650345d21e5c2e7a9bf1810630161089 + 1;
                end else begin
                    I198c055930cb89d0390c336eda8fed4f  <= I650345d21e5c2e7a9bf1810630161089 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I2e78d36bca5bfb016af674c343f9c041 != Ibc0871b3c992fd278815fdbefcd2bac0[16] ) begin
                    I15943aa74e9fbbaebdc0d54eb6a3bffa  <=  ~Ie852635f073dc918e7b1075ffad46f24 + 1;
                end else begin
                    I15943aa74e9fbbaebdc0d54eb6a3bffa  <= Ie852635f073dc918e7b1075ffad46f24 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I2e78d36bca5bfb016af674c343f9c041 != I3d50cfeaa4b69c09bb648b8873a6bc24[6] ) begin
                    Ifb00ae47340bc99669c71da34cccc59e  <=  ~I9ec80c14eb5f0f305e1a9e6107a6001e + 1;
                end else begin
                    Ifb00ae47340bc99669c71da34cccc59e  <= I9ec80c14eb5f0f305e1a9e6107a6001e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I2e78d36bca5bfb016af674c343f9c041 != I14133cbbfa6521c5b81477fa1c229cbf[0] ) begin
                    I688a2c72e69b217d2673e8da75146a83  <=  ~I80ba56447ab19b33610c23105b0b1637 + 1;
                end else begin
                    I688a2c72e69b217d2673e8da75146a83  <= I80ba56447ab19b33610c23105b0b1637 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I17a9a995de58643dbbfb78604f26198b != I8695e1e94cbfcbe4b9eae315b042529e[16] ) begin
                    Ia1a0d8d7dfd6e877f15cce773f85f5b7  <=  ~Ib9132d9fa7180c3fcbacb7c570d6b0f2 + 1;
                end else begin
                    Ia1a0d8d7dfd6e877f15cce773f85f5b7  <= Ib9132d9fa7180c3fcbacb7c570d6b0f2 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I17a9a995de58643dbbfb78604f26198b != I33a6ffad80ddf99a4d316a049078244d[6] ) begin
                    Id4451722e8e2393d627dcd0175dc9903  <=  ~I01621f113f636a9caf9b5ca0bb20ef77 + 1;
                end else begin
                    Id4451722e8e2393d627dcd0175dc9903  <= I01621f113f636a9caf9b5ca0bb20ef77 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I17a9a995de58643dbbfb78604f26198b != I3728e31a7cf48639ce873d9135dc87fb[0] ) begin
                    I3b6fde4ed14cd68af1468ae1d4cc1a22  <=  ~I3eeddb549c6e1f07469c0e0dca68be92 + 1;
                end else begin
                    I3b6fde4ed14cd68af1468ae1d4cc1a22  <= I3eeddb549c6e1f07469c0e0dca68be92 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iad642c4c62766e8f8bd5a1e9e73bdc80 != Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[16] ) begin
                    I57d0920119f8901bd4dea2d5f8fb5d90  <=  ~Ibe664dd203ed4162abcd36eb8d57bfa6 + 1;
                end else begin
                    I57d0920119f8901bd4dea2d5f8fb5d90  <= Ibe664dd203ed4162abcd36eb8d57bfa6 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iad642c4c62766e8f8bd5a1e9e73bdc80 != I980165c1147ac5ff86619c841c6031dc[6] ) begin
                    I80a89644e278e96b1cd1c4b7f764dc34  <=  ~Ia66176893fe306ecfb415d948c50486d + 1;
                end else begin
                    I80a89644e278e96b1cd1c4b7f764dc34  <= Ia66176893fe306ecfb415d948c50486d ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iad642c4c62766e8f8bd5a1e9e73bdc80 != Ic6be12e390bd3c25c66d9b9e7c0532b8[0] ) begin
                    I5d3df1e7563630311f56143ee6d97a8e  <=  ~I8bd4210dcbfc1956381b460fd9ef789b + 1;
                end else begin
                    I5d3df1e7563630311f56143ee6d97a8e  <= I8bd4210dcbfc1956381b460fd9ef789b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I96f92481be1ac6cf985b8ab387d326bf != Iceb64ab2ff8a2e0dfdb74803811d4cfe[18] ) begin
                    Ib57795a63d642a73456324bab41384b6  <=  ~I1ba6328ea9cb7cebcce47d5407d0eae7 + 1;
                end else begin
                    Ib57795a63d642a73456324bab41384b6  <= I1ba6328ea9cb7cebcce47d5407d0eae7 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I96f92481be1ac6cf985b8ab387d326bf != Iec7404bc79c58d4d2538fcdf659e9134[5] ) begin
                    I2370042234b0e93bb66e44b97fca3e43  <=  ~I9e79c17bd782bb7981b4a3623baf96a1 + 1;
                end else begin
                    I2370042234b0e93bb66e44b97fca3e43  <= I9e79c17bd782bb7981b4a3623baf96a1 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I96f92481be1ac6cf985b8ab387d326bf != I82e0e091fba6f79cef97eacac4b43ecb[8] ) begin
                    Ia86740e870d8063f0266b68ad6d7481d  <=  ~I7c6f64d73ff9c6e7f2ed69713e056a2b + 1;
                end else begin
                    Ia86740e870d8063f0266b68ad6d7481d  <= I7c6f64d73ff9c6e7f2ed69713e056a2b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I96f92481be1ac6cf985b8ab387d326bf != Icc50e1923274729fe472ca578b68c0f5[0] ) begin
                    I90a7ea789d3bf7f9126c786474a56da0  <=  ~I00b962a9bf04b62244591051d2dfdbbd + 1;
                end else begin
                    I90a7ea789d3bf7f9126c786474a56da0  <= I00b962a9bf04b62244591051d2dfdbbd ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie03c09039ccafb427153d2347c1caea8 != I5b7caaeb34c43e66e8d095a859e708fe[18] ) begin
                    Ia4b671f3360f3ce55db0dc0e4d78ddbe  <=  ~I3a660b57588325989319701026f658e6 + 1;
                end else begin
                    Ia4b671f3360f3ce55db0dc0e4d78ddbe  <= I3a660b57588325989319701026f658e6 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie03c09039ccafb427153d2347c1caea8 != Ie1cd04c7668d3f450c387a6c1ad778c7[5] ) begin
                    Id96e744d9b10dcddd1ae0115ea57a76a  <=  ~Ibae27cccf3f64e8653c1e244e940e421 + 1;
                end else begin
                    Id96e744d9b10dcddd1ae0115ea57a76a  <= Ibae27cccf3f64e8653c1e244e940e421 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie03c09039ccafb427153d2347c1caea8 != I04302edb2671c5bc0ca2673cd53935e1[8] ) begin
                    I4d226dd2f0bfcdbea6a2e6a6613c1b64  <=  ~I27b89a5001312b2aa48fe385d8a52063 + 1;
                end else begin
                    I4d226dd2f0bfcdbea6a2e6a6613c1b64  <= I27b89a5001312b2aa48fe385d8a52063 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie03c09039ccafb427153d2347c1caea8 != I4d98064f544a41b977ba945d2eecdf21[0] ) begin
                    I5029424c9d9fe923eeb858b1e62cd758  <=  ~Ic6a7476db711a812d146331c562ca7c9 + 1;
                end else begin
                    I5029424c9d9fe923eeb858b1e62cd758  <= Ic6a7476db711a812d146331c562ca7c9 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie7381a8294b4cdf669b9c57cfe4012b5 != I61f0c04673dfb262ef6912eb2df39120[18] ) begin
                    I992e7c551b4aa818606c3465d33eb798  <=  ~I01ca07fe91b5f1edf87300b3583e77c5 + 1;
                end else begin
                    I992e7c551b4aa818606c3465d33eb798  <= I01ca07fe91b5f1edf87300b3583e77c5 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie7381a8294b4cdf669b9c57cfe4012b5 != If511a6ea6aa5cda5353658d8e192791f[5] ) begin
                    I97f2b15ce0a74e68d5a4438111adcb0a  <=  ~I6da707fd74249175d1f68dccb66390c0 + 1;
                end else begin
                    I97f2b15ce0a74e68d5a4438111adcb0a  <= I6da707fd74249175d1f68dccb66390c0 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie7381a8294b4cdf669b9c57cfe4012b5 != I480a0f6d6c3eb936de10a72749f6cd3f[8] ) begin
                    Ia0886ce792e062e22d0c224158cdfb7d  <=  ~I0ae62aae426b75b06d95c46baf33f08e + 1;
                end else begin
                    Ia0886ce792e062e22d0c224158cdfb7d  <= I0ae62aae426b75b06d95c46baf33f08e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie7381a8294b4cdf669b9c57cfe4012b5 != I12f2a9f1e3e715d7e684ff39dd7942f0[0] ) begin
                    I1e805c70d50c2765b4a03ad2982dc421  <=  ~Iec512b5870f295a50921e7e0289a7d35 + 1;
                end else begin
                    I1e805c70d50c2765b4a03ad2982dc421  <= Iec512b5870f295a50921e7e0289a7d35 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I61c9e3f8e42f869f4c9c1386325100b3 != Ibeb5edab51cd6aedad9c2ecedaded6f5[18] ) begin
                    Id9b9a8fe43992ec0793845715dd2226c  <=  ~I3aac84acd9d78070472b1cbc745c80a7 + 1;
                end else begin
                    Id9b9a8fe43992ec0793845715dd2226c  <= I3aac84acd9d78070472b1cbc745c80a7 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I61c9e3f8e42f869f4c9c1386325100b3 != Ib0bf69cc797f330fb2546eb46d2d6f76[5] ) begin
                    Ia6a7f9beaceb08d81012f0e72171252f  <=  ~Ibbb900f56de318bf6e65b49791835ef4 + 1;
                end else begin
                    Ia6a7f9beaceb08d81012f0e72171252f  <= Ibbb900f56de318bf6e65b49791835ef4 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I61c9e3f8e42f869f4c9c1386325100b3 != I50976b0051e84b6a42fc1dbabd7d20ae[8] ) begin
                    I0a9a09b0ab43d2a0f1d1d01e13f0333c  <=  ~I2c2ac1e722fba72c759f1d37b88a9a10 + 1;
                end else begin
                    I0a9a09b0ab43d2a0f1d1d01e13f0333c  <= I2c2ac1e722fba72c759f1d37b88a9a10 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I61c9e3f8e42f869f4c9c1386325100b3 != Iaa4e3c53a0d55e8f42f60ff40893427e[0] ) begin
                    Iba58175a7fd5c5da650222193caff0b3  <=  ~Ida0a18f1b79aff4ddf0e8f7e27794674 + 1;
                end else begin
                    Iba58175a7fd5c5da650222193caff0b3  <= Ida0a18f1b79aff4ddf0e8f7e27794674 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I24c5b2de59eb1f43fe1efe687231c4b7 != I8695e1e94cbfcbe4b9eae315b042529e[17] ) begin
                    I5dd29fd1a73df5662d2b636e7285bad9  <=  ~I9f2029db42c5a968b370587c958c8929 + 1;
                end else begin
                    I5dd29fd1a73df5662d2b636e7285bad9  <= I9f2029db42c5a968b370587c958c8929 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I24c5b2de59eb1f43fe1efe687231c4b7 != I9ef21ef20099af28d9a8c794f70d45a5[4] ) begin
                    I7c19a79f441ecbb73685db5a505e7479  <=  ~If5755f4f61a89d91a91188c17ff5dc5a + 1;
                end else begin
                    I7c19a79f441ecbb73685db5a505e7479  <= If5755f4f61a89d91a91188c17ff5dc5a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I24c5b2de59eb1f43fe1efe687231c4b7 != I26aae317b0b320df86ca4004f64aab88[0] ) begin
                    I7401a0501ba69c5559fbf00c77e58dc5  <=  ~I4419d97c3174ee4610eb6ee9c06cb256 + 1;
                end else begin
                    I7401a0501ba69c5559fbf00c77e58dc5  <= I4419d97c3174ee4610eb6ee9c06cb256 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I43d43acde5f831fc32b7bf5f10b9b3a9 != Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[17] ) begin
                    I89537301987d6da0dbe6cff3caab3ff4  <=  ~Ia964f83676273055e20a2f63c8fffa0d + 1;
                end else begin
                    I89537301987d6da0dbe6cff3caab3ff4  <= Ia964f83676273055e20a2f63c8fffa0d ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I43d43acde5f831fc32b7bf5f10b9b3a9 != Ic2941d16ae6a5cbce70e8546a18ca4ff[4] ) begin
                    I9aaa036a6158d11c235bdc8406d79f4c  <=  ~Iab4fbc811e87df1d1f5821ea732b6a93 + 1;
                end else begin
                    I9aaa036a6158d11c235bdc8406d79f4c  <= Iab4fbc811e87df1d1f5821ea732b6a93 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I43d43acde5f831fc32b7bf5f10b9b3a9 != I9344825cc2e5864f691043a1f94f86a4[0] ) begin
                    Idd9f7ea657ea9cdcb45a7e4b573b9d50  <=  ~I4fbefbb10724b0844c95e85495d4a87f + 1;
                end else begin
                    Idd9f7ea657ea9cdcb45a7e4b573b9d50  <= I4fbefbb10724b0844c95e85495d4a87f ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib06e93161fc8ca3be232f4261b04feb1 != Ib58043c04b5c4c86c1c67e57cc66dcf7[17] ) begin
                    I89013d61c1ea8da8b1c6071cc21c316f  <=  ~I717217d0b5a526f04c7f5ab0835dd5c7 + 1;
                end else begin
                    I89013d61c1ea8da8b1c6071cc21c316f  <= I717217d0b5a526f04c7f5ab0835dd5c7 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib06e93161fc8ca3be232f4261b04feb1 != I8e29ebe9ee25ea8ef3e52ff56fc29157[4] ) begin
                    I1f00849ea055a7893df386aed162a7b6  <=  ~I235937b643e8f2848116dc76c43f47a7 + 1;
                end else begin
                    I1f00849ea055a7893df386aed162a7b6  <= I235937b643e8f2848116dc76c43f47a7 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib06e93161fc8ca3be232f4261b04feb1 != I82988c3879c1de76fe2140c469f6a4c1[0] ) begin
                    I53f275395dd6be17961a5edc3e8da7f2  <=  ~I7481f17d659cce5b4c72a68a9f6be67f + 1;
                end else begin
                    I53f275395dd6be17961a5edc3e8da7f2  <= I7481f17d659cce5b4c72a68a9f6be67f ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ia0dd00f83afc805036f2c6a0e38f725e != Ibc0871b3c992fd278815fdbefcd2bac0[17] ) begin
                    I6ac24c46319a787daa5c545de8c6eeea  <=  ~I5715c21c80992a61bff8aabc3f80415b + 1;
                end else begin
                    I6ac24c46319a787daa5c545de8c6eeea  <= I5715c21c80992a61bff8aabc3f80415b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ia0dd00f83afc805036f2c6a0e38f725e != Ic3742290179b27b9865f9d1f88d66266[4] ) begin
                    If4d5b48882e9e628cf51ad2ac2f38c22  <=  ~I434e3216a615eb46be5c26ef914b9cd2 + 1;
                end else begin
                    If4d5b48882e9e628cf51ad2ac2f38c22  <= I434e3216a615eb46be5c26ef914b9cd2 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ia0dd00f83afc805036f2c6a0e38f725e != I6bdd8334512c7c6a3226ebb4e928a270[0] ) begin
                    Icab010d78cd66b02e089c74f04bf4e75  <=  ~I918326ac0a744d234d74e2c08cf41eb4 + 1;
                end else begin
                    Icab010d78cd66b02e089c74f04bf4e75  <= I918326ac0a744d234d74e2c08cf41eb4 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib0a0f924fe3757a1e0aade7017ad9277 != If511a6ea6aa5cda5353658d8e192791f[6] ) begin
                    I84c88b631bed5311cb6e99e58941149e  <=  ~I966706d314f4c0a7ec842dd699d34926 + 1;
                end else begin
                    I84c88b631bed5311cb6e99e58941149e  <= I966706d314f4c0a7ec842dd699d34926 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib0a0f924fe3757a1e0aade7017ad9277 != I04302edb2671c5bc0ca2673cd53935e1[9] ) begin
                    I5c942076b173cf527e1be2ddb8560e84  <=  ~I5a7d246d88ef12e999f4bdee40e5a585 + 1;
                end else begin
                    I5c942076b173cf527e1be2ddb8560e84  <= I5a7d246d88ef12e999f4bdee40e5a585 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib0a0f924fe3757a1e0aade7017ad9277 != I3c0b6f53f0a5cda5b6758b2ee2c83b92[9] ) begin
                    Ibed2a63af723a7abf96dacf1951e5266  <=  ~Ic2dfaf65c4e17a8dcd55f766c314d6ef + 1;
                end else begin
                    Ibed2a63af723a7abf96dacf1951e5266  <= Ic2dfaf65c4e17a8dcd55f766c314d6ef ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib0a0f924fe3757a1e0aade7017ad9277 != I07930a807994815de45864af579902c4[7] ) begin
                    I242a30bdc8699d8ff550b25dd53d6c59  <=  ~I151831ba6bd0e162275c84815e3c0f12 + 1;
                end else begin
                    I242a30bdc8699d8ff550b25dd53d6c59  <= I151831ba6bd0e162275c84815e3c0f12 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib0a0f924fe3757a1e0aade7017ad9277 != I0debec6ace7160558cce7f111dd1bea6[0] ) begin
                    I376a48b7e0195a5aacc76a0ad8bd14b2  <=  ~I5a8f1675234ebed14d719344b530bbd7 + 1;
                end else begin
                    I376a48b7e0195a5aacc76a0ad8bd14b2  <= I5a8f1675234ebed14d719344b530bbd7 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I1ca949071d734d230cdb8adda46c9d79 != Ib0bf69cc797f330fb2546eb46d2d6f76[6] ) begin
                    I21b062856ced09cb9131c01b5e166f32  <=  ~I95dce76a8d0e729d40fb3f573cfc06ad + 1;
                end else begin
                    I21b062856ced09cb9131c01b5e166f32  <= I95dce76a8d0e729d40fb3f573cfc06ad ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I1ca949071d734d230cdb8adda46c9d79 != I480a0f6d6c3eb936de10a72749f6cd3f[9] ) begin
                    I6b3cd79aa87235ff174c0299b855dd3d  <=  ~I6c26c7918254426c18f2e747c91438c5 + 1;
                end else begin
                    I6b3cd79aa87235ff174c0299b855dd3d  <= I6c26c7918254426c18f2e747c91438c5 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I1ca949071d734d230cdb8adda46c9d79 != I8e591d83170c8ba46d31c61935311b22[9] ) begin
                    I814b62120953991f9da055f118967e05  <=  ~I0414ead2472e42da8a271cb0bd1debf4 + 1;
                end else begin
                    I814b62120953991f9da055f118967e05  <= I0414ead2472e42da8a271cb0bd1debf4 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I1ca949071d734d230cdb8adda46c9d79 != I72a2f42b727a0503d43332c0f22d5ae3[7] ) begin
                    I3f33901c407a87e10d86c13c83dd52eb  <=  ~Ic6a6f5090470a76ddb7315c022ddc104 + 1;
                end else begin
                    I3f33901c407a87e10d86c13c83dd52eb  <= Ic6a6f5090470a76ddb7315c022ddc104 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I1ca949071d734d230cdb8adda46c9d79 != I8ee02e65ce9183683f0f3168bfd755c5[0] ) begin
                    I241622b0367dde514f96ece55c8c3964  <=  ~I2a00ee56a5aa639f45eb3b1bdcffe81c + 1;
                end else begin
                    I241622b0367dde514f96ece55c8c3964  <= I2a00ee56a5aa639f45eb3b1bdcffe81c ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I40170922c652fa7fa42abc6f580b5e3d != Iec7404bc79c58d4d2538fcdf659e9134[6] ) begin
                    If9efe7a1c359ec03014a52870ac13aec  <=  ~Ibceb2b824cd4bc10bb06ee8adc693bd1 + 1;
                end else begin
                    If9efe7a1c359ec03014a52870ac13aec  <= Ibceb2b824cd4bc10bb06ee8adc693bd1 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I40170922c652fa7fa42abc6f580b5e3d != I50976b0051e84b6a42fc1dbabd7d20ae[9] ) begin
                    Ibc73d07e0c97a6fcae791e04106cb082  <=  ~Ia8b9f373fe68ac4cbca35e04376e3cca + 1;
                end else begin
                    Ibc73d07e0c97a6fcae791e04106cb082  <= Ia8b9f373fe68ac4cbca35e04376e3cca ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I40170922c652fa7fa42abc6f580b5e3d != I02b62fafd371de339f299f8aefec6c43[9] ) begin
                    I2f3ab9654e515a54e22e73d6c130ccc3  <=  ~I5d1a89e85f6609b469e73e15aeffcbc4 + 1;
                end else begin
                    I2f3ab9654e515a54e22e73d6c130ccc3  <= I5d1a89e85f6609b469e73e15aeffcbc4 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I40170922c652fa7fa42abc6f580b5e3d != I8b8b9c4777e6df3eb2b9313e69ef2c8c[7] ) begin
                    Idf6875955525d80dc660ce956f4a84e7  <=  ~I677fe06bad241bc8dd6a65a97f6db520 + 1;
                end else begin
                    Idf6875955525d80dc660ce956f4a84e7  <= I677fe06bad241bc8dd6a65a97f6db520 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I40170922c652fa7fa42abc6f580b5e3d != I80e6d2c9c5f7b6bc6bffa063c4959115[0] ) begin
                    If94a1abfb972f63629d07e64dc23863c  <=  ~If3c0f892fd71eb0ed8d1f70b4b33450b + 1;
                end else begin
                    If94a1abfb972f63629d07e64dc23863c  <= If3c0f892fd71eb0ed8d1f70b4b33450b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib1ad0b531ac9028971d68f533e7ae566 != Ie1cd04c7668d3f450c387a6c1ad778c7[6] ) begin
                    I0c0060fe260afa3cdc72f35ffb6938ff  <=  ~Ic65f0f75f56bf85122a89cdf07e98152 + 1;
                end else begin
                    I0c0060fe260afa3cdc72f35ffb6938ff  <= Ic65f0f75f56bf85122a89cdf07e98152 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib1ad0b531ac9028971d68f533e7ae566 != I82e0e091fba6f79cef97eacac4b43ecb[9] ) begin
                    I6627bcdbaa8afb115123777abd45435b  <=  ~I41d22bafaf58e4a6de04640864653a16 + 1;
                end else begin
                    I6627bcdbaa8afb115123777abd45435b  <= I41d22bafaf58e4a6de04640864653a16 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib1ad0b531ac9028971d68f533e7ae566 != I0e0b15868b02ca52b260f17f150d237e[9] ) begin
                    I70d32affde22f9dcb2d77430fca39069  <=  ~I06a46b86f6edede0f5f72658a19910b7 + 1;
                end else begin
                    I70d32affde22f9dcb2d77430fca39069  <= I06a46b86f6edede0f5f72658a19910b7 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib1ad0b531ac9028971d68f533e7ae566 != I4a16e8e7946d9a8220304fc1be3fb362[7] ) begin
                    I76060709de3ea188748849f043c59ac0  <=  ~I8591d0399594adacfeb006c5195c2c71 + 1;
                end else begin
                    I76060709de3ea188748849f043c59ac0  <= I8591d0399594adacfeb006c5195c2c71 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib1ad0b531ac9028971d68f533e7ae566 != I0f21fb041239a7a8895c9506f2754595[0] ) begin
                    I07b9b1f4fa01b16cc69356057d3b6154  <=  ~Id90588b5f82cd32e801fbea04d24e4a5 + 1;
                end else begin
                    I07b9b1f4fa01b16cc69356057d3b6154  <= Id90588b5f82cd32e801fbea04d24e4a5 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I0ab0170c7ceffbb58377b65d2ad92093 != Iceb64ab2ff8a2e0dfdb74803811d4cfe[19] ) begin
                    Iabf572c97b48c6a7dcc19e56676e3a82  <=  ~Ib642d757fae818cd6d713ffb6ce18fc1 + 1;
                end else begin
                    Iabf572c97b48c6a7dcc19e56676e3a82  <= Ib642d757fae818cd6d713ffb6ce18fc1 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I0ab0170c7ceffbb58377b65d2ad92093 != Iedd7d4ea8d082b40244c04946dfb14a0[8] ) begin
                    I5814a85c45fd0f7be21ed325235fe4b7  <=  ~Id76bff2a12cf792e52ccc463647334c0 + 1;
                end else begin
                    I5814a85c45fd0f7be21ed325235fe4b7  <= Id76bff2a12cf792e52ccc463647334c0 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I0ab0170c7ceffbb58377b65d2ad92093 != I8ce37a8e81b54043276835c11e394df5[0] ) begin
                    I2288a6ad3b748b716249f4adc42d52c4  <=  ~I92ffa890ed6d83d4fc543504e4d421c1 + 1;
                end else begin
                    I2288a6ad3b748b716249f4adc42d52c4  <= I92ffa890ed6d83d4fc543504e4d421c1 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9ac68f228a93bbf4aa4a559b1364e42e != I5b7caaeb34c43e66e8d095a859e708fe[19] ) begin
                    I60cbd4369e7ba9b6532f279e5c59084c  <=  ~Ifc4a65edeaf630b3d29437bcd6c20121 + 1;
                end else begin
                    I60cbd4369e7ba9b6532f279e5c59084c  <= Ifc4a65edeaf630b3d29437bcd6c20121 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9ac68f228a93bbf4aa4a559b1364e42e != I56e1fe0c7a62589c123876f2b4e57a26[8] ) begin
                    I95361d5f524ccb9feb42811af5c482e2  <=  ~Id57a11f56fc223501a9b68b8b05ebd3e + 1;
                end else begin
                    I95361d5f524ccb9feb42811af5c482e2  <= Id57a11f56fc223501a9b68b8b05ebd3e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9ac68f228a93bbf4aa4a559b1364e42e != Idf7d1f78735ce1e9695d99a532a7726e[0] ) begin
                    I022df337bcc05ac5648b8ae2e42f3a76  <=  ~I522ba8bfc1949337e8befe82cc1e86e6 + 1;
                end else begin
                    I022df337bcc05ac5648b8ae2e42f3a76  <= I522ba8bfc1949337e8befe82cc1e86e6 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I375c5f7eac92d853e85e0606011f3fb0 != I61f0c04673dfb262ef6912eb2df39120[19] ) begin
                    I2ead0e9941e2280309ab53535b1e1ac1  <=  ~I7153e27c44ebbc2f04e9ba03cf09b5e1 + 1;
                end else begin
                    I2ead0e9941e2280309ab53535b1e1ac1  <= I7153e27c44ebbc2f04e9ba03cf09b5e1 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I375c5f7eac92d853e85e0606011f3fb0 != Ia8a468877c9f96713c8141df9205f92a[8] ) begin
                    I3e5139f24e3d082eb31b0e61ea9fa1aa  <=  ~Id15e4b4f186ec863f12a54acd8ef8963 + 1;
                end else begin
                    I3e5139f24e3d082eb31b0e61ea9fa1aa  <= Id15e4b4f186ec863f12a54acd8ef8963 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I375c5f7eac92d853e85e0606011f3fb0 != I96a552ed2d18c0ba3fc6cb6d6b6a0f44[0] ) begin
                    I60d9a7f95fb8623753002ecaf9a4efcc  <=  ~I95c77eec7575cd7aa93a36f31ea635a2 + 1;
                end else begin
                    I60d9a7f95fb8623753002ecaf9a4efcc  <= I95c77eec7575cd7aa93a36f31ea635a2 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I94f9b1f2e63748c21ec7222c9641366a != Ibeb5edab51cd6aedad9c2ecedaded6f5[19] ) begin
                    I93b69bfb228db4b569a6772179d603be  <=  ~I3c8114dbe0658cc2889c787f1366abfa + 1;
                end else begin
                    I93b69bfb228db4b569a6772179d603be  <= I3c8114dbe0658cc2889c787f1366abfa ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I94f9b1f2e63748c21ec7222c9641366a != I4267622319ca65909a3b40484dc74d3a[8] ) begin
                    I85c4d3d6c8408c6f38741257ed177ca6  <=  ~Ieacf971e9e10fb73c7df9f1da8372f30 + 1;
                end else begin
                    I85c4d3d6c8408c6f38741257ed177ca6  <= Ieacf971e9e10fb73c7df9f1da8372f30 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I94f9b1f2e63748c21ec7222c9641366a != I3c76936e8e3467378210a13645a401d4[0] ) begin
                    I23a74ea5e7174d95e6d16a5e85ac236b  <=  ~I35de1b03ea865f2c6381ce73e03dc220 + 1;
                end else begin
                    I23a74ea5e7174d95e6d16a5e85ac236b  <= I35de1b03ea865f2c6381ce73e03dc220 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I55500c1d85c4970932be67cc5cd2e023 != I8695e1e94cbfcbe4b9eae315b042529e[18] ) begin
                    Ide530e6f4622c8a7b101b6dce9650e42  <=  ~Idec12e02904ea98c7580919584f2dba1 + 1;
                end else begin
                    Ide530e6f4622c8a7b101b6dce9650e42  <= Idec12e02904ea98c7580919584f2dba1 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I55500c1d85c4970932be67cc5cd2e023 != I04302edb2671c5bc0ca2673cd53935e1[10] ) begin
                    Ic95191bccb18e26c10e56be395ca6b1a  <=  ~Ia370c83631a2c1bbf39c7264deafafb5 + 1;
                end else begin
                    Ic95191bccb18e26c10e56be395ca6b1a  <= Ia370c83631a2c1bbf39c7264deafafb5 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I55500c1d85c4970932be67cc5cd2e023 != Id6f07dee3e47f39e3b43329c26f690f7[6] ) begin
                    Id0f75e19b94541ed5c5c352d13390d2d  <=  ~I05b4a07dfc0d2695eae34bea4c1c6565 + 1;
                end else begin
                    Id0f75e19b94541ed5c5c352d13390d2d  <= I05b4a07dfc0d2695eae34bea4c1c6565 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I55500c1d85c4970932be67cc5cd2e023 != Ic9a1d599fcfd5dd51265e5d0989719b6[0] ) begin
                    Ie697d28d757df82b3901564bda43251c  <=  ~If1ecdc27e3419dd1434e403f237c2b58 + 1;
                end else begin
                    Ie697d28d757df82b3901564bda43251c  <= If1ecdc27e3419dd1434e403f237c2b58 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I36b487cd1a57a3a503e587fdefbb19e4 != Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[18] ) begin
                    Iaf0bbbe791bb71d0f557dc71caa5fb87  <=  ~I039c552777d0fb40bebcdd2d4a3394c2 + 1;
                end else begin
                    Iaf0bbbe791bb71d0f557dc71caa5fb87  <= I039c552777d0fb40bebcdd2d4a3394c2 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I36b487cd1a57a3a503e587fdefbb19e4 != I480a0f6d6c3eb936de10a72749f6cd3f[10] ) begin
                    Ie4ae993ddb776bdffec843db0def2f5c  <=  ~Iaa52fb63184514b6d754bcc896235150 + 1;
                end else begin
                    Ie4ae993ddb776bdffec843db0def2f5c  <= Iaa52fb63184514b6d754bcc896235150 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I36b487cd1a57a3a503e587fdefbb19e4 != Ic7f04c065f8ff82c2288f1de77d37189[6] ) begin
                    I4dca2dd40a7127ce44f83b430a34c738  <=  ~Ied9781e625c1fa8741853dd6b8b3a9e7 + 1;
                end else begin
                    I4dca2dd40a7127ce44f83b430a34c738  <= Ied9781e625c1fa8741853dd6b8b3a9e7 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I36b487cd1a57a3a503e587fdefbb19e4 != I60156470e631268c392040d3c5582eca[0] ) begin
                    I8572aedc94f7243ce5eacb332c81eae2  <=  ~I767272262e9d2e85dba1aa93f578f25c + 1;
                end else begin
                    I8572aedc94f7243ce5eacb332c81eae2  <= I767272262e9d2e85dba1aa93f578f25c ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Icb5350e8c55a2adb370078a7575e28f8 != Ib58043c04b5c4c86c1c67e57cc66dcf7[18] ) begin
                    I4102100fa5f1dd299af0190862efcc42  <=  ~Ib3b4cd6d8ab17869a2278552c02635c8 + 1;
                end else begin
                    I4102100fa5f1dd299af0190862efcc42  <= Ib3b4cd6d8ab17869a2278552c02635c8 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Icb5350e8c55a2adb370078a7575e28f8 != I50976b0051e84b6a42fc1dbabd7d20ae[10] ) begin
                    I224bbdf94ac86c5c376d1db4f4d4e060  <=  ~Ie7a5cb2ecb3fce35825785b9bca6b3bd + 1;
                end else begin
                    I224bbdf94ac86c5c376d1db4f4d4e060  <= Ie7a5cb2ecb3fce35825785b9bca6b3bd ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Icb5350e8c55a2adb370078a7575e28f8 != Ieb244944e7ee8236a207924f56fbc689[6] ) begin
                    I6d83efa9f988328f487e9232bf2633a2  <=  ~Ib9a0f8efd3dad427f247ce90fdfb94a4 + 1;
                end else begin
                    I6d83efa9f988328f487e9232bf2633a2  <= Ib9a0f8efd3dad427f247ce90fdfb94a4 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Icb5350e8c55a2adb370078a7575e28f8 != I821126d1516ad7e8191a7b2a3b5e4b47[0] ) begin
                    I6734123aaf6320da75638b212812732f  <=  ~I69a221a1bd95a588aa74b9bed0357762 + 1;
                end else begin
                    I6734123aaf6320da75638b212812732f  <= I69a221a1bd95a588aa74b9bed0357762 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I8a7a31327c9e4cbd88ce39fea8971caf != Ibc0871b3c992fd278815fdbefcd2bac0[18] ) begin
                    I52403a0454e5fa002e79eaab7ea497bd  <=  ~I64f125cf2ca6a6da8a9cdae9e246c24a + 1;
                end else begin
                    I52403a0454e5fa002e79eaab7ea497bd  <= I64f125cf2ca6a6da8a9cdae9e246c24a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I8a7a31327c9e4cbd88ce39fea8971caf != I82e0e091fba6f79cef97eacac4b43ecb[10] ) begin
                    I96fe3eb633eff6958ac575b997460bb9  <=  ~Ifac9dd60dd6c543aa94b39c599f0819a + 1;
                end else begin
                    I96fe3eb633eff6958ac575b997460bb9  <= Ifac9dd60dd6c543aa94b39c599f0819a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I8a7a31327c9e4cbd88ce39fea8971caf != Ie9b2be4c32334220e134e041ca8dfc06[6] ) begin
                    I69f563e7b7ad483893ac9c4684349769  <=  ~Icf062382a1e462571569ccee75b0a3ee + 1;
                end else begin
                    I69f563e7b7ad483893ac9c4684349769  <= Icf062382a1e462571569ccee75b0a3ee ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I8a7a31327c9e4cbd88ce39fea8971caf != Ibe72e9f6d2c3cbbcf98f6b5aa6a4f93b[0] ) begin
                    I7f6dc6f0f403c58f9aaaa70c2383a666  <=  ~Ieed8b94295bed265961c4f52c3379914 + 1;
                end else begin
                    I7f6dc6f0f403c58f9aaaa70c2383a666  <= Ieed8b94295bed265961c4f52c3379914 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ied069655ed3775819d0bcb722d6d0488 != Ib0bf69cc797f330fb2546eb46d2d6f76[7] ) begin
                    I4f1221ce7880729fe584b42ef3afe6b2  <=  ~I165eabcdde76821fdc308ff7a8c6d2ea + 1;
                end else begin
                    I4f1221ce7880729fe584b42ef3afe6b2  <= I165eabcdde76821fdc308ff7a8c6d2ea ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ied069655ed3775819d0bcb722d6d0488 != I0e0b15868b02ca52b260f17f150d237e[10] ) begin
                    Ic08e85346f61da036a15345a13ac12f0  <=  ~I8b3542a6d64d6a7ebba4124bc6702f3e + 1;
                end else begin
                    Ic08e85346f61da036a15345a13ac12f0  <= I8b3542a6d64d6a7ebba4124bc6702f3e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ied069655ed3775819d0bcb722d6d0488 != I651d700a00d7004d8728bc7356f30926[6] ) begin
                    I9160d11439c5140c0109b5190eb82e6b  <=  ~I7b68afec199be705d766c169f1ece981 + 1;
                end else begin
                    I9160d11439c5140c0109b5190eb82e6b  <= I7b68afec199be705d766c169f1ece981 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ied069655ed3775819d0bcb722d6d0488 != I1e8b6306d2dfde4a36ee9b9c2caf1c85[0] ) begin
                    I66391978843c39b6acbdb4847a01050a  <=  ~I4b6c8226ef2bc20dbd31d242bdb98b8c + 1;
                end else begin
                    I66391978843c39b6acbdb4847a01050a  <= I4b6c8226ef2bc20dbd31d242bdb98b8c ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I78a5fc80d42e8db1b56cce5f4c97e325 != Iec7404bc79c58d4d2538fcdf659e9134[7] ) begin
                    I6a6eb62960b616043415406ebfc21346  <=  ~Ic3b4a86f22caf5b6103d52b6c9d2a991 + 1;
                end else begin
                    I6a6eb62960b616043415406ebfc21346  <= Ic3b4a86f22caf5b6103d52b6c9d2a991 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I78a5fc80d42e8db1b56cce5f4c97e325 != I3c0b6f53f0a5cda5b6758b2ee2c83b92[10] ) begin
                    Id667c80003b5541de9f84d3b8709c828  <=  ~Ia37592b207086f63e2d94e3d7d26c740 + 1;
                end else begin
                    Id667c80003b5541de9f84d3b8709c828  <= Ia37592b207086f63e2d94e3d7d26c740 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I78a5fc80d42e8db1b56cce5f4c97e325 != Ic2580cbeec8c11a19bd1e2ebc29d255e[6] ) begin
                    Ia030c08757123aae947f86ab8bfb6d94  <=  ~Id0d786026e3ab0ddbffbc20e4d409857 + 1;
                end else begin
                    Ia030c08757123aae947f86ab8bfb6d94  <= Id0d786026e3ab0ddbffbc20e4d409857 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I78a5fc80d42e8db1b56cce5f4c97e325 != I48ed92480f457fc3cc2ff0dd7d177a10[0] ) begin
                    I4f756e4125c8af5c412944b273e01cb0  <=  ~I333837f976cfc7f90ab0a6dcd8c1ce79 + 1;
                end else begin
                    I4f756e4125c8af5c412944b273e01cb0  <= I333837f976cfc7f90ab0a6dcd8c1ce79 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I3ade7e345432319c1a9c91d4068b3ec9 != Ie1cd04c7668d3f450c387a6c1ad778c7[7] ) begin
                    Iaec1f186cb4a65da21d41e637fc628f7  <=  ~Id115b4708a49dcfd167e79ef6993e371 + 1;
                end else begin
                    Iaec1f186cb4a65da21d41e637fc628f7  <= Id115b4708a49dcfd167e79ef6993e371 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I3ade7e345432319c1a9c91d4068b3ec9 != I8e591d83170c8ba46d31c61935311b22[10] ) begin
                    I123a212546a8ac394051425db4924812  <=  ~I666da645400344644e848ee6f7592d3c + 1;
                end else begin
                    I123a212546a8ac394051425db4924812  <= I666da645400344644e848ee6f7592d3c ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I3ade7e345432319c1a9c91d4068b3ec9 != If79ed5ee2b8710da0608c1e245d07d55[6] ) begin
                    I730634ea15ac94d241f3ad2d6393a227  <=  ~Ibafeadd691eee03f855ed657c01022c9 + 1;
                end else begin
                    I730634ea15ac94d241f3ad2d6393a227  <= Ibafeadd691eee03f855ed657c01022c9 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I3ade7e345432319c1a9c91d4068b3ec9 != Iaed28d88a651f0151501ec4ea6ee3346[0] ) begin
                    Id2c9f7ac95de07148c54803f69347f56  <=  ~I10ec5c43a3fb65273053063001307280 + 1;
                end else begin
                    Id2c9f7ac95de07148c54803f69347f56  <= I10ec5c43a3fb65273053063001307280 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I88aed46f6dad7a81006562a720670654 != If511a6ea6aa5cda5353658d8e192791f[7] ) begin
                    I45c5e6710240685bf54b73b0d7a64271  <=  ~I05c778eb3588bdaccf714ba456f534c2 + 1;
                end else begin
                    I45c5e6710240685bf54b73b0d7a64271  <= I05c778eb3588bdaccf714ba456f534c2 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I88aed46f6dad7a81006562a720670654 != I02b62fafd371de339f299f8aefec6c43[10] ) begin
                    Iebdc41368d57498a04fa73e30b10a966  <=  ~Icd11e8d97a6ac6c0a73e8adee1f98c4e + 1;
                end else begin
                    Iebdc41368d57498a04fa73e30b10a966  <= Icd11e8d97a6ac6c0a73e8adee1f98c4e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I88aed46f6dad7a81006562a720670654 != I9497bbb4f746969a95cff948a3ee9ade[6] ) begin
                    I47b878f27c30f79a37e97e022307e9e9  <=  ~If07c2223d4262e22cca9b77c3ed5ee01 + 1;
                end else begin
                    I47b878f27c30f79a37e97e022307e9e9  <= If07c2223d4262e22cca9b77c3ed5ee01 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I88aed46f6dad7a81006562a720670654 != I9d94d9b5414662de841443d7866e66b1[0] ) begin
                    I5061e13a179d27e1ba5f89ce8ee0fd4a  <=  ~If0c8ce0ff66fe2806448f1c819d58ec8 + 1;
                end else begin
                    I5061e13a179d27e1ba5f89ce8ee0fd4a  <= If0c8ce0ff66fe2806448f1c819d58ec8 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I79e574dc9c7e18b695c9a2619b71b995 != Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[19] ) begin
                    Ic7ff9cde71054c1ee9eef81eabdd7061  <=  ~Iccdc2371dfd9fda3e506adc2b1681ba3 + 1;
                end else begin
                    Ic7ff9cde71054c1ee9eef81eabdd7061  <= Iccdc2371dfd9fda3e506adc2b1681ba3 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I79e574dc9c7e18b695c9a2619b71b995 != Ie9b2be4c32334220e134e041ca8dfc06[7] ) begin
                    Ia0a02781c674fe5d769206448d475245  <=  ~I26e61dca9d045c4661b97afe346152c8 + 1;
                end else begin
                    Ia0a02781c674fe5d769206448d475245  <= I26e61dca9d045c4661b97afe346152c8 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I79e574dc9c7e18b695c9a2619b71b995 != I4267622319ca65909a3b40484dc74d3a[9] ) begin
                    Id66c47fd69c175a4393e975a269cf053  <=  ~Id488d650b86f5def0668f4a1ef841b6a + 1;
                end else begin
                    Id66c47fd69c175a4393e975a269cf053  <= Id488d650b86f5def0668f4a1ef841b6a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I79e574dc9c7e18b695c9a2619b71b995 != I870b8a3b11be215a8704ba05568f05e2[0] ) begin
                    I0f7c32fc1548fb49b8041f55c157498a  <=  ~I479365266255d2228ecd86c350e8d38b + 1;
                end else begin
                    I0f7c32fc1548fb49b8041f55c157498a  <= I479365266255d2228ecd86c350e8d38b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I800ef583bec1d46d3d4ffdea6b312ef9 != Ib58043c04b5c4c86c1c67e57cc66dcf7[19] ) begin
                    I4939f69abb1eac56d5021e06406a93b5  <=  ~I08d9c488fd85db45344e649699196263 + 1;
                end else begin
                    I4939f69abb1eac56d5021e06406a93b5  <= I08d9c488fd85db45344e649699196263 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I800ef583bec1d46d3d4ffdea6b312ef9 != Id6f07dee3e47f39e3b43329c26f690f7[7] ) begin
                    Ife1190f76c2e251704c2960c23330a48  <=  ~Icde86d0ead44385b07e9a29057417417 + 1;
                end else begin
                    Ife1190f76c2e251704c2960c23330a48  <= Icde86d0ead44385b07e9a29057417417 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I800ef583bec1d46d3d4ffdea6b312ef9 != Iedd7d4ea8d082b40244c04946dfb14a0[9] ) begin
                    Ib06b60cf9933dd8952206c5f3ccced8e  <=  ~I21feecd24d912ef3d0aec0e375958f3f + 1;
                end else begin
                    Ib06b60cf9933dd8952206c5f3ccced8e  <= I21feecd24d912ef3d0aec0e375958f3f ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I800ef583bec1d46d3d4ffdea6b312ef9 != Ia8bbf21e040b326058a9acb7d198a835[0] ) begin
                    I89ffab735ee30423c82e079ed98216c5  <=  ~I59f419b3bc183a5fe743be3878fac587 + 1;
                end else begin
                    I89ffab735ee30423c82e079ed98216c5  <= I59f419b3bc183a5fe743be3878fac587 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I56cc5cd6d0a5a4e4601fd48e838fdaf3 != Ibc0871b3c992fd278815fdbefcd2bac0[19] ) begin
                    I634f0ce28934600a1a31ab0d8e59b4a9  <=  ~Ib0804d8bdda49ecd0024300eed52be53 + 1;
                end else begin
                    I634f0ce28934600a1a31ab0d8e59b4a9  <= Ib0804d8bdda49ecd0024300eed52be53 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I56cc5cd6d0a5a4e4601fd48e838fdaf3 != Ic7f04c065f8ff82c2288f1de77d37189[7] ) begin
                    I1a24e98165afa62bd14986911a36fb6e  <=  ~I37b0efdee34647a5111d698a5a80f367 + 1;
                end else begin
                    I1a24e98165afa62bd14986911a36fb6e  <= I37b0efdee34647a5111d698a5a80f367 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I56cc5cd6d0a5a4e4601fd48e838fdaf3 != I56e1fe0c7a62589c123876f2b4e57a26[9] ) begin
                    I9c4b34b5fb1d59c132bcaeb6258675df  <=  ~Id382a04e94d0749d0858041bdc5861be + 1;
                end else begin
                    I9c4b34b5fb1d59c132bcaeb6258675df  <= Id382a04e94d0749d0858041bdc5861be ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I56cc5cd6d0a5a4e4601fd48e838fdaf3 != Ie852f207c8f537621b080ffa0a89bfdc[0] ) begin
                    I9494921d8487ee0b314f75cf0380fd2f  <=  ~I368be992a21201268c41506396dcdcf6 + 1;
                end else begin
                    I9494921d8487ee0b314f75cf0380fd2f  <= I368be992a21201268c41506396dcdcf6 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I21047a3955b8b89bdb9013d571b2bd0d != I8695e1e94cbfcbe4b9eae315b042529e[19] ) begin
                    Ibaf00a6780325882067a79f0c4d693d2  <=  ~I603a008893b5196d9f273b47a9d63144 + 1;
                end else begin
                    Ibaf00a6780325882067a79f0c4d693d2  <= I603a008893b5196d9f273b47a9d63144 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I21047a3955b8b89bdb9013d571b2bd0d != Ieb244944e7ee8236a207924f56fbc689[7] ) begin
                    Ic23e01562c8a753fd70c343297be288a  <=  ~Ie70d3a768bc09ddff6ac68aaba7d9f2c + 1;
                end else begin
                    Ic23e01562c8a753fd70c343297be288a  <= Ie70d3a768bc09ddff6ac68aaba7d9f2c ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I21047a3955b8b89bdb9013d571b2bd0d != Ia8a468877c9f96713c8141df9205f92a[9] ) begin
                    I61cc8a0f49e393721a62a776e4793deb  <=  ~Ifb8bd837ada3d8ed5116db29da82d2a9 + 1;
                end else begin
                    I61cc8a0f49e393721a62a776e4793deb  <= Ifb8bd837ada3d8ed5116db29da82d2a9 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I21047a3955b8b89bdb9013d571b2bd0d != If53029b05bea46d656a6ef72fb6d6642[0] ) begin
                    If2b3e7d1541cbd8ffc2b4cfc3ad13a57  <=  ~I978b93d46e20cb3eda70e5a976d62348 + 1;
                end else begin
                    If2b3e7d1541cbd8ffc2b4cfc3ad13a57  <= I978b93d46e20cb3eda70e5a976d62348 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I56eb529a34b484cd20e29958cd6878eb != Ibeb5edab51cd6aedad9c2ecedaded6f5[20] ) begin
                    I71afab29cdb962e1f1ca21b61dfb50c6  <=  ~Ib404040d4fb58f47f245184c3be01789 + 1;
                end else begin
                    I71afab29cdb962e1f1ca21b61dfb50c6  <= Ib404040d4fb58f47f245184c3be01789 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I56eb529a34b484cd20e29958cd6878eb != I04302edb2671c5bc0ca2673cd53935e1[11] ) begin
                    Ia284f974dd8a526f31eb81ed71a06e94  <=  ~I9c664265c53ebffaad097b70ff3cbbce + 1;
                end else begin
                    Ia284f974dd8a526f31eb81ed71a06e94  <= I9c664265c53ebffaad097b70ff3cbbce ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I56eb529a34b484cd20e29958cd6878eb != I872f61d20baf011e867b44dc5539fc37[13] ) begin
                    I3e3ce8b4ead150a6eae2e5c701c7b598  <=  ~I781306c6b1ce0741d9c2fa06865f7a19 + 1;
                end else begin
                    I3e3ce8b4ead150a6eae2e5c701c7b598  <= I781306c6b1ce0741d9c2fa06865f7a19 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I56eb529a34b484cd20e29958cd6878eb != I8e8a740d09e000444ba1f4931b5cccf4[0] ) begin
                    Idf3d79da44f2d686f5bd43c3c1427430  <=  ~I16fa2e3dc0b3eddbc72811b51d6ac8ed + 1;
                end else begin
                    Idf3d79da44f2d686f5bd43c3c1427430  <= I16fa2e3dc0b3eddbc72811b51d6ac8ed ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I74588df6399af2c1112e3fa557e89e17 != Iceb64ab2ff8a2e0dfdb74803811d4cfe[20] ) begin
                    Iefd370d0df1a93639af482f78a1e8706  <=  ~Ia6f232495726806d01b702b0e248b2f2 + 1;
                end else begin
                    Iefd370d0df1a93639af482f78a1e8706  <= Ia6f232495726806d01b702b0e248b2f2 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I74588df6399af2c1112e3fa557e89e17 != I480a0f6d6c3eb936de10a72749f6cd3f[11] ) begin
                    I3ed2da9b53daac0852a06ad1acfad21b  <=  ~I66b3734060600caa45d699508c5083d2 + 1;
                end else begin
                    I3ed2da9b53daac0852a06ad1acfad21b  <= I66b3734060600caa45d699508c5083d2 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I74588df6399af2c1112e3fa557e89e17 != I6f5c991e5fdcf56d582c6f80eb6731df[13] ) begin
                    I453fdf4fbb5af5bd28a20d7643da9eb2  <=  ~I85fae6b23d086235a94a0162e2fb5310 + 1;
                end else begin
                    I453fdf4fbb5af5bd28a20d7643da9eb2  <= I85fae6b23d086235a94a0162e2fb5310 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I74588df6399af2c1112e3fa557e89e17 != I46605d823e06af5485e50b256b5c3f22[0] ) begin
                    If8125ad3c9e7f0a2b84106064d320996  <=  ~I8d6443d1be42203cb834345ae7e5aff5 + 1;
                end else begin
                    If8125ad3c9e7f0a2b84106064d320996  <= I8d6443d1be42203cb834345ae7e5aff5 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ic8eae1a92f46db040eb22d726c3a0e6d != I5b7caaeb34c43e66e8d095a859e708fe[20] ) begin
                    Ifb6c65a00d9a2c31d8b1119b949828d8  <=  ~I717332b7f76e9caf9351f1aa69b72a12 + 1;
                end else begin
                    Ifb6c65a00d9a2c31d8b1119b949828d8  <= I717332b7f76e9caf9351f1aa69b72a12 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ic8eae1a92f46db040eb22d726c3a0e6d != I50976b0051e84b6a42fc1dbabd7d20ae[11] ) begin
                    I43f2b69c6b427de3095c44d4166b77cd  <=  ~Ieebd34db071409288f489129b70ab599 + 1;
                end else begin
                    I43f2b69c6b427de3095c44d4166b77cd  <= Ieebd34db071409288f489129b70ab599 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ic8eae1a92f46db040eb22d726c3a0e6d != Ia5cc3055ba3365e64cf59c4d4fd3f093[13] ) begin
                    Ie9cce5746a83479a567bbaeac6dbf497  <=  ~I917c874137d64a9a495335c8f8ef5374 + 1;
                end else begin
                    Ie9cce5746a83479a567bbaeac6dbf497  <= I917c874137d64a9a495335c8f8ef5374 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ic8eae1a92f46db040eb22d726c3a0e6d != I38344d68127f5c035193bb9030ce4d4d[0] ) begin
                    Ic9018b88fa91fb638bbab0613795ae13  <=  ~I15fb4fb838d4a614c468f7d49261bda3 + 1;
                end else begin
                    Ic9018b88fa91fb638bbab0613795ae13  <= I15fb4fb838d4a614c468f7d49261bda3 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I854a15bc7e9728b01c9a1960f6248dc9 != I61f0c04673dfb262ef6912eb2df39120[20] ) begin
                    I56873feb8418005b5661c7382f2dbeec  <=  ~I2eb093d2a38ba8cf4be47d1d7f54ecc4 + 1;
                end else begin
                    I56873feb8418005b5661c7382f2dbeec  <= I2eb093d2a38ba8cf4be47d1d7f54ecc4 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I854a15bc7e9728b01c9a1960f6248dc9 != I82e0e091fba6f79cef97eacac4b43ecb[11] ) begin
                    Iefdcb71f2903b11f5cb0b8857f7a1727  <=  ~I8f9affdc5cda0fecc35dd15fc5aeb244 + 1;
                end else begin
                    Iefdcb71f2903b11f5cb0b8857f7a1727  <= I8f9affdc5cda0fecc35dd15fc5aeb244 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I854a15bc7e9728b01c9a1960f6248dc9 != Iea7da1f43ba202d753b0edb0be8b3fcf[13] ) begin
                    Ic57eb4a034247a4c952d8224ea9f2bac  <=  ~I615a443d49d1479338d033d2a2cab51f + 1;
                end else begin
                    Ic57eb4a034247a4c952d8224ea9f2bac  <= I615a443d49d1479338d033d2a2cab51f ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I854a15bc7e9728b01c9a1960f6248dc9 != Iba9f33c08db89a7f120cc1e3eaf05dec[0] ) begin
                    Iad4ea0196eb32f9a152c9e6fe5059e46  <=  ~I0635a3270a9653ca0f23c116fd5b2f97 + 1;
                end else begin
                    Iad4ea0196eb32f9a152c9e6fe5059e46  <= I0635a3270a9653ca0f23c116fd5b2f97 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iae332cfd000fd0529684ab787041b5dc != Ib58043c04b5c4c86c1c67e57cc66dcf7[20] ) begin
                    Iadbd245bf842aebb456417579a3e6296  <=  ~I93a7c75ebce8fbf4c613b4d11dc98b72 + 1;
                end else begin
                    Iadbd245bf842aebb456417579a3e6296  <= I93a7c75ebce8fbf4c613b4d11dc98b72 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iae332cfd000fd0529684ab787041b5dc != Ie1cd04c7668d3f450c387a6c1ad778c7[8] ) begin
                    I9c15a6a5c0db11ede80ff6d04c9a56d8  <=  ~I39334aa9d55bcc001ece37ce2a6c329c + 1;
                end else begin
                    I9c15a6a5c0db11ede80ff6d04c9a56d8  <= I39334aa9d55bcc001ece37ce2a6c329c ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iae332cfd000fd0529684ab787041b5dc != I8e591d83170c8ba46d31c61935311b22[11] ) begin
                    Ie95f1a7e0effcec0aa423dc803056a13  <=  ~I07e328d23da9383a296ecb03679ec74b + 1;
                end else begin
                    Ie95f1a7e0effcec0aa423dc803056a13  <= I07e328d23da9383a296ecb03679ec74b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iae332cfd000fd0529684ab787041b5dc != Ibde51eb91b3ca50a8a0513c94bd7be15[0] ) begin
                    Ia8ff29ed728e7f2ae4213f00328b495d  <=  ~I8a6e1eace6152af5c98c415804cb60fa + 1;
                end else begin
                    Ia8ff29ed728e7f2ae4213f00328b495d  <= I8a6e1eace6152af5c98c415804cb60fa ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I70148fe95244eebf7f0ec953703398de != Ibc0871b3c992fd278815fdbefcd2bac0[20] ) begin
                    I7103aa739616a39c03e675ea0efb0335  <=  ~I6ed4d6c350e8691b3a12ab51419cfa65 + 1;
                end else begin
                    I7103aa739616a39c03e675ea0efb0335  <= I6ed4d6c350e8691b3a12ab51419cfa65 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I70148fe95244eebf7f0ec953703398de != If511a6ea6aa5cda5353658d8e192791f[8] ) begin
                    I5827bc87b5db1801b7db16e1e61515db  <=  ~Ie2b9ed680dac51ac866cb830ca17ef84 + 1;
                end else begin
                    I5827bc87b5db1801b7db16e1e61515db  <= Ie2b9ed680dac51ac866cb830ca17ef84 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I70148fe95244eebf7f0ec953703398de != I02b62fafd371de339f299f8aefec6c43[11] ) begin
                    I5b4305bef5b4350c1d7ae143667afddd  <=  ~Ie439b520bbb0c8b29a5ecea167acb1c9 + 1;
                end else begin
                    I5b4305bef5b4350c1d7ae143667afddd  <= Ie439b520bbb0c8b29a5ecea167acb1c9 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I70148fe95244eebf7f0ec953703398de != Ifb94196d1653a0166567e170f06ec0db[0] ) begin
                    I70717726200ec02929f679ef05496455  <=  ~I9f8ef3295578acf5b0a42d074a15a70b + 1;
                end else begin
                    I70717726200ec02929f679ef05496455  <= I9f8ef3295578acf5b0a42d074a15a70b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I24ee2d953e65fefdc73b3d3c4c0ddd05 != I8695e1e94cbfcbe4b9eae315b042529e[20] ) begin
                    I16e3559c63ebfed83d6698fc9a9cd93a  <=  ~Ief01b06341d489e36ee344fd52084ccf + 1;
                end else begin
                    I16e3559c63ebfed83d6698fc9a9cd93a  <= Ief01b06341d489e36ee344fd52084ccf ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I24ee2d953e65fefdc73b3d3c4c0ddd05 != Ib0bf69cc797f330fb2546eb46d2d6f76[8] ) begin
                    Ie7f3f1d6cee7f02ae1b17740ed54c049  <=  ~I3b72a085b104e17dca3d8b2824f84e97 + 1;
                end else begin
                    Ie7f3f1d6cee7f02ae1b17740ed54c049  <= I3b72a085b104e17dca3d8b2824f84e97 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I24ee2d953e65fefdc73b3d3c4c0ddd05 != I0e0b15868b02ca52b260f17f150d237e[11] ) begin
                    If5dfdadb3868ed5a495007362f7db648  <=  ~I5e1f41e23887493db1d723e1e2cbd996 + 1;
                end else begin
                    If5dfdadb3868ed5a495007362f7db648  <= I5e1f41e23887493db1d723e1e2cbd996 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I24ee2d953e65fefdc73b3d3c4c0ddd05 != I9cf7557e2cac4532a77fcb212712db0f[0] ) begin
                    Iaf1e4c7dae6ad89567836877c08f57d2  <=  ~I0e6f4c7bdc39bd22833f3d9fcfa55f1d + 1;
                end else begin
                    Iaf1e4c7dae6ad89567836877c08f57d2  <= I0e6f4c7bdc39bd22833f3d9fcfa55f1d ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie3a5f8eec283fd4f682b5d0f909b051c != Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[20] ) begin
                    I88c10c47ae424fbdcb852fbf1e94127c  <=  ~Ie346802a8898b4b075be289e062b462c + 1;
                end else begin
                    I88c10c47ae424fbdcb852fbf1e94127c  <= Ie346802a8898b4b075be289e062b462c ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie3a5f8eec283fd4f682b5d0f909b051c != Iec7404bc79c58d4d2538fcdf659e9134[8] ) begin
                    I06c7728ef64be8311f48d10d766d0c44  <=  ~I82ea6f21706a97166ef11af548e80392 + 1;
                end else begin
                    I06c7728ef64be8311f48d10d766d0c44  <= I82ea6f21706a97166ef11af548e80392 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie3a5f8eec283fd4f682b5d0f909b051c != I3c0b6f53f0a5cda5b6758b2ee2c83b92[11] ) begin
                    I02cbb4255db2b21ea32140f9e9ddb36b  <=  ~I5f38764f6ecc2dcd1fdd5316102f1f82 + 1;
                end else begin
                    I02cbb4255db2b21ea32140f9e9ddb36b  <= I5f38764f6ecc2dcd1fdd5316102f1f82 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie3a5f8eec283fd4f682b5d0f909b051c != I3159d7faeee1a904c409bde1967d2c21[0] ) begin
                    Icd09aa81e9b43528af73e23b2f0f80cb  <=  ~Id4034bf7a0e92a6c92d0187e00d3df99 + 1;
                end else begin
                    Icd09aa81e9b43528af73e23b2f0f80cb  <= Id4034bf7a0e92a6c92d0187e00d3df99 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I781d986d7fd6c2fec3a8cf3f29545174 != I651d700a00d7004d8728bc7356f30926[7] ) begin
                    I6ff7b86cd7f63f9243646f1be10b2577  <=  ~I44692fd63388c57268ea9035a7e4c3ef + 1;
                end else begin
                    I6ff7b86cd7f63f9243646f1be10b2577  <= I44692fd63388c57268ea9035a7e4c3ef ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I781d986d7fd6c2fec3a8cf3f29545174 != Ia8a468877c9f96713c8141df9205f92a[10] ) begin
                    Ie631e40caade823a196370fc3358f042  <=  ~I0c2892a34e5236f1366959eadfd83825 + 1;
                end else begin
                    Ie631e40caade823a196370fc3358f042  <= I0c2892a34e5236f1366959eadfd83825 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I781d986d7fd6c2fec3a8cf3f29545174 != I35dfb5ece5e04504d6e74739ae99c9cc[0] ) begin
                    I6ebb2b94f0f80425f8401ae823d92a1d  <=  ~Iccef2754044e7066e191bc5e1a3805f1 + 1;
                end else begin
                    I6ebb2b94f0f80425f8401ae823d92a1d  <= Iccef2754044e7066e191bc5e1a3805f1 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib4db8131350f8605e00907234aff901d != Ic2580cbeec8c11a19bd1e2ebc29d255e[7] ) begin
                    I8c35c5b343b552c22000e194c517ca12  <=  ~I8ace46f1c56cfb3f4773324e0f8cae58 + 1;
                end else begin
                    I8c35c5b343b552c22000e194c517ca12  <= I8ace46f1c56cfb3f4773324e0f8cae58 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib4db8131350f8605e00907234aff901d != I4267622319ca65909a3b40484dc74d3a[10] ) begin
                    I37dca40506d61bdeab1255ed4892ca20  <=  ~I94ec0139bd827ef5dce2c5ee9eb9aded + 1;
                end else begin
                    I37dca40506d61bdeab1255ed4892ca20  <= I94ec0139bd827ef5dce2c5ee9eb9aded ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib4db8131350f8605e00907234aff901d != Iabff939ae4acf7d7b038e028c29b6166[0] ) begin
                    I4a2c3204a6a9936d4a215b46c0ffd045  <=  ~Ied62b116607c549ff5918d5b95e2118f + 1;
                end else begin
                    I4a2c3204a6a9936d4a215b46c0ffd045  <= Ied62b116607c549ff5918d5b95e2118f ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie093f0750b60d3aed75705637933f34c != If79ed5ee2b8710da0608c1e245d07d55[7] ) begin
                    Iee367c535d9c39f872d2ec043e7e7b33  <=  ~I9efa5796297bc922bc5fe17f8319a515 + 1;
                end else begin
                    Iee367c535d9c39f872d2ec043e7e7b33  <= I9efa5796297bc922bc5fe17f8319a515 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie093f0750b60d3aed75705637933f34c != Iedd7d4ea8d082b40244c04946dfb14a0[10] ) begin
                    I67347c413b5efd8ff9e0d5bc7ab2a047  <=  ~Ifa6908d8fda29713d7c1bbaa69b72b53 + 1;
                end else begin
                    I67347c413b5efd8ff9e0d5bc7ab2a047  <= Ifa6908d8fda29713d7c1bbaa69b72b53 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ie093f0750b60d3aed75705637933f34c != Ia14159444578c6dc88f2d5ea0317774b[0] ) begin
                    Ib02c0694762c4815448b2c8d3df767c2  <=  ~Ieb46857229186ce0391cddb2d30f434e + 1;
                end else begin
                    Ib02c0694762c4815448b2c8d3df767c2  <= Ieb46857229186ce0391cddb2d30f434e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Id2fba7c1b3dc7a75a5e0d90494d56962 != I9497bbb4f746969a95cff948a3ee9ade[7] ) begin
                    Ie76b0739aec66f8860870e66e87a6445  <=  ~I67fa03f808026b38ca5b4e71e21588bf + 1;
                end else begin
                    Ie76b0739aec66f8860870e66e87a6445  <= I67fa03f808026b38ca5b4e71e21588bf ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Id2fba7c1b3dc7a75a5e0d90494d56962 != I56e1fe0c7a62589c123876f2b4e57a26[10] ) begin
                    I613d4b1e3b9e812b785c9cf14fefdfe6  <=  ~I70938dfe09b0da9d87dafed6af3fa05c + 1;
                end else begin
                    I613d4b1e3b9e812b785c9cf14fefdfe6  <= I70938dfe09b0da9d87dafed6af3fa05c ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Id2fba7c1b3dc7a75a5e0d90494d56962 != Ie2306a5c441d621388b73195027fc118[0] ) begin
                    I98cee6efbbe565d3a4de16703189782f  <=  ~Iff30a4e14b6282e9ef92e7f58230b516 + 1;
                end else begin
                    I98cee6efbbe565d3a4de16703189782f  <= Iff30a4e14b6282e9ef92e7f58230b516 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9ecee74c445711a376133636ef414666 != I5b7caaeb34c43e66e8d095a859e708fe[21] ) begin
                    I4a777f0dd62b19dd340ad31517c4e789  <=  ~I43e0faf8070869ab0528a7a4a5cdc103 + 1;
                end else begin
                    I4a777f0dd62b19dd340ad31517c4e789  <= I43e0faf8070869ab0528a7a4a5cdc103 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9ecee74c445711a376133636ef414666 != I50976b0051e84b6a42fc1dbabd7d20ae[12] ) begin
                    I1e50c90010a3df1a8ce1cff811cc7a0c  <=  ~Ib2f0333fac7701ae4a5589d54005b8f3 + 1;
                end else begin
                    I1e50c90010a3df1a8ce1cff811cc7a0c  <= Ib2f0333fac7701ae4a5589d54005b8f3 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9ecee74c445711a376133636ef414666 != Iea7da1f43ba202d753b0edb0be8b3fcf[14] ) begin
                    Ia642db613c0ec1ca4e69afde7a14a839  <=  ~Ie4e1491da700923e81b2c1a246e528b1 + 1;
                end else begin
                    Ia642db613c0ec1ca4e69afde7a14a839  <= Ie4e1491da700923e81b2c1a246e528b1 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9ecee74c445711a376133636ef414666 != I700a0fbf81e57d4970ce07090ec4f2e2[0] ) begin
                    Ibf981c01a9d44cbea3c6d8ead92bc2ab  <=  ~Ie8602467de2ece2013878a6b8d3129a1 + 1;
                end else begin
                    Ibf981c01a9d44cbea3c6d8ead92bc2ab  <= Ie8602467de2ece2013878a6b8d3129a1 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ifb3cf6b88835d27220df837682c4dc93 != I61f0c04673dfb262ef6912eb2df39120[21] ) begin
                    Ib6ea4a822da2ea32e0abf6cf8a33d295  <=  ~I85c93c62f79b1703cb6928f96737cf27 + 1;
                end else begin
                    Ib6ea4a822da2ea32e0abf6cf8a33d295  <= I85c93c62f79b1703cb6928f96737cf27 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ifb3cf6b88835d27220df837682c4dc93 != I82e0e091fba6f79cef97eacac4b43ecb[12] ) begin
                    I2eb90278aaa54b9c8212b3b4af7c3617  <=  ~I3dc816ee6c2a818b32f6d4e1228704bf + 1;
                end else begin
                    I2eb90278aaa54b9c8212b3b4af7c3617  <= I3dc816ee6c2a818b32f6d4e1228704bf ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ifb3cf6b88835d27220df837682c4dc93 != I872f61d20baf011e867b44dc5539fc37[14] ) begin
                    I45bc13ae0e0554a79c62cd9c6aa8f2a5  <=  ~Id34d83701e815c01359bc5cd1b9c993c + 1;
                end else begin
                    I45bc13ae0e0554a79c62cd9c6aa8f2a5  <= Id34d83701e815c01359bc5cd1b9c993c ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ifb3cf6b88835d27220df837682c4dc93 != I6007914b3fb3011c3ab2f9a9d7794ab2[0] ) begin
                    I864c33e8ea204d20a9baef4584f22d4e  <=  ~I0a20e3e26261ba558d681346649cf0b3 + 1;
                end else begin
                    I864c33e8ea204d20a9baef4584f22d4e  <= I0a20e3e26261ba558d681346649cf0b3 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I386fbb3bd550891d682e137044e8773a != Ibeb5edab51cd6aedad9c2ecedaded6f5[21] ) begin
                    I9905e2686b350e8a6e7f790563a91294  <=  ~I331c6e8dbe2ea1e2232f82766926d0e6 + 1;
                end else begin
                    I9905e2686b350e8a6e7f790563a91294  <= I331c6e8dbe2ea1e2232f82766926d0e6 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I386fbb3bd550891d682e137044e8773a != I04302edb2671c5bc0ca2673cd53935e1[12] ) begin
                    Icc93450a007cee4c0a42717ed7600528  <=  ~Ie27046fd2751357e4a81dc62086f00be + 1;
                end else begin
                    Icc93450a007cee4c0a42717ed7600528  <= Ie27046fd2751357e4a81dc62086f00be ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I386fbb3bd550891d682e137044e8773a != I6f5c991e5fdcf56d582c6f80eb6731df[14] ) begin
                    Ic4a6c02880a9aead7353332708e3f388  <=  ~I0897ceba8201bc14a49ab30318183875 + 1;
                end else begin
                    Ic4a6c02880a9aead7353332708e3f388  <= I0897ceba8201bc14a49ab30318183875 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I386fbb3bd550891d682e137044e8773a != I2096f40fe62e9d6f1ff96f258ffdbe33[0] ) begin
                    I6ad3228e0e2e1f19648d73e83ba5a229  <=  ~Ie7b15aa8ce2492bfb433894efeb967f3 + 1;
                end else begin
                    I6ad3228e0e2e1f19648d73e83ba5a229  <= Ie7b15aa8ce2492bfb433894efeb967f3 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I7ede7d2e1c2730b3b71340b11e880f5b != Iceb64ab2ff8a2e0dfdb74803811d4cfe[21] ) begin
                    I995d2809ffaf0ecda6a004d01cb9c8c4  <=  ~I255add08e982f701508a98db221e617d + 1;
                end else begin
                    I995d2809ffaf0ecda6a004d01cb9c8c4  <= I255add08e982f701508a98db221e617d ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I7ede7d2e1c2730b3b71340b11e880f5b != I480a0f6d6c3eb936de10a72749f6cd3f[12] ) begin
                    Idefa29d4d4e2a6e9147f84893520096f  <=  ~If7ca4919fa1449f38777f742ee1fb875 + 1;
                end else begin
                    Idefa29d4d4e2a6e9147f84893520096f  <= If7ca4919fa1449f38777f742ee1fb875 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I7ede7d2e1c2730b3b71340b11e880f5b != Ia5cc3055ba3365e64cf59c4d4fd3f093[14] ) begin
                    Ic044d7419cc43736d278c2df33b4a3cc  <=  ~I24cafcb5b9825321c54e84827a662fdc + 1;
                end else begin
                    Ic044d7419cc43736d278c2df33b4a3cc  <= I24cafcb5b9825321c54e84827a662fdc ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I7ede7d2e1c2730b3b71340b11e880f5b != I93d8b7a24702bacbfc528242991516a9[0] ) begin
                    Ie099210a99a4899c53baf39559592690  <=  ~I3ede71cb7cb39774aedb9889240a2462 + 1;
                end else begin
                    Ie099210a99a4899c53baf39559592690  <= I3ede71cb7cb39774aedb9889240a2462 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I64c65fad4a7d958d625c783626808175 != Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[21] ) begin
                    Icd2e75e47cab1d539ba9ff1b6e1d7155  <=  ~I24da9598a6840d3ba7b12fe4f638219b + 1;
                end else begin
                    Icd2e75e47cab1d539ba9ff1b6e1d7155  <= I24da9598a6840d3ba7b12fe4f638219b ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I64c65fad4a7d958d625c783626808175 != I0e0b15868b02ca52b260f17f150d237e[12] ) begin
                    Ia1ee5579358b564de06c08ca418a9bf4  <=  ~I0358ca8833007cec4ce5047db32ab7a3 + 1;
                end else begin
                    Ia1ee5579358b564de06c08ca418a9bf4  <= I0358ca8833007cec4ce5047db32ab7a3 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I64c65fad4a7d958d625c783626808175 != Id6f07dee3e47f39e3b43329c26f690f7[8] ) begin
                    Id3e0c98bff2636e216b4d3a0ffd51054  <=  ~I85b5354463c1c15f91ed67292da912c1 + 1;
                end else begin
                    Id3e0c98bff2636e216b4d3a0ffd51054  <= I85b5354463c1c15f91ed67292da912c1 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I64c65fad4a7d958d625c783626808175 != If0863fae91b2ec980ebdb26cfc90ae2e[0] ) begin
                    Ieeec71d9df4613555fade2ced7b3baf1  <=  ~Ie93731739ace44811198d0fd95b04a6a + 1;
                end else begin
                    Ieeec71d9df4613555fade2ced7b3baf1  <= Ie93731739ace44811198d0fd95b04a6a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib2e0cd0a2b51c3a265bdd20834c0ed2d != Ib58043c04b5c4c86c1c67e57cc66dcf7[21] ) begin
                    Ifc8ece44a4e68c3117eda9e65f3084d2  <=  ~I464926faf4e005ad491b0bf93a365e07 + 1;
                end else begin
                    Ifc8ece44a4e68c3117eda9e65f3084d2  <= I464926faf4e005ad491b0bf93a365e07 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib2e0cd0a2b51c3a265bdd20834c0ed2d != I3c0b6f53f0a5cda5b6758b2ee2c83b92[12] ) begin
                    I65354f2069de0c25bbe7cd50fbe892aa  <=  ~Icdaaccfead6f2d5ac2ce19caf1104d57 + 1;
                end else begin
                    I65354f2069de0c25bbe7cd50fbe892aa  <= Icdaaccfead6f2d5ac2ce19caf1104d57 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib2e0cd0a2b51c3a265bdd20834c0ed2d != Ic7f04c065f8ff82c2288f1de77d37189[8] ) begin
                    Ife1164cad7cda4aa9a08d94dfe86add6  <=  ~I916d6f9429f2b0cc1bd6fb900484cde5 + 1;
                end else begin
                    Ife1164cad7cda4aa9a08d94dfe86add6  <= I916d6f9429f2b0cc1bd6fb900484cde5 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ib2e0cd0a2b51c3a265bdd20834c0ed2d != I9ec29a319384efd562c2337e1857cb4e[0] ) begin
                    I4931884e3544af182bcda9061091a42d  <=  ~I0142f9b3d361a0d88522f1c5f54aca84 + 1;
                end else begin
                    I4931884e3544af182bcda9061091a42d  <= I0142f9b3d361a0d88522f1c5f54aca84 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I67be0b66c8d0680eb23290a4b3885af3 != Ibc0871b3c992fd278815fdbefcd2bac0[21] ) begin
                    I0296d01fd3f9a269a617efd4beea9b8b  <=  ~Ie6871983b4f81b5321519647e628bd0e + 1;
                end else begin
                    I0296d01fd3f9a269a617efd4beea9b8b  <= Ie6871983b4f81b5321519647e628bd0e ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I67be0b66c8d0680eb23290a4b3885af3 != I8e591d83170c8ba46d31c61935311b22[12] ) begin
                    I106deaff50b8480eac31ddbae2ec7c61  <=  ~I17d7be125df22153fc1ed051d4e0770a + 1;
                end else begin
                    I106deaff50b8480eac31ddbae2ec7c61  <= I17d7be125df22153fc1ed051d4e0770a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I67be0b66c8d0680eb23290a4b3885af3 != Ieb244944e7ee8236a207924f56fbc689[8] ) begin
                    I5669856f88f5e2c98f64df696db76414  <=  ~I50b13959e06243e54fad2088eaf65aa7 + 1;
                end else begin
                    I5669856f88f5e2c98f64df696db76414  <= I50b13959e06243e54fad2088eaf65aa7 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I67be0b66c8d0680eb23290a4b3885af3 != Ia56ecc024eae608d7de1509d75139dc2[0] ) begin
                    Ib3fb10da528d450251764a9b9ede0dba  <=  ~I7a423d609b492f73d5a322849b4b1cce + 1;
                end else begin
                    Ib3fb10da528d450251764a9b9ede0dba  <= I7a423d609b492f73d5a322849b4b1cce ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I01148401f7d058614dc1ae6ed3c8bd94 != I8695e1e94cbfcbe4b9eae315b042529e[21] ) begin
                    I9747a02384abb1c2dd1f52b3a5a999cc  <=  ~Iefec67e214d1868670a34a7297d4a1c8 + 1;
                end else begin
                    I9747a02384abb1c2dd1f52b3a5a999cc  <= Iefec67e214d1868670a34a7297d4a1c8 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I01148401f7d058614dc1ae6ed3c8bd94 != I02b62fafd371de339f299f8aefec6c43[12] ) begin
                    I2795d21d343b83a69146314a2407cfa2  <=  ~Iae7da7fdc002b635ce4285d6916d8156 + 1;
                end else begin
                    I2795d21d343b83a69146314a2407cfa2  <= Iae7da7fdc002b635ce4285d6916d8156 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I01148401f7d058614dc1ae6ed3c8bd94 != Ie9b2be4c32334220e134e041ca8dfc06[8] ) begin
                    I1b7a401bc11741e6f011fb9895b5c797  <=  ~Ic561e44b2caeae84df6720f1afa3e8f6 + 1;
                end else begin
                    I1b7a401bc11741e6f011fb9895b5c797  <= Ic561e44b2caeae84df6720f1afa3e8f6 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I01148401f7d058614dc1ae6ed3c8bd94 != Iebcd65ea41cd38bfe3c8577277809acd[0] ) begin
                    Icdc9e676957b2223d60c413331fa982f  <=  ~I5be062f5b52e104ca67e615ce75a7c80 + 1;
                end else begin
                    Icdc9e676957b2223d60c413331fa982f  <= I5be062f5b52e104ca67e615ce75a7c80 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I3394319c370daf6102be00d938d55769 != Ib0bf69cc797f330fb2546eb46d2d6f76[9] ) begin
                    Ib196f5bcf9152703dc32c5101076600a  <=  ~Iecdde23e34c34ee0055be41f44959a19 + 1;
                end else begin
                    Ib196f5bcf9152703dc32c5101076600a  <= Iecdde23e34c34ee0055be41f44959a19 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I3394319c370daf6102be00d938d55769 != I651d700a00d7004d8728bc7356f30926[8] ) begin
                    I165653ab165cfafe2b74cd441331f9e1  <=  ~Ibe09be9cad0e56d5403868d072d7d628 + 1;
                end else begin
                    I165653ab165cfafe2b74cd441331f9e1  <= Ibe09be9cad0e56d5403868d072d7d628 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I3394319c370daf6102be00d938d55769 != I4267622319ca65909a3b40484dc74d3a[11] ) begin
                    I340c98b886123c541a1b8d9fc8a6d48c  <=  ~I464e1f3c13acaf466afb354a9b35ba0a + 1;
                end else begin
                    I340c98b886123c541a1b8d9fc8a6d48c  <= I464e1f3c13acaf466afb354a9b35ba0a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I3394319c370daf6102be00d938d55769 != I75be12b14694ebcb5aff6e5d3e576315[0] ) begin
                    I381f6051282c062ccf53866830344cd4  <=  ~I160a465c22073a53510e8a4c489c3321 + 1;
                end else begin
                    I381f6051282c062ccf53866830344cd4  <= I160a465c22073a53510e8a4c489c3321 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I24d6a334dd15ccdea558f32cd029e6d1 != Iec7404bc79c58d4d2538fcdf659e9134[9] ) begin
                    I9fe11f6c8147391aa4a5afd1a4e4f731  <=  ~I9e86d3e49827861b24f4fbeb308ad3a4 + 1;
                end else begin
                    I9fe11f6c8147391aa4a5afd1a4e4f731  <= I9e86d3e49827861b24f4fbeb308ad3a4 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I24d6a334dd15ccdea558f32cd029e6d1 != Ic2580cbeec8c11a19bd1e2ebc29d255e[8] ) begin
                    Ibf80bb564263ea85bd886a8617f09bb2  <=  ~Ib96b7d796e20967e89a47e01bf424e59 + 1;
                end else begin
                    Ibf80bb564263ea85bd886a8617f09bb2  <= Ib96b7d796e20967e89a47e01bf424e59 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I24d6a334dd15ccdea558f32cd029e6d1 != Iedd7d4ea8d082b40244c04946dfb14a0[11] ) begin
                    I72b1bb104bf2843f161448baf7aab44b  <=  ~I565e666f6ba14b4c25e0dd402a3266e1 + 1;
                end else begin
                    I72b1bb104bf2843f161448baf7aab44b  <= I565e666f6ba14b4c25e0dd402a3266e1 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I24d6a334dd15ccdea558f32cd029e6d1 != I8e06fe414cd04103baf3882771a63e2c[0] ) begin
                    Icfc21935c007fbbceb2a67ebe1a68a0b  <=  ~I97e8bac5becd5128bc70f3bb48f73e6c + 1;
                end else begin
                    Icfc21935c007fbbceb2a67ebe1a68a0b  <= I97e8bac5becd5128bc70f3bb48f73e6c ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I3a41f68bca2d7edd1f5738c4fda8e73c != Ie1cd04c7668d3f450c387a6c1ad778c7[9] ) begin
                    I8922487573e02d684a3d71448c3828f5  <=  ~Iced39475c6e5e3d8f36d2a5c5a80f146 + 1;
                end else begin
                    I8922487573e02d684a3d71448c3828f5  <= Iced39475c6e5e3d8f36d2a5c5a80f146 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I3a41f68bca2d7edd1f5738c4fda8e73c != If79ed5ee2b8710da0608c1e245d07d55[8] ) begin
                    I68bb1f26f878862f288c1f57049cf58b  <=  ~Idcbd423c2b963c1f693dea2ddf428195 + 1;
                end else begin
                    I68bb1f26f878862f288c1f57049cf58b  <= Idcbd423c2b963c1f693dea2ddf428195 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I3a41f68bca2d7edd1f5738c4fda8e73c != I56e1fe0c7a62589c123876f2b4e57a26[11] ) begin
                    I848ed394bd4f0b199d11c0ff458394a7  <=  ~If1640e294bdcc51ee12fca5b3a33be6d + 1;
                end else begin
                    I848ed394bd4f0b199d11c0ff458394a7  <= If1640e294bdcc51ee12fca5b3a33be6d ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I3a41f68bca2d7edd1f5738c4fda8e73c != I0fe8574049166c363c7cc816b1435009[0] ) begin
                    I120d597a80158374726e064fb0f099fb  <=  ~I4754c6c355e632d2ed1336b5a88c3b46 + 1;
                end else begin
                    I120d597a80158374726e064fb0f099fb  <= I4754c6c355e632d2ed1336b5a88c3b46 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9ef1784d165492f3482d14f475732451 != If511a6ea6aa5cda5353658d8e192791f[9] ) begin
                    I1c85c8f73ef80a6808c6aec0c8eca8ab  <=  ~I1634d703ad5d6e58a97b13ef957bdbec + 1;
                end else begin
                    I1c85c8f73ef80a6808c6aec0c8eca8ab  <= I1634d703ad5d6e58a97b13ef957bdbec ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9ef1784d165492f3482d14f475732451 != I9497bbb4f746969a95cff948a3ee9ade[8] ) begin
                    I50383e3d7c172eedfa00aa50a9faac4c  <=  ~I804e1e6a01edeb780b0159ecae707b71 + 1;
                end else begin
                    I50383e3d7c172eedfa00aa50a9faac4c  <= I804e1e6a01edeb780b0159ecae707b71 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9ef1784d165492f3482d14f475732451 != Ia8a468877c9f96713c8141df9205f92a[11] ) begin
                    I4c971e714427664c59c6371e14781bae  <=  ~Iea3c0f3c3c3017fe87a3b01647189fe0 + 1;
                end else begin
                    I4c971e714427664c59c6371e14781bae  <= Iea3c0f3c3c3017fe87a3b01647189fe0 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9ef1784d165492f3482d14f475732451 != Id5f435c07240d5fe4a0e48c8f25ad0b7[0] ) begin
                    I2520aa556aadf851f58f0b1820498730  <=  ~I756b7d7e6bd3e71afa472e7e4727264a + 1;
                end else begin
                    I2520aa556aadf851f58f0b1820498730  <= I756b7d7e6bd3e71afa472e7e4727264a ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9d9378337a77515a4e8d04fb88938808 != Ibeb5edab51cd6aedad9c2ecedaded6f5[22] ) begin
                    I524e78ae6a4204e17ba4532dba047d4b  <=  ~Ifbeae0a2acf80eda6ffd050d3bb07eb3 + 1;
                end else begin
                    I524e78ae6a4204e17ba4532dba047d4b  <= Ifbeae0a2acf80eda6ffd050d3bb07eb3 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9d9378337a77515a4e8d04fb88938808 != I480a0f6d6c3eb936de10a72749f6cd3f[13] ) begin
                    Id1fbbe0594dae272856566522633bb3d  <=  ~I990ab4dcb70ee860c2c40f306ef314d3 + 1;
                end else begin
                    Id1fbbe0594dae272856566522633bb3d  <= I990ab4dcb70ee860c2c40f306ef314d3 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9d9378337a77515a4e8d04fb88938808 != Iea7da1f43ba202d753b0edb0be8b3fcf[15] ) begin
                    I432aa7cb844286c442356954f8814260  <=  ~Ib131087ea9ccc4bd161c3f9ac2c72303 + 1;
                end else begin
                    I432aa7cb844286c442356954f8814260  <= Ib131087ea9ccc4bd161c3f9ac2c72303 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (I9d9378337a77515a4e8d04fb88938808 != I1ae21e0db88f955c4f08f6d52f58974d[0] ) begin
                    I6203f49a08107f7185ebadeecf2c16b0  <=  ~I9a967ac9d11583faaa783984229aeb2c + 1;
                end else begin
                    I6203f49a08107f7185ebadeecf2c16b0  <= I9a967ac9d11583faaa783984229aeb2c ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (If0e20ef9aa69b77ae0e58ca3dfc9998f != Iceb64ab2ff8a2e0dfdb74803811d4cfe[22] ) begin
                    I4e8ebc46bc068c3f9889d970db131112  <=  ~Ib9921dfcf121e5f4ac4d8be83a868210 + 1;
                end else begin
                    I4e8ebc46bc068c3f9889d970db131112  <= Ib9921dfcf121e5f4ac4d8be83a868210 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (If0e20ef9aa69b77ae0e58ca3dfc9998f != I50976b0051e84b6a42fc1dbabd7d20ae[13] ) begin
                    Ie1817cbf3a80dae435a5571dfbd2f5ad  <=  ~If22d8fd45caed08b2c7cee8b7349700f + 1;
                end else begin
                    Ie1817cbf3a80dae435a5571dfbd2f5ad  <= If22d8fd45caed08b2c7cee8b7349700f ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (If0e20ef9aa69b77ae0e58ca3dfc9998f != I872f61d20baf011e867b44dc5539fc37[15] ) begin
                    I92678f5b52c9c55556ff7f17f0f607b7  <=  ~Iabf029e67c7f827faf17b6518cd1bfa3 + 1;
                end else begin
                    I92678f5b52c9c55556ff7f17f0f607b7  <= Iabf029e67c7f827faf17b6518cd1bfa3 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (If0e20ef9aa69b77ae0e58ca3dfc9998f != I92efddd59e1ea92902a295c0b8385c68[0] ) begin
                    Ia706fb593b63cebbee0321c154cb859b  <=  ~Iaeab83001c6285630e3404ae67227f46 + 1;
                end else begin
                    Ia706fb593b63cebbee0321c154cb859b  <= Iaeab83001c6285630e3404ae67227f46 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iec2cb48bb1b58f268bf164d5e8a8120f != I5b7caaeb34c43e66e8d095a859e708fe[22] ) begin
                    Ib75747cb32130d44b338ed8c8af8ca11  <=  ~I53ac6d02d2bfc9aca9469148753070a7 + 1;
                end else begin
                    Ib75747cb32130d44b338ed8c8af8ca11  <= I53ac6d02d2bfc9aca9469148753070a7 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iec2cb48bb1b58f268bf164d5e8a8120f != I82e0e091fba6f79cef97eacac4b43ecb[13] ) begin
                    I43493f70f0336453d77caf7f27503daa  <=  ~I61992979f60b26d313efd1dc23bb54ab + 1;
                end else begin
                    I43493f70f0336453d77caf7f27503daa  <= I61992979f60b26d313efd1dc23bb54ab ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iec2cb48bb1b58f268bf164d5e8a8120f != I6f5c991e5fdcf56d582c6f80eb6731df[15] ) begin
                    I7fb3b66cb48521f8715f66bf5642cdb2  <=  ~I8b46b3f0835310114208963de7ac8e97 + 1;
                end else begin
                    I7fb3b66cb48521f8715f66bf5642cdb2  <= I8b46b3f0835310114208963de7ac8e97 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Iec2cb48bb1b58f268bf164d5e8a8120f != I56948ad2b2cc245bb1003fd71ae5f899[0] ) begin
                    Ia4b5f2b07556629673fc6576bc49a5dc  <=  ~Icda26ba6f5c7f77a80776b2c1bbc975d + 1;
                end else begin
                    Ia4b5f2b07556629673fc6576bc49a5dc  <= Icda26ba6f5c7f77a80776b2c1bbc975d ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ia4ae7c98720d43a604f28dfc5dd67d50 != I61f0c04673dfb262ef6912eb2df39120[22] ) begin
                    Id1659ccdeaea3e59eb2d3f65a65ebd05  <=  ~I0863565b3ae88137a2384750436f9e19 + 1;
                end else begin
                    Id1659ccdeaea3e59eb2d3f65a65ebd05  <= I0863565b3ae88137a2384750436f9e19 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ia4ae7c98720d43a604f28dfc5dd67d50 != I04302edb2671c5bc0ca2673cd53935e1[13] ) begin
                    I9ec9f389d0489908d497487e44c6edcd  <=  ~Id646110f8d09cd47dc7695e05f73efc6 + 1;
                end else begin
                    I9ec9f389d0489908d497487e44c6edcd  <= Id646110f8d09cd47dc7695e05f73efc6 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ia4ae7c98720d43a604f28dfc5dd67d50 != Ia5cc3055ba3365e64cf59c4d4fd3f093[15] ) begin
                    I6714551e8885ef5e4490673fe1b2dad1  <=  ~I5999eef2304e579a3d47e4f15ba336e1 + 1;
                end else begin
                    I6714551e8885ef5e4490673fe1b2dad1  <= I5999eef2304e579a3d47e4f15ba336e1 ;
                end
             end
             if (Iac11baea9832d6493626d2fe40fd385f) begin
                if (Ia4ae7c98720d43a604f28dfc5dd67d50 != I5fb5081b7a2da89115c0080b0967974d[0] ) begin
                    Ic532c6b85b156f821e0742f47239a65c  <=  ~Idd302bdc6ff8368a6b73d53bbc8f8425 + 1;
                end else begin
                    Ic532c6b85b156f821e0742f47239a65c  <= Idd302bdc6ff8368a6b73d53bbc8f8425 ;
                end
             end
       end
   end


   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
            I748f85f6680918a2e992df339b4b6558                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I95878a848ec38c4f334bc1915576e6d6[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib58043c04b5c4c86c1c67e57cc66dcf7[0]  <= 1'b0;
            I95878a848ec38c4f334bc1915576e6d6[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib58043c04b5c4c86c1c67e57cc66dcf7[1]  <= 1'b0;
            I95878a848ec38c4f334bc1915576e6d6[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib58043c04b5c4c86c1c67e57cc66dcf7[2]  <= 1'b0;
            I95878a848ec38c4f334bc1915576e6d6[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib58043c04b5c4c86c1c67e57cc66dcf7[3]  <= 1'b0;
            I95878a848ec38c4f334bc1915576e6d6[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib58043c04b5c4c86c1c67e57cc66dcf7[4]  <= 1'b0;
            I95878a848ec38c4f334bc1915576e6d6[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib58043c04b5c4c86c1c67e57cc66dcf7[5]  <= 1'b0;
            I95878a848ec38c4f334bc1915576e6d6[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib58043c04b5c4c86c1c67e57cc66dcf7[6]  <= 1'b0;
            I95878a848ec38c4f334bc1915576e6d6[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib58043c04b5c4c86c1c67e57cc66dcf7[7]  <= 1'b0;
            I95878a848ec38c4f334bc1915576e6d6[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib58043c04b5c4c86c1c67e57cc66dcf7[8]  <= 1'b0;
            I95878a848ec38c4f334bc1915576e6d6[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib58043c04b5c4c86c1c67e57cc66dcf7[9]  <= 1'b0;
            I95878a848ec38c4f334bc1915576e6d6[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib58043c04b5c4c86c1c67e57cc66dcf7[10]  <= 1'b0;
            I95878a848ec38c4f334bc1915576e6d6[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib58043c04b5c4c86c1c67e57cc66dcf7[11]  <= 1'b0;
            I95878a848ec38c4f334bc1915576e6d6[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib58043c04b5c4c86c1c67e57cc66dcf7[12]  <= 1'b0;
            I95878a848ec38c4f334bc1915576e6d6[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib58043c04b5c4c86c1c67e57cc66dcf7[13]  <= 1'b0;
            I95878a848ec38c4f334bc1915576e6d6[14]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib58043c04b5c4c86c1c67e57cc66dcf7[14]  <= 1'b0;
            I95878a848ec38c4f334bc1915576e6d6[15]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib58043c04b5c4c86c1c67e57cc66dcf7[15]  <= 1'b0;
            I95878a848ec38c4f334bc1915576e6d6[16]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib58043c04b5c4c86c1c67e57cc66dcf7[16]  <= 1'b0;
            I95878a848ec38c4f334bc1915576e6d6[17]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib58043c04b5c4c86c1c67e57cc66dcf7[17]  <= 1'b0;
            I95878a848ec38c4f334bc1915576e6d6[18]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib58043c04b5c4c86c1c67e57cc66dcf7[18]  <= 1'b0;
            I95878a848ec38c4f334bc1915576e6d6[19]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib58043c04b5c4c86c1c67e57cc66dcf7[19]  <= 1'b0;
            I95878a848ec38c4f334bc1915576e6d6[20]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib58043c04b5c4c86c1c67e57cc66dcf7[20]  <= 1'b0;
            I95878a848ec38c4f334bc1915576e6d6[21]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib58043c04b5c4c86c1c67e57cc66dcf7[21]  <= 1'b0;
            Ib0f57837099e3fdf1b908d78bcda4a43                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I3eb1902edf9266038f39c281d134c26c[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibc0871b3c992fd278815fdbefcd2bac0[0]  <= 1'b0;
            I3eb1902edf9266038f39c281d134c26c[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibc0871b3c992fd278815fdbefcd2bac0[1]  <= 1'b0;
            I3eb1902edf9266038f39c281d134c26c[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibc0871b3c992fd278815fdbefcd2bac0[2]  <= 1'b0;
            I3eb1902edf9266038f39c281d134c26c[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibc0871b3c992fd278815fdbefcd2bac0[3]  <= 1'b0;
            I3eb1902edf9266038f39c281d134c26c[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibc0871b3c992fd278815fdbefcd2bac0[4]  <= 1'b0;
            I3eb1902edf9266038f39c281d134c26c[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibc0871b3c992fd278815fdbefcd2bac0[5]  <= 1'b0;
            I3eb1902edf9266038f39c281d134c26c[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibc0871b3c992fd278815fdbefcd2bac0[6]  <= 1'b0;
            I3eb1902edf9266038f39c281d134c26c[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibc0871b3c992fd278815fdbefcd2bac0[7]  <= 1'b0;
            I3eb1902edf9266038f39c281d134c26c[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibc0871b3c992fd278815fdbefcd2bac0[8]  <= 1'b0;
            I3eb1902edf9266038f39c281d134c26c[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibc0871b3c992fd278815fdbefcd2bac0[9]  <= 1'b0;
            I3eb1902edf9266038f39c281d134c26c[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibc0871b3c992fd278815fdbefcd2bac0[10]  <= 1'b0;
            I3eb1902edf9266038f39c281d134c26c[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibc0871b3c992fd278815fdbefcd2bac0[11]  <= 1'b0;
            I3eb1902edf9266038f39c281d134c26c[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibc0871b3c992fd278815fdbefcd2bac0[12]  <= 1'b0;
            I3eb1902edf9266038f39c281d134c26c[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibc0871b3c992fd278815fdbefcd2bac0[13]  <= 1'b0;
            I3eb1902edf9266038f39c281d134c26c[14]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibc0871b3c992fd278815fdbefcd2bac0[14]  <= 1'b0;
            I3eb1902edf9266038f39c281d134c26c[15]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibc0871b3c992fd278815fdbefcd2bac0[15]  <= 1'b0;
            I3eb1902edf9266038f39c281d134c26c[16]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibc0871b3c992fd278815fdbefcd2bac0[16]  <= 1'b0;
            I3eb1902edf9266038f39c281d134c26c[17]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibc0871b3c992fd278815fdbefcd2bac0[17]  <= 1'b0;
            I3eb1902edf9266038f39c281d134c26c[18]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibc0871b3c992fd278815fdbefcd2bac0[18]  <= 1'b0;
            I3eb1902edf9266038f39c281d134c26c[19]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibc0871b3c992fd278815fdbefcd2bac0[19]  <= 1'b0;
            I3eb1902edf9266038f39c281d134c26c[20]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibc0871b3c992fd278815fdbefcd2bac0[20]  <= 1'b0;
            I3eb1902edf9266038f39c281d134c26c[21]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibc0871b3c992fd278815fdbefcd2bac0[21]  <= 1'b0;
            If75e99660e3997f53f7b903bc366f47f                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ie791b43e8d5c9d1669743ea4d6e3139c[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8695e1e94cbfcbe4b9eae315b042529e[0]  <= 1'b0;
            Ie791b43e8d5c9d1669743ea4d6e3139c[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8695e1e94cbfcbe4b9eae315b042529e[1]  <= 1'b0;
            Ie791b43e8d5c9d1669743ea4d6e3139c[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8695e1e94cbfcbe4b9eae315b042529e[2]  <= 1'b0;
            Ie791b43e8d5c9d1669743ea4d6e3139c[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8695e1e94cbfcbe4b9eae315b042529e[3]  <= 1'b0;
            Ie791b43e8d5c9d1669743ea4d6e3139c[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8695e1e94cbfcbe4b9eae315b042529e[4]  <= 1'b0;
            Ie791b43e8d5c9d1669743ea4d6e3139c[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8695e1e94cbfcbe4b9eae315b042529e[5]  <= 1'b0;
            Ie791b43e8d5c9d1669743ea4d6e3139c[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8695e1e94cbfcbe4b9eae315b042529e[6]  <= 1'b0;
            Ie791b43e8d5c9d1669743ea4d6e3139c[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8695e1e94cbfcbe4b9eae315b042529e[7]  <= 1'b0;
            Ie791b43e8d5c9d1669743ea4d6e3139c[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8695e1e94cbfcbe4b9eae315b042529e[8]  <= 1'b0;
            Ie791b43e8d5c9d1669743ea4d6e3139c[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8695e1e94cbfcbe4b9eae315b042529e[9]  <= 1'b0;
            Ie791b43e8d5c9d1669743ea4d6e3139c[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8695e1e94cbfcbe4b9eae315b042529e[10]  <= 1'b0;
            Ie791b43e8d5c9d1669743ea4d6e3139c[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8695e1e94cbfcbe4b9eae315b042529e[11]  <= 1'b0;
            Ie791b43e8d5c9d1669743ea4d6e3139c[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8695e1e94cbfcbe4b9eae315b042529e[12]  <= 1'b0;
            Ie791b43e8d5c9d1669743ea4d6e3139c[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8695e1e94cbfcbe4b9eae315b042529e[13]  <= 1'b0;
            Ie791b43e8d5c9d1669743ea4d6e3139c[14]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8695e1e94cbfcbe4b9eae315b042529e[14]  <= 1'b0;
            Ie791b43e8d5c9d1669743ea4d6e3139c[15]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8695e1e94cbfcbe4b9eae315b042529e[15]  <= 1'b0;
            Ie791b43e8d5c9d1669743ea4d6e3139c[16]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8695e1e94cbfcbe4b9eae315b042529e[16]  <= 1'b0;
            Ie791b43e8d5c9d1669743ea4d6e3139c[17]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8695e1e94cbfcbe4b9eae315b042529e[17]  <= 1'b0;
            Ie791b43e8d5c9d1669743ea4d6e3139c[18]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8695e1e94cbfcbe4b9eae315b042529e[18]  <= 1'b0;
            Ie791b43e8d5c9d1669743ea4d6e3139c[19]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8695e1e94cbfcbe4b9eae315b042529e[19]  <= 1'b0;
            Ie791b43e8d5c9d1669743ea4d6e3139c[20]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8695e1e94cbfcbe4b9eae315b042529e[20]  <= 1'b0;
            Ie791b43e8d5c9d1669743ea4d6e3139c[21]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8695e1e94cbfcbe4b9eae315b042529e[21]  <= 1'b0;
            I3253481bee7dbfc0f3eac94c3252ee4e                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I5b892f00b2642ca102f7755ab512d067[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[0]  <= 1'b0;
            I5b892f00b2642ca102f7755ab512d067[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[1]  <= 1'b0;
            I5b892f00b2642ca102f7755ab512d067[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[2]  <= 1'b0;
            I5b892f00b2642ca102f7755ab512d067[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[3]  <= 1'b0;
            I5b892f00b2642ca102f7755ab512d067[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[4]  <= 1'b0;
            I5b892f00b2642ca102f7755ab512d067[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[5]  <= 1'b0;
            I5b892f00b2642ca102f7755ab512d067[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[6]  <= 1'b0;
            I5b892f00b2642ca102f7755ab512d067[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[7]  <= 1'b0;
            I5b892f00b2642ca102f7755ab512d067[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[8]  <= 1'b0;
            I5b892f00b2642ca102f7755ab512d067[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[9]  <= 1'b0;
            I5b892f00b2642ca102f7755ab512d067[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[10]  <= 1'b0;
            I5b892f00b2642ca102f7755ab512d067[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[11]  <= 1'b0;
            I5b892f00b2642ca102f7755ab512d067[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[12]  <= 1'b0;
            I5b892f00b2642ca102f7755ab512d067[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[13]  <= 1'b0;
            I5b892f00b2642ca102f7755ab512d067[14]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[14]  <= 1'b0;
            I5b892f00b2642ca102f7755ab512d067[15]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[15]  <= 1'b0;
            I5b892f00b2642ca102f7755ab512d067[16]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[16]  <= 1'b0;
            I5b892f00b2642ca102f7755ab512d067[17]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[17]  <= 1'b0;
            I5b892f00b2642ca102f7755ab512d067[18]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[18]  <= 1'b0;
            I5b892f00b2642ca102f7755ab512d067[19]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[19]  <= 1'b0;
            I5b892f00b2642ca102f7755ab512d067[20]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[20]  <= 1'b0;
            I5b892f00b2642ca102f7755ab512d067[21]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[21]  <= 1'b0;
            Ia80693da8182ee2c3708b6ec21d397d2                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I8f906015dba99b4a73dcf767cbd948ee[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I61f0c04673dfb262ef6912eb2df39120[0]  <= 1'b0;
            I8f906015dba99b4a73dcf767cbd948ee[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I61f0c04673dfb262ef6912eb2df39120[1]  <= 1'b0;
            I8f906015dba99b4a73dcf767cbd948ee[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I61f0c04673dfb262ef6912eb2df39120[2]  <= 1'b0;
            I8f906015dba99b4a73dcf767cbd948ee[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I61f0c04673dfb262ef6912eb2df39120[3]  <= 1'b0;
            I8f906015dba99b4a73dcf767cbd948ee[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I61f0c04673dfb262ef6912eb2df39120[4]  <= 1'b0;
            I8f906015dba99b4a73dcf767cbd948ee[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I61f0c04673dfb262ef6912eb2df39120[5]  <= 1'b0;
            I8f906015dba99b4a73dcf767cbd948ee[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I61f0c04673dfb262ef6912eb2df39120[6]  <= 1'b0;
            I8f906015dba99b4a73dcf767cbd948ee[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I61f0c04673dfb262ef6912eb2df39120[7]  <= 1'b0;
            I8f906015dba99b4a73dcf767cbd948ee[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I61f0c04673dfb262ef6912eb2df39120[8]  <= 1'b0;
            I8f906015dba99b4a73dcf767cbd948ee[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I61f0c04673dfb262ef6912eb2df39120[9]  <= 1'b0;
            I8f906015dba99b4a73dcf767cbd948ee[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I61f0c04673dfb262ef6912eb2df39120[10]  <= 1'b0;
            I8f906015dba99b4a73dcf767cbd948ee[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I61f0c04673dfb262ef6912eb2df39120[11]  <= 1'b0;
            I8f906015dba99b4a73dcf767cbd948ee[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I61f0c04673dfb262ef6912eb2df39120[12]  <= 1'b0;
            I8f906015dba99b4a73dcf767cbd948ee[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I61f0c04673dfb262ef6912eb2df39120[13]  <= 1'b0;
            I8f906015dba99b4a73dcf767cbd948ee[14]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I61f0c04673dfb262ef6912eb2df39120[14]  <= 1'b0;
            I8f906015dba99b4a73dcf767cbd948ee[15]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I61f0c04673dfb262ef6912eb2df39120[15]  <= 1'b0;
            I8f906015dba99b4a73dcf767cbd948ee[16]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I61f0c04673dfb262ef6912eb2df39120[16]  <= 1'b0;
            I8f906015dba99b4a73dcf767cbd948ee[17]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I61f0c04673dfb262ef6912eb2df39120[17]  <= 1'b0;
            I8f906015dba99b4a73dcf767cbd948ee[18]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I61f0c04673dfb262ef6912eb2df39120[18]  <= 1'b0;
            I8f906015dba99b4a73dcf767cbd948ee[19]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I61f0c04673dfb262ef6912eb2df39120[19]  <= 1'b0;
            I8f906015dba99b4a73dcf767cbd948ee[20]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I61f0c04673dfb262ef6912eb2df39120[20]  <= 1'b0;
            I8f906015dba99b4a73dcf767cbd948ee[21]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I61f0c04673dfb262ef6912eb2df39120[21]  <= 1'b0;
            I8f906015dba99b4a73dcf767cbd948ee[22]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I61f0c04673dfb262ef6912eb2df39120[22]  <= 1'b0;
            I7fa3f2648baacebf9e4b59c179601fa6                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I9ab4bbe4191d0f284defcdce6b885054[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibeb5edab51cd6aedad9c2ecedaded6f5[0]  <= 1'b0;
            I9ab4bbe4191d0f284defcdce6b885054[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibeb5edab51cd6aedad9c2ecedaded6f5[1]  <= 1'b0;
            I9ab4bbe4191d0f284defcdce6b885054[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibeb5edab51cd6aedad9c2ecedaded6f5[2]  <= 1'b0;
            I9ab4bbe4191d0f284defcdce6b885054[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibeb5edab51cd6aedad9c2ecedaded6f5[3]  <= 1'b0;
            I9ab4bbe4191d0f284defcdce6b885054[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibeb5edab51cd6aedad9c2ecedaded6f5[4]  <= 1'b0;
            I9ab4bbe4191d0f284defcdce6b885054[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibeb5edab51cd6aedad9c2ecedaded6f5[5]  <= 1'b0;
            I9ab4bbe4191d0f284defcdce6b885054[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibeb5edab51cd6aedad9c2ecedaded6f5[6]  <= 1'b0;
            I9ab4bbe4191d0f284defcdce6b885054[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibeb5edab51cd6aedad9c2ecedaded6f5[7]  <= 1'b0;
            I9ab4bbe4191d0f284defcdce6b885054[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibeb5edab51cd6aedad9c2ecedaded6f5[8]  <= 1'b0;
            I9ab4bbe4191d0f284defcdce6b885054[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibeb5edab51cd6aedad9c2ecedaded6f5[9]  <= 1'b0;
            I9ab4bbe4191d0f284defcdce6b885054[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibeb5edab51cd6aedad9c2ecedaded6f5[10]  <= 1'b0;
            I9ab4bbe4191d0f284defcdce6b885054[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibeb5edab51cd6aedad9c2ecedaded6f5[11]  <= 1'b0;
            I9ab4bbe4191d0f284defcdce6b885054[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibeb5edab51cd6aedad9c2ecedaded6f5[12]  <= 1'b0;
            I9ab4bbe4191d0f284defcdce6b885054[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibeb5edab51cd6aedad9c2ecedaded6f5[13]  <= 1'b0;
            I9ab4bbe4191d0f284defcdce6b885054[14]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibeb5edab51cd6aedad9c2ecedaded6f5[14]  <= 1'b0;
            I9ab4bbe4191d0f284defcdce6b885054[15]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibeb5edab51cd6aedad9c2ecedaded6f5[15]  <= 1'b0;
            I9ab4bbe4191d0f284defcdce6b885054[16]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibeb5edab51cd6aedad9c2ecedaded6f5[16]  <= 1'b0;
            I9ab4bbe4191d0f284defcdce6b885054[17]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibeb5edab51cd6aedad9c2ecedaded6f5[17]  <= 1'b0;
            I9ab4bbe4191d0f284defcdce6b885054[18]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibeb5edab51cd6aedad9c2ecedaded6f5[18]  <= 1'b0;
            I9ab4bbe4191d0f284defcdce6b885054[19]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibeb5edab51cd6aedad9c2ecedaded6f5[19]  <= 1'b0;
            I9ab4bbe4191d0f284defcdce6b885054[20]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibeb5edab51cd6aedad9c2ecedaded6f5[20]  <= 1'b0;
            I9ab4bbe4191d0f284defcdce6b885054[21]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibeb5edab51cd6aedad9c2ecedaded6f5[21]  <= 1'b0;
            I9ab4bbe4191d0f284defcdce6b885054[22]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibeb5edab51cd6aedad9c2ecedaded6f5[22]  <= 1'b0;
            Id7699f8f89380c315303644fdebacb32                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[0]  <= 1'b0;
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[1]  <= 1'b0;
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[2]  <= 1'b0;
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[3]  <= 1'b0;
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[4]  <= 1'b0;
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[5]  <= 1'b0;
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[6]  <= 1'b0;
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[7]  <= 1'b0;
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[8]  <= 1'b0;
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[9]  <= 1'b0;
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[10]  <= 1'b0;
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[11]  <= 1'b0;
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[12]  <= 1'b0;
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[13]  <= 1'b0;
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[14]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[14]  <= 1'b0;
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[15]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[15]  <= 1'b0;
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[16]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[16]  <= 1'b0;
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[17]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[17]  <= 1'b0;
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[18]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[18]  <= 1'b0;
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[19]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[19]  <= 1'b0;
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[20]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[20]  <= 1'b0;
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[21]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[21]  <= 1'b0;
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[22]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[22]  <= 1'b0;
            Ibf3e1ead3776901898d4b154aeb61267                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I6ff6fafd1a3364131b269724ad273ba5[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b7caaeb34c43e66e8d095a859e708fe[0]  <= 1'b0;
            I6ff6fafd1a3364131b269724ad273ba5[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b7caaeb34c43e66e8d095a859e708fe[1]  <= 1'b0;
            I6ff6fafd1a3364131b269724ad273ba5[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b7caaeb34c43e66e8d095a859e708fe[2]  <= 1'b0;
            I6ff6fafd1a3364131b269724ad273ba5[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b7caaeb34c43e66e8d095a859e708fe[3]  <= 1'b0;
            I6ff6fafd1a3364131b269724ad273ba5[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b7caaeb34c43e66e8d095a859e708fe[4]  <= 1'b0;
            I6ff6fafd1a3364131b269724ad273ba5[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b7caaeb34c43e66e8d095a859e708fe[5]  <= 1'b0;
            I6ff6fafd1a3364131b269724ad273ba5[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b7caaeb34c43e66e8d095a859e708fe[6]  <= 1'b0;
            I6ff6fafd1a3364131b269724ad273ba5[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b7caaeb34c43e66e8d095a859e708fe[7]  <= 1'b0;
            I6ff6fafd1a3364131b269724ad273ba5[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b7caaeb34c43e66e8d095a859e708fe[8]  <= 1'b0;
            I6ff6fafd1a3364131b269724ad273ba5[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b7caaeb34c43e66e8d095a859e708fe[9]  <= 1'b0;
            I6ff6fafd1a3364131b269724ad273ba5[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b7caaeb34c43e66e8d095a859e708fe[10]  <= 1'b0;
            I6ff6fafd1a3364131b269724ad273ba5[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b7caaeb34c43e66e8d095a859e708fe[11]  <= 1'b0;
            I6ff6fafd1a3364131b269724ad273ba5[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b7caaeb34c43e66e8d095a859e708fe[12]  <= 1'b0;
            I6ff6fafd1a3364131b269724ad273ba5[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b7caaeb34c43e66e8d095a859e708fe[13]  <= 1'b0;
            I6ff6fafd1a3364131b269724ad273ba5[14]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b7caaeb34c43e66e8d095a859e708fe[14]  <= 1'b0;
            I6ff6fafd1a3364131b269724ad273ba5[15]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b7caaeb34c43e66e8d095a859e708fe[15]  <= 1'b0;
            I6ff6fafd1a3364131b269724ad273ba5[16]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b7caaeb34c43e66e8d095a859e708fe[16]  <= 1'b0;
            I6ff6fafd1a3364131b269724ad273ba5[17]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b7caaeb34c43e66e8d095a859e708fe[17]  <= 1'b0;
            I6ff6fafd1a3364131b269724ad273ba5[18]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b7caaeb34c43e66e8d095a859e708fe[18]  <= 1'b0;
            I6ff6fafd1a3364131b269724ad273ba5[19]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b7caaeb34c43e66e8d095a859e708fe[19]  <= 1'b0;
            I6ff6fafd1a3364131b269724ad273ba5[20]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b7caaeb34c43e66e8d095a859e708fe[20]  <= 1'b0;
            I6ff6fafd1a3364131b269724ad273ba5[21]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b7caaeb34c43e66e8d095a859e708fe[21]  <= 1'b0;
            I6ff6fafd1a3364131b269724ad273ba5[22]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b7caaeb34c43e66e8d095a859e708fe[22]  <= 1'b0;
            Ie486617fc1d6354c7f347692cdbd894d                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I154fcd3171f1231e825ee603d53ecfe8[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib0bf69cc797f330fb2546eb46d2d6f76[0]  <= 1'b0;
            I154fcd3171f1231e825ee603d53ecfe8[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib0bf69cc797f330fb2546eb46d2d6f76[1]  <= 1'b0;
            I154fcd3171f1231e825ee603d53ecfe8[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib0bf69cc797f330fb2546eb46d2d6f76[2]  <= 1'b0;
            I154fcd3171f1231e825ee603d53ecfe8[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib0bf69cc797f330fb2546eb46d2d6f76[3]  <= 1'b0;
            I154fcd3171f1231e825ee603d53ecfe8[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib0bf69cc797f330fb2546eb46d2d6f76[4]  <= 1'b0;
            I154fcd3171f1231e825ee603d53ecfe8[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib0bf69cc797f330fb2546eb46d2d6f76[5]  <= 1'b0;
            I154fcd3171f1231e825ee603d53ecfe8[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib0bf69cc797f330fb2546eb46d2d6f76[6]  <= 1'b0;
            I154fcd3171f1231e825ee603d53ecfe8[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib0bf69cc797f330fb2546eb46d2d6f76[7]  <= 1'b0;
            I154fcd3171f1231e825ee603d53ecfe8[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib0bf69cc797f330fb2546eb46d2d6f76[8]  <= 1'b0;
            I154fcd3171f1231e825ee603d53ecfe8[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib0bf69cc797f330fb2546eb46d2d6f76[9]  <= 1'b0;
            I7ba403c6745e7d026282ad704e065702                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I489e70342dbba4a551097e3064dc9835[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iec7404bc79c58d4d2538fcdf659e9134[0]  <= 1'b0;
            I489e70342dbba4a551097e3064dc9835[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iec7404bc79c58d4d2538fcdf659e9134[1]  <= 1'b0;
            I489e70342dbba4a551097e3064dc9835[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iec7404bc79c58d4d2538fcdf659e9134[2]  <= 1'b0;
            I489e70342dbba4a551097e3064dc9835[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iec7404bc79c58d4d2538fcdf659e9134[3]  <= 1'b0;
            I489e70342dbba4a551097e3064dc9835[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iec7404bc79c58d4d2538fcdf659e9134[4]  <= 1'b0;
            I489e70342dbba4a551097e3064dc9835[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iec7404bc79c58d4d2538fcdf659e9134[5]  <= 1'b0;
            I489e70342dbba4a551097e3064dc9835[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iec7404bc79c58d4d2538fcdf659e9134[6]  <= 1'b0;
            I489e70342dbba4a551097e3064dc9835[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iec7404bc79c58d4d2538fcdf659e9134[7]  <= 1'b0;
            I489e70342dbba4a551097e3064dc9835[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iec7404bc79c58d4d2538fcdf659e9134[8]  <= 1'b0;
            I489e70342dbba4a551097e3064dc9835[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iec7404bc79c58d4d2538fcdf659e9134[9]  <= 1'b0;
            I93cb3974b8594665b2e7ce5593fde69b                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I0b0a1f577a212bd9024c8b9a44c92e00[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie1cd04c7668d3f450c387a6c1ad778c7[0]  <= 1'b0;
            I0b0a1f577a212bd9024c8b9a44c92e00[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie1cd04c7668d3f450c387a6c1ad778c7[1]  <= 1'b0;
            I0b0a1f577a212bd9024c8b9a44c92e00[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie1cd04c7668d3f450c387a6c1ad778c7[2]  <= 1'b0;
            I0b0a1f577a212bd9024c8b9a44c92e00[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie1cd04c7668d3f450c387a6c1ad778c7[3]  <= 1'b0;
            I0b0a1f577a212bd9024c8b9a44c92e00[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie1cd04c7668d3f450c387a6c1ad778c7[4]  <= 1'b0;
            I0b0a1f577a212bd9024c8b9a44c92e00[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie1cd04c7668d3f450c387a6c1ad778c7[5]  <= 1'b0;
            I0b0a1f577a212bd9024c8b9a44c92e00[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie1cd04c7668d3f450c387a6c1ad778c7[6]  <= 1'b0;
            I0b0a1f577a212bd9024c8b9a44c92e00[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie1cd04c7668d3f450c387a6c1ad778c7[7]  <= 1'b0;
            I0b0a1f577a212bd9024c8b9a44c92e00[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie1cd04c7668d3f450c387a6c1ad778c7[8]  <= 1'b0;
            I0b0a1f577a212bd9024c8b9a44c92e00[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie1cd04c7668d3f450c387a6c1ad778c7[9]  <= 1'b0;
            Id6a9ab06d58c3a01e1fe04fcf61406fd                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I40d311bab75b73e3788c50115a205270[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If511a6ea6aa5cda5353658d8e192791f[0]  <= 1'b0;
            I40d311bab75b73e3788c50115a205270[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If511a6ea6aa5cda5353658d8e192791f[1]  <= 1'b0;
            I40d311bab75b73e3788c50115a205270[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If511a6ea6aa5cda5353658d8e192791f[2]  <= 1'b0;
            I40d311bab75b73e3788c50115a205270[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If511a6ea6aa5cda5353658d8e192791f[3]  <= 1'b0;
            I40d311bab75b73e3788c50115a205270[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If511a6ea6aa5cda5353658d8e192791f[4]  <= 1'b0;
            I40d311bab75b73e3788c50115a205270[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If511a6ea6aa5cda5353658d8e192791f[5]  <= 1'b0;
            I40d311bab75b73e3788c50115a205270[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If511a6ea6aa5cda5353658d8e192791f[6]  <= 1'b0;
            I40d311bab75b73e3788c50115a205270[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If511a6ea6aa5cda5353658d8e192791f[7]  <= 1'b0;
            I40d311bab75b73e3788c50115a205270[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If511a6ea6aa5cda5353658d8e192791f[8]  <= 1'b0;
            I40d311bab75b73e3788c50115a205270[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If511a6ea6aa5cda5353658d8e192791f[9]  <= 1'b0;
            I261bd53528b82128acabd405389c8d60                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I5fa015a360308bffc46921d119b60c1b[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id88b9265ff08e0730e6a41abe1f80a32[0]  <= 1'b0;
            I5fa015a360308bffc46921d119b60c1b[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id88b9265ff08e0730e6a41abe1f80a32[1]  <= 1'b0;
            I5fa015a360308bffc46921d119b60c1b[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id88b9265ff08e0730e6a41abe1f80a32[2]  <= 1'b0;
            I5fa015a360308bffc46921d119b60c1b[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id88b9265ff08e0730e6a41abe1f80a32[3]  <= 1'b0;
            I5fa015a360308bffc46921d119b60c1b[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id88b9265ff08e0730e6a41abe1f80a32[4]  <= 1'b0;
            If7fa833bf1b1438e7a5bc783ee745252                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I9e42bc767599ce3cc4e2d886e5ef2e62[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6330943c9295298c53e889d47c7904d9[0]  <= 1'b0;
            I9e42bc767599ce3cc4e2d886e5ef2e62[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6330943c9295298c53e889d47c7904d9[1]  <= 1'b0;
            I9e42bc767599ce3cc4e2d886e5ef2e62[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6330943c9295298c53e889d47c7904d9[2]  <= 1'b0;
            I9e42bc767599ce3cc4e2d886e5ef2e62[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6330943c9295298c53e889d47c7904d9[3]  <= 1'b0;
            I9e42bc767599ce3cc4e2d886e5ef2e62[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6330943c9295298c53e889d47c7904d9[4]  <= 1'b0;
            Ibb103853fc21f8f3d466ca16557ccd3e                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Iea43b150eabf3c7781275821eee3e0c1[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5686b595177e07dd5bf231a35ee41659[0]  <= 1'b0;
            Iea43b150eabf3c7781275821eee3e0c1[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5686b595177e07dd5bf231a35ee41659[1]  <= 1'b0;
            Iea43b150eabf3c7781275821eee3e0c1[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5686b595177e07dd5bf231a35ee41659[2]  <= 1'b0;
            Iea43b150eabf3c7781275821eee3e0c1[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5686b595177e07dd5bf231a35ee41659[3]  <= 1'b0;
            Iea43b150eabf3c7781275821eee3e0c1[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5686b595177e07dd5bf231a35ee41659[4]  <= 1'b0;
            I37446eb66ccfd268cb418655b8160fe1                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I8012eea3d53fa4e000eb28b121e02ada[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9c0b88a0be66d62f8ab061aeaee7e60f[0]  <= 1'b0;
            I8012eea3d53fa4e000eb28b121e02ada[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9c0b88a0be66d62f8ab061aeaee7e60f[1]  <= 1'b0;
            I8012eea3d53fa4e000eb28b121e02ada[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9c0b88a0be66d62f8ab061aeaee7e60f[2]  <= 1'b0;
            I8012eea3d53fa4e000eb28b121e02ada[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9c0b88a0be66d62f8ab061aeaee7e60f[3]  <= 1'b0;
            I8012eea3d53fa4e000eb28b121e02ada[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9c0b88a0be66d62f8ab061aeaee7e60f[4]  <= 1'b0;
            Id17f6250f8c7f1d7f75fd27f92698da3                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I49804415d20c0c087f802b25dd609887[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9ef21ef20099af28d9a8c794f70d45a5[0]  <= 1'b0;
            I49804415d20c0c087f802b25dd609887[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9ef21ef20099af28d9a8c794f70d45a5[1]  <= 1'b0;
            I49804415d20c0c087f802b25dd609887[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9ef21ef20099af28d9a8c794f70d45a5[2]  <= 1'b0;
            I49804415d20c0c087f802b25dd609887[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9ef21ef20099af28d9a8c794f70d45a5[3]  <= 1'b0;
            I49804415d20c0c087f802b25dd609887[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9ef21ef20099af28d9a8c794f70d45a5[4]  <= 1'b0;
            I9957b02e8d0d888e6950eb553d9084d7                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Id270f05bf5c3fc0bb211d1665d149044[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic2941d16ae6a5cbce70e8546a18ca4ff[0]  <= 1'b0;
            Id270f05bf5c3fc0bb211d1665d149044[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic2941d16ae6a5cbce70e8546a18ca4ff[1]  <= 1'b0;
            Id270f05bf5c3fc0bb211d1665d149044[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic2941d16ae6a5cbce70e8546a18ca4ff[2]  <= 1'b0;
            Id270f05bf5c3fc0bb211d1665d149044[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic2941d16ae6a5cbce70e8546a18ca4ff[3]  <= 1'b0;
            Id270f05bf5c3fc0bb211d1665d149044[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic2941d16ae6a5cbce70e8546a18ca4ff[4]  <= 1'b0;
            Ic71258b745437bc8463fb4f847c55e27                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            If091fe044c792be711325c103b84cf1d[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8e29ebe9ee25ea8ef3e52ff56fc29157[0]  <= 1'b0;
            If091fe044c792be711325c103b84cf1d[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8e29ebe9ee25ea8ef3e52ff56fc29157[1]  <= 1'b0;
            If091fe044c792be711325c103b84cf1d[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8e29ebe9ee25ea8ef3e52ff56fc29157[2]  <= 1'b0;
            If091fe044c792be711325c103b84cf1d[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8e29ebe9ee25ea8ef3e52ff56fc29157[3]  <= 1'b0;
            If091fe044c792be711325c103b84cf1d[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8e29ebe9ee25ea8ef3e52ff56fc29157[4]  <= 1'b0;
            I24bb5c315eacf0f4e8c86f6582389e39                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I1550db301291ab131a5536147fb938f6[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic3742290179b27b9865f9d1f88d66266[0]  <= 1'b0;
            I1550db301291ab131a5536147fb938f6[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic3742290179b27b9865f9d1f88d66266[1]  <= 1'b0;
            I1550db301291ab131a5536147fb938f6[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic3742290179b27b9865f9d1f88d66266[2]  <= 1'b0;
            I1550db301291ab131a5536147fb938f6[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic3742290179b27b9865f9d1f88d66266[3]  <= 1'b0;
            I1550db301291ab131a5536147fb938f6[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic3742290179b27b9865f9d1f88d66266[4]  <= 1'b0;
            I607f203694ff76930cfee4103cb73c30                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I74d1345ee56f5688f875823a5d7c1f4f[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I04302edb2671c5bc0ca2673cd53935e1[0]  <= 1'b0;
            I74d1345ee56f5688f875823a5d7c1f4f[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I04302edb2671c5bc0ca2673cd53935e1[1]  <= 1'b0;
            I74d1345ee56f5688f875823a5d7c1f4f[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I04302edb2671c5bc0ca2673cd53935e1[2]  <= 1'b0;
            I74d1345ee56f5688f875823a5d7c1f4f[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I04302edb2671c5bc0ca2673cd53935e1[3]  <= 1'b0;
            I74d1345ee56f5688f875823a5d7c1f4f[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I04302edb2671c5bc0ca2673cd53935e1[4]  <= 1'b0;
            I74d1345ee56f5688f875823a5d7c1f4f[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I04302edb2671c5bc0ca2673cd53935e1[5]  <= 1'b0;
            I74d1345ee56f5688f875823a5d7c1f4f[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I04302edb2671c5bc0ca2673cd53935e1[6]  <= 1'b0;
            I74d1345ee56f5688f875823a5d7c1f4f[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I04302edb2671c5bc0ca2673cd53935e1[7]  <= 1'b0;
            I74d1345ee56f5688f875823a5d7c1f4f[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I04302edb2671c5bc0ca2673cd53935e1[8]  <= 1'b0;
            I74d1345ee56f5688f875823a5d7c1f4f[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I04302edb2671c5bc0ca2673cd53935e1[9]  <= 1'b0;
            I74d1345ee56f5688f875823a5d7c1f4f[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I04302edb2671c5bc0ca2673cd53935e1[10]  <= 1'b0;
            I74d1345ee56f5688f875823a5d7c1f4f[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I04302edb2671c5bc0ca2673cd53935e1[11]  <= 1'b0;
            I74d1345ee56f5688f875823a5d7c1f4f[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I04302edb2671c5bc0ca2673cd53935e1[12]  <= 1'b0;
            I74d1345ee56f5688f875823a5d7c1f4f[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I04302edb2671c5bc0ca2673cd53935e1[13]  <= 1'b0;
            Ica8e4c56ebb37e189ca8e6b3daafdb80                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I187371a49a27a988920854b2bb61bea5[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I480a0f6d6c3eb936de10a72749f6cd3f[0]  <= 1'b0;
            I187371a49a27a988920854b2bb61bea5[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I480a0f6d6c3eb936de10a72749f6cd3f[1]  <= 1'b0;
            I187371a49a27a988920854b2bb61bea5[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I480a0f6d6c3eb936de10a72749f6cd3f[2]  <= 1'b0;
            I187371a49a27a988920854b2bb61bea5[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I480a0f6d6c3eb936de10a72749f6cd3f[3]  <= 1'b0;
            I187371a49a27a988920854b2bb61bea5[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I480a0f6d6c3eb936de10a72749f6cd3f[4]  <= 1'b0;
            I187371a49a27a988920854b2bb61bea5[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I480a0f6d6c3eb936de10a72749f6cd3f[5]  <= 1'b0;
            I187371a49a27a988920854b2bb61bea5[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I480a0f6d6c3eb936de10a72749f6cd3f[6]  <= 1'b0;
            I187371a49a27a988920854b2bb61bea5[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I480a0f6d6c3eb936de10a72749f6cd3f[7]  <= 1'b0;
            I187371a49a27a988920854b2bb61bea5[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I480a0f6d6c3eb936de10a72749f6cd3f[8]  <= 1'b0;
            I187371a49a27a988920854b2bb61bea5[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I480a0f6d6c3eb936de10a72749f6cd3f[9]  <= 1'b0;
            I187371a49a27a988920854b2bb61bea5[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I480a0f6d6c3eb936de10a72749f6cd3f[10]  <= 1'b0;
            I187371a49a27a988920854b2bb61bea5[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I480a0f6d6c3eb936de10a72749f6cd3f[11]  <= 1'b0;
            I187371a49a27a988920854b2bb61bea5[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I480a0f6d6c3eb936de10a72749f6cd3f[12]  <= 1'b0;
            I187371a49a27a988920854b2bb61bea5[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I480a0f6d6c3eb936de10a72749f6cd3f[13]  <= 1'b0;
            I7089386c94261e0febf3b4f7dc1aec30                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I48c4c6e7414394e3aeff9d17ec25d020[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I50976b0051e84b6a42fc1dbabd7d20ae[0]  <= 1'b0;
            I48c4c6e7414394e3aeff9d17ec25d020[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I50976b0051e84b6a42fc1dbabd7d20ae[1]  <= 1'b0;
            I48c4c6e7414394e3aeff9d17ec25d020[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I50976b0051e84b6a42fc1dbabd7d20ae[2]  <= 1'b0;
            I48c4c6e7414394e3aeff9d17ec25d020[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I50976b0051e84b6a42fc1dbabd7d20ae[3]  <= 1'b0;
            I48c4c6e7414394e3aeff9d17ec25d020[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I50976b0051e84b6a42fc1dbabd7d20ae[4]  <= 1'b0;
            I48c4c6e7414394e3aeff9d17ec25d020[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I50976b0051e84b6a42fc1dbabd7d20ae[5]  <= 1'b0;
            I48c4c6e7414394e3aeff9d17ec25d020[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I50976b0051e84b6a42fc1dbabd7d20ae[6]  <= 1'b0;
            I48c4c6e7414394e3aeff9d17ec25d020[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I50976b0051e84b6a42fc1dbabd7d20ae[7]  <= 1'b0;
            I48c4c6e7414394e3aeff9d17ec25d020[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I50976b0051e84b6a42fc1dbabd7d20ae[8]  <= 1'b0;
            I48c4c6e7414394e3aeff9d17ec25d020[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I50976b0051e84b6a42fc1dbabd7d20ae[9]  <= 1'b0;
            I48c4c6e7414394e3aeff9d17ec25d020[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I50976b0051e84b6a42fc1dbabd7d20ae[10]  <= 1'b0;
            I48c4c6e7414394e3aeff9d17ec25d020[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I50976b0051e84b6a42fc1dbabd7d20ae[11]  <= 1'b0;
            I48c4c6e7414394e3aeff9d17ec25d020[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I50976b0051e84b6a42fc1dbabd7d20ae[12]  <= 1'b0;
            I48c4c6e7414394e3aeff9d17ec25d020[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I50976b0051e84b6a42fc1dbabd7d20ae[13]  <= 1'b0;
            Ia1e4f20f32f7371cb0078d6e80fe8b7e                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I3cba0f4c2ca8c7c200df8e1071ab429d[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I82e0e091fba6f79cef97eacac4b43ecb[0]  <= 1'b0;
            I3cba0f4c2ca8c7c200df8e1071ab429d[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I82e0e091fba6f79cef97eacac4b43ecb[1]  <= 1'b0;
            I3cba0f4c2ca8c7c200df8e1071ab429d[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I82e0e091fba6f79cef97eacac4b43ecb[2]  <= 1'b0;
            I3cba0f4c2ca8c7c200df8e1071ab429d[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I82e0e091fba6f79cef97eacac4b43ecb[3]  <= 1'b0;
            I3cba0f4c2ca8c7c200df8e1071ab429d[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I82e0e091fba6f79cef97eacac4b43ecb[4]  <= 1'b0;
            I3cba0f4c2ca8c7c200df8e1071ab429d[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I82e0e091fba6f79cef97eacac4b43ecb[5]  <= 1'b0;
            I3cba0f4c2ca8c7c200df8e1071ab429d[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I82e0e091fba6f79cef97eacac4b43ecb[6]  <= 1'b0;
            I3cba0f4c2ca8c7c200df8e1071ab429d[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I82e0e091fba6f79cef97eacac4b43ecb[7]  <= 1'b0;
            I3cba0f4c2ca8c7c200df8e1071ab429d[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I82e0e091fba6f79cef97eacac4b43ecb[8]  <= 1'b0;
            I3cba0f4c2ca8c7c200df8e1071ab429d[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I82e0e091fba6f79cef97eacac4b43ecb[9]  <= 1'b0;
            I3cba0f4c2ca8c7c200df8e1071ab429d[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I82e0e091fba6f79cef97eacac4b43ecb[10]  <= 1'b0;
            I3cba0f4c2ca8c7c200df8e1071ab429d[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I82e0e091fba6f79cef97eacac4b43ecb[11]  <= 1'b0;
            I3cba0f4c2ca8c7c200df8e1071ab429d[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I82e0e091fba6f79cef97eacac4b43ecb[12]  <= 1'b0;
            I3cba0f4c2ca8c7c200df8e1071ab429d[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I82e0e091fba6f79cef97eacac4b43ecb[13]  <= 1'b0;
            I790cbca796af58b1726d0a4680cc164f                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I35688678e1a83ec39d737d9cdfd44ba3[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I3d50cfeaa4b69c09bb648b8873a6bc24[0]  <= 1'b0;
            I35688678e1a83ec39d737d9cdfd44ba3[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I3d50cfeaa4b69c09bb648b8873a6bc24[1]  <= 1'b0;
            I35688678e1a83ec39d737d9cdfd44ba3[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I3d50cfeaa4b69c09bb648b8873a6bc24[2]  <= 1'b0;
            I35688678e1a83ec39d737d9cdfd44ba3[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I3d50cfeaa4b69c09bb648b8873a6bc24[3]  <= 1'b0;
            I35688678e1a83ec39d737d9cdfd44ba3[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I3d50cfeaa4b69c09bb648b8873a6bc24[4]  <= 1'b0;
            I35688678e1a83ec39d737d9cdfd44ba3[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I3d50cfeaa4b69c09bb648b8873a6bc24[5]  <= 1'b0;
            I35688678e1a83ec39d737d9cdfd44ba3[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I3d50cfeaa4b69c09bb648b8873a6bc24[6]  <= 1'b0;
            I0a93f095f9efb1542116a295c0db9c8b                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I94b86d31e8226723950096e91855b6d3[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I33a6ffad80ddf99a4d316a049078244d[0]  <= 1'b0;
            I94b86d31e8226723950096e91855b6d3[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I33a6ffad80ddf99a4d316a049078244d[1]  <= 1'b0;
            I94b86d31e8226723950096e91855b6d3[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I33a6ffad80ddf99a4d316a049078244d[2]  <= 1'b0;
            I94b86d31e8226723950096e91855b6d3[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I33a6ffad80ddf99a4d316a049078244d[3]  <= 1'b0;
            I94b86d31e8226723950096e91855b6d3[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I33a6ffad80ddf99a4d316a049078244d[4]  <= 1'b0;
            I94b86d31e8226723950096e91855b6d3[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I33a6ffad80ddf99a4d316a049078244d[5]  <= 1'b0;
            I94b86d31e8226723950096e91855b6d3[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I33a6ffad80ddf99a4d316a049078244d[6]  <= 1'b0;
            I989ba39f188a44475a83e65a4960d2af                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I0ea7c4721ee0c13ad15a9b0fa7b15ad3[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I980165c1147ac5ff86619c841c6031dc[0]  <= 1'b0;
            I0ea7c4721ee0c13ad15a9b0fa7b15ad3[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I980165c1147ac5ff86619c841c6031dc[1]  <= 1'b0;
            I0ea7c4721ee0c13ad15a9b0fa7b15ad3[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I980165c1147ac5ff86619c841c6031dc[2]  <= 1'b0;
            I0ea7c4721ee0c13ad15a9b0fa7b15ad3[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I980165c1147ac5ff86619c841c6031dc[3]  <= 1'b0;
            I0ea7c4721ee0c13ad15a9b0fa7b15ad3[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I980165c1147ac5ff86619c841c6031dc[4]  <= 1'b0;
            I0ea7c4721ee0c13ad15a9b0fa7b15ad3[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I980165c1147ac5ff86619c841c6031dc[5]  <= 1'b0;
            I0ea7c4721ee0c13ad15a9b0fa7b15ad3[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I980165c1147ac5ff86619c841c6031dc[6]  <= 1'b0;
            I9bcc1d9b3dd258fa7b6042f0185d48cb                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I29dd5fb1c2673cd4daa9cafaf24d8e7c[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I19df055705f322292a3601fa63f0e5f9[0]  <= 1'b0;
            I29dd5fb1c2673cd4daa9cafaf24d8e7c[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I19df055705f322292a3601fa63f0e5f9[1]  <= 1'b0;
            I29dd5fb1c2673cd4daa9cafaf24d8e7c[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I19df055705f322292a3601fa63f0e5f9[2]  <= 1'b0;
            I29dd5fb1c2673cd4daa9cafaf24d8e7c[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I19df055705f322292a3601fa63f0e5f9[3]  <= 1'b0;
            I29dd5fb1c2673cd4daa9cafaf24d8e7c[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I19df055705f322292a3601fa63f0e5f9[4]  <= 1'b0;
            I29dd5fb1c2673cd4daa9cafaf24d8e7c[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I19df055705f322292a3601fa63f0e5f9[5]  <= 1'b0;
            I29dd5fb1c2673cd4daa9cafaf24d8e7c[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I19df055705f322292a3601fa63f0e5f9[6]  <= 1'b0;
            I9ba14715d9f33ef45681ad52f5be9593                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Iead4c81d836e3befae55049797c30d6b[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0e0b15868b02ca52b260f17f150d237e[0]  <= 1'b0;
            Iead4c81d836e3befae55049797c30d6b[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0e0b15868b02ca52b260f17f150d237e[1]  <= 1'b0;
            Iead4c81d836e3befae55049797c30d6b[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0e0b15868b02ca52b260f17f150d237e[2]  <= 1'b0;
            Iead4c81d836e3befae55049797c30d6b[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0e0b15868b02ca52b260f17f150d237e[3]  <= 1'b0;
            Iead4c81d836e3befae55049797c30d6b[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0e0b15868b02ca52b260f17f150d237e[4]  <= 1'b0;
            Iead4c81d836e3befae55049797c30d6b[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0e0b15868b02ca52b260f17f150d237e[5]  <= 1'b0;
            Iead4c81d836e3befae55049797c30d6b[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0e0b15868b02ca52b260f17f150d237e[6]  <= 1'b0;
            Iead4c81d836e3befae55049797c30d6b[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0e0b15868b02ca52b260f17f150d237e[7]  <= 1'b0;
            Iead4c81d836e3befae55049797c30d6b[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0e0b15868b02ca52b260f17f150d237e[8]  <= 1'b0;
            Iead4c81d836e3befae55049797c30d6b[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0e0b15868b02ca52b260f17f150d237e[9]  <= 1'b0;
            Iead4c81d836e3befae55049797c30d6b[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0e0b15868b02ca52b260f17f150d237e[10]  <= 1'b0;
            Iead4c81d836e3befae55049797c30d6b[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0e0b15868b02ca52b260f17f150d237e[11]  <= 1'b0;
            Iead4c81d836e3befae55049797c30d6b[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0e0b15868b02ca52b260f17f150d237e[12]  <= 1'b0;
            I396a897f79b519f4fa02af39d0274f64                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I23e22f44791c167acaba27c91ef3b497[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[0]  <= 1'b0;
            I23e22f44791c167acaba27c91ef3b497[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[1]  <= 1'b0;
            I23e22f44791c167acaba27c91ef3b497[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[2]  <= 1'b0;
            I23e22f44791c167acaba27c91ef3b497[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[3]  <= 1'b0;
            I23e22f44791c167acaba27c91ef3b497[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[4]  <= 1'b0;
            I23e22f44791c167acaba27c91ef3b497[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[5]  <= 1'b0;
            I23e22f44791c167acaba27c91ef3b497[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[6]  <= 1'b0;
            I23e22f44791c167acaba27c91ef3b497[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[7]  <= 1'b0;
            I23e22f44791c167acaba27c91ef3b497[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[8]  <= 1'b0;
            I23e22f44791c167acaba27c91ef3b497[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[9]  <= 1'b0;
            I23e22f44791c167acaba27c91ef3b497[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[10]  <= 1'b0;
            I23e22f44791c167acaba27c91ef3b497[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[11]  <= 1'b0;
            I23e22f44791c167acaba27c91ef3b497[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[12]  <= 1'b0;
            I197c0cd576e16ee2197a28c86397f801                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ic91f087829e0b9e0c964229a2dc567bc[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8e591d83170c8ba46d31c61935311b22[0]  <= 1'b0;
            Ic91f087829e0b9e0c964229a2dc567bc[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8e591d83170c8ba46d31c61935311b22[1]  <= 1'b0;
            Ic91f087829e0b9e0c964229a2dc567bc[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8e591d83170c8ba46d31c61935311b22[2]  <= 1'b0;
            Ic91f087829e0b9e0c964229a2dc567bc[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8e591d83170c8ba46d31c61935311b22[3]  <= 1'b0;
            Ic91f087829e0b9e0c964229a2dc567bc[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8e591d83170c8ba46d31c61935311b22[4]  <= 1'b0;
            Ic91f087829e0b9e0c964229a2dc567bc[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8e591d83170c8ba46d31c61935311b22[5]  <= 1'b0;
            Ic91f087829e0b9e0c964229a2dc567bc[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8e591d83170c8ba46d31c61935311b22[6]  <= 1'b0;
            Ic91f087829e0b9e0c964229a2dc567bc[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8e591d83170c8ba46d31c61935311b22[7]  <= 1'b0;
            Ic91f087829e0b9e0c964229a2dc567bc[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8e591d83170c8ba46d31c61935311b22[8]  <= 1'b0;
            Ic91f087829e0b9e0c964229a2dc567bc[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8e591d83170c8ba46d31c61935311b22[9]  <= 1'b0;
            Ic91f087829e0b9e0c964229a2dc567bc[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8e591d83170c8ba46d31c61935311b22[10]  <= 1'b0;
            Ic91f087829e0b9e0c964229a2dc567bc[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8e591d83170c8ba46d31c61935311b22[11]  <= 1'b0;
            Ic91f087829e0b9e0c964229a2dc567bc[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8e591d83170c8ba46d31c61935311b22[12]  <= 1'b0;
            I094a178e55425f27ac1ff6195217396b                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I0fd9bcdcf8faaaabf94649881419c66f[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I02b62fafd371de339f299f8aefec6c43[0]  <= 1'b0;
            I0fd9bcdcf8faaaabf94649881419c66f[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I02b62fafd371de339f299f8aefec6c43[1]  <= 1'b0;
            I0fd9bcdcf8faaaabf94649881419c66f[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I02b62fafd371de339f299f8aefec6c43[2]  <= 1'b0;
            I0fd9bcdcf8faaaabf94649881419c66f[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I02b62fafd371de339f299f8aefec6c43[3]  <= 1'b0;
            I0fd9bcdcf8faaaabf94649881419c66f[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I02b62fafd371de339f299f8aefec6c43[4]  <= 1'b0;
            I0fd9bcdcf8faaaabf94649881419c66f[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I02b62fafd371de339f299f8aefec6c43[5]  <= 1'b0;
            I0fd9bcdcf8faaaabf94649881419c66f[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I02b62fafd371de339f299f8aefec6c43[6]  <= 1'b0;
            I0fd9bcdcf8faaaabf94649881419c66f[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I02b62fafd371de339f299f8aefec6c43[7]  <= 1'b0;
            I0fd9bcdcf8faaaabf94649881419c66f[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I02b62fafd371de339f299f8aefec6c43[8]  <= 1'b0;
            I0fd9bcdcf8faaaabf94649881419c66f[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I02b62fafd371de339f299f8aefec6c43[9]  <= 1'b0;
            I0fd9bcdcf8faaaabf94649881419c66f[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I02b62fafd371de339f299f8aefec6c43[10]  <= 1'b0;
            I0fd9bcdcf8faaaabf94649881419c66f[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I02b62fafd371de339f299f8aefec6c43[11]  <= 1'b0;
            I0fd9bcdcf8faaaabf94649881419c66f[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I02b62fafd371de339f299f8aefec6c43[12]  <= 1'b0;
            I3177408f7d08b431be99297fb10586e6                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I7cbcdd5018de9ceb49554b140e5665e8[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6ebab438dc55ccf6c1600313891d9c38[0]  <= 1'b0;
            I7cbcdd5018de9ceb49554b140e5665e8[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6ebab438dc55ccf6c1600313891d9c38[1]  <= 1'b0;
            I7cbcdd5018de9ceb49554b140e5665e8[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6ebab438dc55ccf6c1600313891d9c38[2]  <= 1'b0;
            I7cbcdd5018de9ceb49554b140e5665e8[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6ebab438dc55ccf6c1600313891d9c38[3]  <= 1'b0;
            I7cbcdd5018de9ceb49554b140e5665e8[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6ebab438dc55ccf6c1600313891d9c38[4]  <= 1'b0;
            I7cbcdd5018de9ceb49554b140e5665e8[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6ebab438dc55ccf6c1600313891d9c38[5]  <= 1'b0;
            Id4948c876d48bdbf317d32f135e645b4                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I5a79c19fd2093d974b574e85245b5617[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I2fbf89398a148c47810456812dbee5a6[0]  <= 1'b0;
            I5a79c19fd2093d974b574e85245b5617[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I2fbf89398a148c47810456812dbee5a6[1]  <= 1'b0;
            I5a79c19fd2093d974b574e85245b5617[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I2fbf89398a148c47810456812dbee5a6[2]  <= 1'b0;
            I5a79c19fd2093d974b574e85245b5617[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I2fbf89398a148c47810456812dbee5a6[3]  <= 1'b0;
            I5a79c19fd2093d974b574e85245b5617[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I2fbf89398a148c47810456812dbee5a6[4]  <= 1'b0;
            I5a79c19fd2093d974b574e85245b5617[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I2fbf89398a148c47810456812dbee5a6[5]  <= 1'b0;
            Ice5ff01d4fb4583898498651a0ac0171                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ica937143b618734fa099683949153130[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icac5a9001ee113e612e3457b4b49ee68[0]  <= 1'b0;
            Ica937143b618734fa099683949153130[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icac5a9001ee113e612e3457b4b49ee68[1]  <= 1'b0;
            Ica937143b618734fa099683949153130[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icac5a9001ee113e612e3457b4b49ee68[2]  <= 1'b0;
            Ica937143b618734fa099683949153130[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icac5a9001ee113e612e3457b4b49ee68[3]  <= 1'b0;
            Ica937143b618734fa099683949153130[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icac5a9001ee113e612e3457b4b49ee68[4]  <= 1'b0;
            Ica937143b618734fa099683949153130[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icac5a9001ee113e612e3457b4b49ee68[5]  <= 1'b0;
            I0fb33a5ced3d15622c9aefa188052e24                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I2d4d5d2694718b39e80b89b422d690cc[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9461e92a5880cb9e04fcece2ef4674f0[0]  <= 1'b0;
            I2d4d5d2694718b39e80b89b422d690cc[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9461e92a5880cb9e04fcece2ef4674f0[1]  <= 1'b0;
            I2d4d5d2694718b39e80b89b422d690cc[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9461e92a5880cb9e04fcece2ef4674f0[2]  <= 1'b0;
            I2d4d5d2694718b39e80b89b422d690cc[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9461e92a5880cb9e04fcece2ef4674f0[3]  <= 1'b0;
            I2d4d5d2694718b39e80b89b422d690cc[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9461e92a5880cb9e04fcece2ef4674f0[4]  <= 1'b0;
            I2d4d5d2694718b39e80b89b422d690cc[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9461e92a5880cb9e04fcece2ef4674f0[5]  <= 1'b0;
            I0074e1c3ca0ff903a9201ac5fe7ca841                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ic2faea3d4bb97dda16ecc29c27939ca6[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I07930a807994815de45864af579902c4[0]  <= 1'b0;
            Ic2faea3d4bb97dda16ecc29c27939ca6[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I07930a807994815de45864af579902c4[1]  <= 1'b0;
            Ic2faea3d4bb97dda16ecc29c27939ca6[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I07930a807994815de45864af579902c4[2]  <= 1'b0;
            Ic2faea3d4bb97dda16ecc29c27939ca6[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I07930a807994815de45864af579902c4[3]  <= 1'b0;
            Ic2faea3d4bb97dda16ecc29c27939ca6[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I07930a807994815de45864af579902c4[4]  <= 1'b0;
            Ic2faea3d4bb97dda16ecc29c27939ca6[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I07930a807994815de45864af579902c4[5]  <= 1'b0;
            Ic2faea3d4bb97dda16ecc29c27939ca6[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I07930a807994815de45864af579902c4[6]  <= 1'b0;
            Ic2faea3d4bb97dda16ecc29c27939ca6[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I07930a807994815de45864af579902c4[7]  <= 1'b0;
            If65f587e987a51c093e8dd4df532e26c                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I503e83a1146c42d5c1ef011ecb280807[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I72a2f42b727a0503d43332c0f22d5ae3[0]  <= 1'b0;
            I503e83a1146c42d5c1ef011ecb280807[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I72a2f42b727a0503d43332c0f22d5ae3[1]  <= 1'b0;
            I503e83a1146c42d5c1ef011ecb280807[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I72a2f42b727a0503d43332c0f22d5ae3[2]  <= 1'b0;
            I503e83a1146c42d5c1ef011ecb280807[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I72a2f42b727a0503d43332c0f22d5ae3[3]  <= 1'b0;
            I503e83a1146c42d5c1ef011ecb280807[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I72a2f42b727a0503d43332c0f22d5ae3[4]  <= 1'b0;
            I503e83a1146c42d5c1ef011ecb280807[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I72a2f42b727a0503d43332c0f22d5ae3[5]  <= 1'b0;
            I503e83a1146c42d5c1ef011ecb280807[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I72a2f42b727a0503d43332c0f22d5ae3[6]  <= 1'b0;
            I503e83a1146c42d5c1ef011ecb280807[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I72a2f42b727a0503d43332c0f22d5ae3[7]  <= 1'b0;
            I33d7e77d08590f0dfb1867e741dd8b6b                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ib9886c1fcd27ceb24afb2d0d7da85c26[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8b8b9c4777e6df3eb2b9313e69ef2c8c[0]  <= 1'b0;
            Ib9886c1fcd27ceb24afb2d0d7da85c26[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8b8b9c4777e6df3eb2b9313e69ef2c8c[1]  <= 1'b0;
            Ib9886c1fcd27ceb24afb2d0d7da85c26[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8b8b9c4777e6df3eb2b9313e69ef2c8c[2]  <= 1'b0;
            Ib9886c1fcd27ceb24afb2d0d7da85c26[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8b8b9c4777e6df3eb2b9313e69ef2c8c[3]  <= 1'b0;
            Ib9886c1fcd27ceb24afb2d0d7da85c26[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8b8b9c4777e6df3eb2b9313e69ef2c8c[4]  <= 1'b0;
            Ib9886c1fcd27ceb24afb2d0d7da85c26[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8b8b9c4777e6df3eb2b9313e69ef2c8c[5]  <= 1'b0;
            Ib9886c1fcd27ceb24afb2d0d7da85c26[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8b8b9c4777e6df3eb2b9313e69ef2c8c[6]  <= 1'b0;
            Ib9886c1fcd27ceb24afb2d0d7da85c26[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8b8b9c4777e6df3eb2b9313e69ef2c8c[7]  <= 1'b0;
            I678c22563e0273403b046df4261f21cf                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Icd90612c09423a2817a72f750e585309[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4a16e8e7946d9a8220304fc1be3fb362[0]  <= 1'b0;
            Icd90612c09423a2817a72f750e585309[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4a16e8e7946d9a8220304fc1be3fb362[1]  <= 1'b0;
            Icd90612c09423a2817a72f750e585309[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4a16e8e7946d9a8220304fc1be3fb362[2]  <= 1'b0;
            Icd90612c09423a2817a72f750e585309[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4a16e8e7946d9a8220304fc1be3fb362[3]  <= 1'b0;
            Icd90612c09423a2817a72f750e585309[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4a16e8e7946d9a8220304fc1be3fb362[4]  <= 1'b0;
            Icd90612c09423a2817a72f750e585309[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4a16e8e7946d9a8220304fc1be3fb362[5]  <= 1'b0;
            Icd90612c09423a2817a72f750e585309[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4a16e8e7946d9a8220304fc1be3fb362[6]  <= 1'b0;
            Icd90612c09423a2817a72f750e585309[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4a16e8e7946d9a8220304fc1be3fb362[7]  <= 1'b0;
            Icca700c12ae2e8155ca6b41e692e8a8c                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ib7b7884d2653893806af34579f7c0760[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic2580cbeec8c11a19bd1e2ebc29d255e[0]  <= 1'b0;
            Ib7b7884d2653893806af34579f7c0760[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic2580cbeec8c11a19bd1e2ebc29d255e[1]  <= 1'b0;
            Ib7b7884d2653893806af34579f7c0760[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic2580cbeec8c11a19bd1e2ebc29d255e[2]  <= 1'b0;
            Ib7b7884d2653893806af34579f7c0760[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic2580cbeec8c11a19bd1e2ebc29d255e[3]  <= 1'b0;
            Ib7b7884d2653893806af34579f7c0760[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic2580cbeec8c11a19bd1e2ebc29d255e[4]  <= 1'b0;
            Ib7b7884d2653893806af34579f7c0760[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic2580cbeec8c11a19bd1e2ebc29d255e[5]  <= 1'b0;
            Ib7b7884d2653893806af34579f7c0760[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic2580cbeec8c11a19bd1e2ebc29d255e[6]  <= 1'b0;
            Ib7b7884d2653893806af34579f7c0760[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic2580cbeec8c11a19bd1e2ebc29d255e[7]  <= 1'b0;
            Ib7b7884d2653893806af34579f7c0760[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic2580cbeec8c11a19bd1e2ebc29d255e[8]  <= 1'b0;
            I5ed74e81d2497681af5a0ca13fe23088                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ic3f0ad21d8a446c31afec49309a18133[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If79ed5ee2b8710da0608c1e245d07d55[0]  <= 1'b0;
            Ic3f0ad21d8a446c31afec49309a18133[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If79ed5ee2b8710da0608c1e245d07d55[1]  <= 1'b0;
            Ic3f0ad21d8a446c31afec49309a18133[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If79ed5ee2b8710da0608c1e245d07d55[2]  <= 1'b0;
            Ic3f0ad21d8a446c31afec49309a18133[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If79ed5ee2b8710da0608c1e245d07d55[3]  <= 1'b0;
            Ic3f0ad21d8a446c31afec49309a18133[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If79ed5ee2b8710da0608c1e245d07d55[4]  <= 1'b0;
            Ic3f0ad21d8a446c31afec49309a18133[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If79ed5ee2b8710da0608c1e245d07d55[5]  <= 1'b0;
            Ic3f0ad21d8a446c31afec49309a18133[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If79ed5ee2b8710da0608c1e245d07d55[6]  <= 1'b0;
            Ic3f0ad21d8a446c31afec49309a18133[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If79ed5ee2b8710da0608c1e245d07d55[7]  <= 1'b0;
            Ic3f0ad21d8a446c31afec49309a18133[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If79ed5ee2b8710da0608c1e245d07d55[8]  <= 1'b0;
            Ic7fa6b8cdfcf7d83d4e101d9c8b7b34f                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I2dd65bec7d2bc4778b7fc48a413d2ba7[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9497bbb4f746969a95cff948a3ee9ade[0]  <= 1'b0;
            I2dd65bec7d2bc4778b7fc48a413d2ba7[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9497bbb4f746969a95cff948a3ee9ade[1]  <= 1'b0;
            I2dd65bec7d2bc4778b7fc48a413d2ba7[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9497bbb4f746969a95cff948a3ee9ade[2]  <= 1'b0;
            I2dd65bec7d2bc4778b7fc48a413d2ba7[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9497bbb4f746969a95cff948a3ee9ade[3]  <= 1'b0;
            I2dd65bec7d2bc4778b7fc48a413d2ba7[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9497bbb4f746969a95cff948a3ee9ade[4]  <= 1'b0;
            I2dd65bec7d2bc4778b7fc48a413d2ba7[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9497bbb4f746969a95cff948a3ee9ade[5]  <= 1'b0;
            I2dd65bec7d2bc4778b7fc48a413d2ba7[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9497bbb4f746969a95cff948a3ee9ade[6]  <= 1'b0;
            I2dd65bec7d2bc4778b7fc48a413d2ba7[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9497bbb4f746969a95cff948a3ee9ade[7]  <= 1'b0;
            I2dd65bec7d2bc4778b7fc48a413d2ba7[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9497bbb4f746969a95cff948a3ee9ade[8]  <= 1'b0;
            I26010e26e22d8a2ea831e86fae34a24e                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I36b5867a3da6f2ed529e791166640d3f[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I651d700a00d7004d8728bc7356f30926[0]  <= 1'b0;
            I36b5867a3da6f2ed529e791166640d3f[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I651d700a00d7004d8728bc7356f30926[1]  <= 1'b0;
            I36b5867a3da6f2ed529e791166640d3f[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I651d700a00d7004d8728bc7356f30926[2]  <= 1'b0;
            I36b5867a3da6f2ed529e791166640d3f[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I651d700a00d7004d8728bc7356f30926[3]  <= 1'b0;
            I36b5867a3da6f2ed529e791166640d3f[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I651d700a00d7004d8728bc7356f30926[4]  <= 1'b0;
            I36b5867a3da6f2ed529e791166640d3f[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I651d700a00d7004d8728bc7356f30926[5]  <= 1'b0;
            I36b5867a3da6f2ed529e791166640d3f[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I651d700a00d7004d8728bc7356f30926[6]  <= 1'b0;
            I36b5867a3da6f2ed529e791166640d3f[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I651d700a00d7004d8728bc7356f30926[7]  <= 1'b0;
            I36b5867a3da6f2ed529e791166640d3f[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I651d700a00d7004d8728bc7356f30926[8]  <= 1'b0;
            I578efe5c2c504f12c8f2466a7f734215                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Iedc20522d3322bbe3f55e2aa611d76df[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6f5c991e5fdcf56d582c6f80eb6731df[0]  <= 1'b0;
            Iedc20522d3322bbe3f55e2aa611d76df[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6f5c991e5fdcf56d582c6f80eb6731df[1]  <= 1'b0;
            Iedc20522d3322bbe3f55e2aa611d76df[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6f5c991e5fdcf56d582c6f80eb6731df[2]  <= 1'b0;
            Iedc20522d3322bbe3f55e2aa611d76df[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6f5c991e5fdcf56d582c6f80eb6731df[3]  <= 1'b0;
            Iedc20522d3322bbe3f55e2aa611d76df[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6f5c991e5fdcf56d582c6f80eb6731df[4]  <= 1'b0;
            Iedc20522d3322bbe3f55e2aa611d76df[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6f5c991e5fdcf56d582c6f80eb6731df[5]  <= 1'b0;
            Iedc20522d3322bbe3f55e2aa611d76df[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6f5c991e5fdcf56d582c6f80eb6731df[6]  <= 1'b0;
            Iedc20522d3322bbe3f55e2aa611d76df[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6f5c991e5fdcf56d582c6f80eb6731df[7]  <= 1'b0;
            Iedc20522d3322bbe3f55e2aa611d76df[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6f5c991e5fdcf56d582c6f80eb6731df[8]  <= 1'b0;
            Iedc20522d3322bbe3f55e2aa611d76df[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6f5c991e5fdcf56d582c6f80eb6731df[9]  <= 1'b0;
            Iedc20522d3322bbe3f55e2aa611d76df[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6f5c991e5fdcf56d582c6f80eb6731df[10]  <= 1'b0;
            Iedc20522d3322bbe3f55e2aa611d76df[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6f5c991e5fdcf56d582c6f80eb6731df[11]  <= 1'b0;
            Iedc20522d3322bbe3f55e2aa611d76df[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6f5c991e5fdcf56d582c6f80eb6731df[12]  <= 1'b0;
            Iedc20522d3322bbe3f55e2aa611d76df[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6f5c991e5fdcf56d582c6f80eb6731df[13]  <= 1'b0;
            Iedc20522d3322bbe3f55e2aa611d76df[14]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6f5c991e5fdcf56d582c6f80eb6731df[14]  <= 1'b0;
            Iedc20522d3322bbe3f55e2aa611d76df[15]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6f5c991e5fdcf56d582c6f80eb6731df[15]  <= 1'b0;
            Ida86d05f907d23ff9fed06927c2ec9d9                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I6821e897aea31f7c237ca1a553bf0cd1[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia5cc3055ba3365e64cf59c4d4fd3f093[0]  <= 1'b0;
            I6821e897aea31f7c237ca1a553bf0cd1[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia5cc3055ba3365e64cf59c4d4fd3f093[1]  <= 1'b0;
            I6821e897aea31f7c237ca1a553bf0cd1[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia5cc3055ba3365e64cf59c4d4fd3f093[2]  <= 1'b0;
            I6821e897aea31f7c237ca1a553bf0cd1[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia5cc3055ba3365e64cf59c4d4fd3f093[3]  <= 1'b0;
            I6821e897aea31f7c237ca1a553bf0cd1[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia5cc3055ba3365e64cf59c4d4fd3f093[4]  <= 1'b0;
            I6821e897aea31f7c237ca1a553bf0cd1[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia5cc3055ba3365e64cf59c4d4fd3f093[5]  <= 1'b0;
            I6821e897aea31f7c237ca1a553bf0cd1[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia5cc3055ba3365e64cf59c4d4fd3f093[6]  <= 1'b0;
            I6821e897aea31f7c237ca1a553bf0cd1[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia5cc3055ba3365e64cf59c4d4fd3f093[7]  <= 1'b0;
            I6821e897aea31f7c237ca1a553bf0cd1[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia5cc3055ba3365e64cf59c4d4fd3f093[8]  <= 1'b0;
            I6821e897aea31f7c237ca1a553bf0cd1[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia5cc3055ba3365e64cf59c4d4fd3f093[9]  <= 1'b0;
            I6821e897aea31f7c237ca1a553bf0cd1[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia5cc3055ba3365e64cf59c4d4fd3f093[10]  <= 1'b0;
            I6821e897aea31f7c237ca1a553bf0cd1[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia5cc3055ba3365e64cf59c4d4fd3f093[11]  <= 1'b0;
            I6821e897aea31f7c237ca1a553bf0cd1[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia5cc3055ba3365e64cf59c4d4fd3f093[12]  <= 1'b0;
            I6821e897aea31f7c237ca1a553bf0cd1[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia5cc3055ba3365e64cf59c4d4fd3f093[13]  <= 1'b0;
            I6821e897aea31f7c237ca1a553bf0cd1[14]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia5cc3055ba3365e64cf59c4d4fd3f093[14]  <= 1'b0;
            I6821e897aea31f7c237ca1a553bf0cd1[15]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia5cc3055ba3365e64cf59c4d4fd3f093[15]  <= 1'b0;
            I9d9f8c7a23d9750ec44e706bf763df76                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I290499340d94dd8e234f53f9962a182b[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iea7da1f43ba202d753b0edb0be8b3fcf[0]  <= 1'b0;
            I290499340d94dd8e234f53f9962a182b[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iea7da1f43ba202d753b0edb0be8b3fcf[1]  <= 1'b0;
            I290499340d94dd8e234f53f9962a182b[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iea7da1f43ba202d753b0edb0be8b3fcf[2]  <= 1'b0;
            I290499340d94dd8e234f53f9962a182b[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iea7da1f43ba202d753b0edb0be8b3fcf[3]  <= 1'b0;
            I290499340d94dd8e234f53f9962a182b[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iea7da1f43ba202d753b0edb0be8b3fcf[4]  <= 1'b0;
            I290499340d94dd8e234f53f9962a182b[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iea7da1f43ba202d753b0edb0be8b3fcf[5]  <= 1'b0;
            I290499340d94dd8e234f53f9962a182b[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iea7da1f43ba202d753b0edb0be8b3fcf[6]  <= 1'b0;
            I290499340d94dd8e234f53f9962a182b[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iea7da1f43ba202d753b0edb0be8b3fcf[7]  <= 1'b0;
            I290499340d94dd8e234f53f9962a182b[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iea7da1f43ba202d753b0edb0be8b3fcf[8]  <= 1'b0;
            I290499340d94dd8e234f53f9962a182b[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iea7da1f43ba202d753b0edb0be8b3fcf[9]  <= 1'b0;
            I290499340d94dd8e234f53f9962a182b[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iea7da1f43ba202d753b0edb0be8b3fcf[10]  <= 1'b0;
            I290499340d94dd8e234f53f9962a182b[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iea7da1f43ba202d753b0edb0be8b3fcf[11]  <= 1'b0;
            I290499340d94dd8e234f53f9962a182b[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iea7da1f43ba202d753b0edb0be8b3fcf[12]  <= 1'b0;
            I290499340d94dd8e234f53f9962a182b[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iea7da1f43ba202d753b0edb0be8b3fcf[13]  <= 1'b0;
            I290499340d94dd8e234f53f9962a182b[14]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iea7da1f43ba202d753b0edb0be8b3fcf[14]  <= 1'b0;
            I290499340d94dd8e234f53f9962a182b[15]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iea7da1f43ba202d753b0edb0be8b3fcf[15]  <= 1'b0;
            I0b41b002a32b8e9e2fe68e819f228fb7                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I5ce387684404cf922955e4af33ed2367[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I872f61d20baf011e867b44dc5539fc37[0]  <= 1'b0;
            I5ce387684404cf922955e4af33ed2367[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I872f61d20baf011e867b44dc5539fc37[1]  <= 1'b0;
            I5ce387684404cf922955e4af33ed2367[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I872f61d20baf011e867b44dc5539fc37[2]  <= 1'b0;
            I5ce387684404cf922955e4af33ed2367[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I872f61d20baf011e867b44dc5539fc37[3]  <= 1'b0;
            I5ce387684404cf922955e4af33ed2367[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I872f61d20baf011e867b44dc5539fc37[4]  <= 1'b0;
            I5ce387684404cf922955e4af33ed2367[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I872f61d20baf011e867b44dc5539fc37[5]  <= 1'b0;
            I5ce387684404cf922955e4af33ed2367[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I872f61d20baf011e867b44dc5539fc37[6]  <= 1'b0;
            I5ce387684404cf922955e4af33ed2367[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I872f61d20baf011e867b44dc5539fc37[7]  <= 1'b0;
            I5ce387684404cf922955e4af33ed2367[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I872f61d20baf011e867b44dc5539fc37[8]  <= 1'b0;
            I5ce387684404cf922955e4af33ed2367[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I872f61d20baf011e867b44dc5539fc37[9]  <= 1'b0;
            I5ce387684404cf922955e4af33ed2367[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I872f61d20baf011e867b44dc5539fc37[10]  <= 1'b0;
            I5ce387684404cf922955e4af33ed2367[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I872f61d20baf011e867b44dc5539fc37[11]  <= 1'b0;
            I5ce387684404cf922955e4af33ed2367[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I872f61d20baf011e867b44dc5539fc37[12]  <= 1'b0;
            I5ce387684404cf922955e4af33ed2367[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I872f61d20baf011e867b44dc5539fc37[13]  <= 1'b0;
            I5ce387684404cf922955e4af33ed2367[14]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I872f61d20baf011e867b44dc5539fc37[14]  <= 1'b0;
            I5ce387684404cf922955e4af33ed2367[15]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I872f61d20baf011e867b44dc5539fc37[15]  <= 1'b0;
            I0e872d4c07169cac84549178fa144274                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I1ae87f851f8bd64e6e1428a143e82151[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ieb244944e7ee8236a207924f56fbc689[0]  <= 1'b0;
            I1ae87f851f8bd64e6e1428a143e82151[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ieb244944e7ee8236a207924f56fbc689[1]  <= 1'b0;
            I1ae87f851f8bd64e6e1428a143e82151[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ieb244944e7ee8236a207924f56fbc689[2]  <= 1'b0;
            I1ae87f851f8bd64e6e1428a143e82151[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ieb244944e7ee8236a207924f56fbc689[3]  <= 1'b0;
            I1ae87f851f8bd64e6e1428a143e82151[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ieb244944e7ee8236a207924f56fbc689[4]  <= 1'b0;
            I1ae87f851f8bd64e6e1428a143e82151[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ieb244944e7ee8236a207924f56fbc689[5]  <= 1'b0;
            I1ae87f851f8bd64e6e1428a143e82151[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ieb244944e7ee8236a207924f56fbc689[6]  <= 1'b0;
            I1ae87f851f8bd64e6e1428a143e82151[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ieb244944e7ee8236a207924f56fbc689[7]  <= 1'b0;
            I1ae87f851f8bd64e6e1428a143e82151[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ieb244944e7ee8236a207924f56fbc689[8]  <= 1'b0;
            I6f4ef0f404ae046519b8436171d51e09                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I646767a2d4b3029ed7acb73a15af1682[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie9b2be4c32334220e134e041ca8dfc06[0]  <= 1'b0;
            I646767a2d4b3029ed7acb73a15af1682[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie9b2be4c32334220e134e041ca8dfc06[1]  <= 1'b0;
            I646767a2d4b3029ed7acb73a15af1682[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie9b2be4c32334220e134e041ca8dfc06[2]  <= 1'b0;
            I646767a2d4b3029ed7acb73a15af1682[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie9b2be4c32334220e134e041ca8dfc06[3]  <= 1'b0;
            I646767a2d4b3029ed7acb73a15af1682[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie9b2be4c32334220e134e041ca8dfc06[4]  <= 1'b0;
            I646767a2d4b3029ed7acb73a15af1682[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie9b2be4c32334220e134e041ca8dfc06[5]  <= 1'b0;
            I646767a2d4b3029ed7acb73a15af1682[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie9b2be4c32334220e134e041ca8dfc06[6]  <= 1'b0;
            I646767a2d4b3029ed7acb73a15af1682[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie9b2be4c32334220e134e041ca8dfc06[7]  <= 1'b0;
            I646767a2d4b3029ed7acb73a15af1682[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie9b2be4c32334220e134e041ca8dfc06[8]  <= 1'b0;
            I4d04e66ad9103a685fbe088b74517452                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I48001f5c6554999a2178308ae271b70e[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id6f07dee3e47f39e3b43329c26f690f7[0]  <= 1'b0;
            I48001f5c6554999a2178308ae271b70e[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id6f07dee3e47f39e3b43329c26f690f7[1]  <= 1'b0;
            I48001f5c6554999a2178308ae271b70e[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id6f07dee3e47f39e3b43329c26f690f7[2]  <= 1'b0;
            I48001f5c6554999a2178308ae271b70e[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id6f07dee3e47f39e3b43329c26f690f7[3]  <= 1'b0;
            I48001f5c6554999a2178308ae271b70e[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id6f07dee3e47f39e3b43329c26f690f7[4]  <= 1'b0;
            I48001f5c6554999a2178308ae271b70e[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id6f07dee3e47f39e3b43329c26f690f7[5]  <= 1'b0;
            I48001f5c6554999a2178308ae271b70e[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id6f07dee3e47f39e3b43329c26f690f7[6]  <= 1'b0;
            I48001f5c6554999a2178308ae271b70e[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id6f07dee3e47f39e3b43329c26f690f7[7]  <= 1'b0;
            I48001f5c6554999a2178308ae271b70e[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id6f07dee3e47f39e3b43329c26f690f7[8]  <= 1'b0;
            I988e525020c1e43d238fad41dab4e6ea                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I7fe6d853fc1c11142b64ff8f40783246[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic7f04c065f8ff82c2288f1de77d37189[0]  <= 1'b0;
            I7fe6d853fc1c11142b64ff8f40783246[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic7f04c065f8ff82c2288f1de77d37189[1]  <= 1'b0;
            I7fe6d853fc1c11142b64ff8f40783246[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic7f04c065f8ff82c2288f1de77d37189[2]  <= 1'b0;
            I7fe6d853fc1c11142b64ff8f40783246[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic7f04c065f8ff82c2288f1de77d37189[3]  <= 1'b0;
            I7fe6d853fc1c11142b64ff8f40783246[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic7f04c065f8ff82c2288f1de77d37189[4]  <= 1'b0;
            I7fe6d853fc1c11142b64ff8f40783246[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic7f04c065f8ff82c2288f1de77d37189[5]  <= 1'b0;
            I7fe6d853fc1c11142b64ff8f40783246[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic7f04c065f8ff82c2288f1de77d37189[6]  <= 1'b0;
            I7fe6d853fc1c11142b64ff8f40783246[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic7f04c065f8ff82c2288f1de77d37189[7]  <= 1'b0;
            I7fe6d853fc1c11142b64ff8f40783246[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic7f04c065f8ff82c2288f1de77d37189[8]  <= 1'b0;
            I90d92887cb2526a2956d5e8c9fad760c                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Iadc98deb917f599574e99a90e3230e88[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4267622319ca65909a3b40484dc74d3a[0]  <= 1'b0;
            Iadc98deb917f599574e99a90e3230e88[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4267622319ca65909a3b40484dc74d3a[1]  <= 1'b0;
            Iadc98deb917f599574e99a90e3230e88[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4267622319ca65909a3b40484dc74d3a[2]  <= 1'b0;
            Iadc98deb917f599574e99a90e3230e88[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4267622319ca65909a3b40484dc74d3a[3]  <= 1'b0;
            Iadc98deb917f599574e99a90e3230e88[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4267622319ca65909a3b40484dc74d3a[4]  <= 1'b0;
            Iadc98deb917f599574e99a90e3230e88[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4267622319ca65909a3b40484dc74d3a[5]  <= 1'b0;
            Iadc98deb917f599574e99a90e3230e88[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4267622319ca65909a3b40484dc74d3a[6]  <= 1'b0;
            Iadc98deb917f599574e99a90e3230e88[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4267622319ca65909a3b40484dc74d3a[7]  <= 1'b0;
            Iadc98deb917f599574e99a90e3230e88[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4267622319ca65909a3b40484dc74d3a[8]  <= 1'b0;
            Iadc98deb917f599574e99a90e3230e88[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4267622319ca65909a3b40484dc74d3a[9]  <= 1'b0;
            Iadc98deb917f599574e99a90e3230e88[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4267622319ca65909a3b40484dc74d3a[10]  <= 1'b0;
            Iadc98deb917f599574e99a90e3230e88[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4267622319ca65909a3b40484dc74d3a[11]  <= 1'b0;
            I00fe3792cde1eeab36e576fd6634c4fa                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I3d79461a85cd6a58bf9f96f6e0d704ac[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iedd7d4ea8d082b40244c04946dfb14a0[0]  <= 1'b0;
            I3d79461a85cd6a58bf9f96f6e0d704ac[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iedd7d4ea8d082b40244c04946dfb14a0[1]  <= 1'b0;
            I3d79461a85cd6a58bf9f96f6e0d704ac[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iedd7d4ea8d082b40244c04946dfb14a0[2]  <= 1'b0;
            I3d79461a85cd6a58bf9f96f6e0d704ac[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iedd7d4ea8d082b40244c04946dfb14a0[3]  <= 1'b0;
            I3d79461a85cd6a58bf9f96f6e0d704ac[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iedd7d4ea8d082b40244c04946dfb14a0[4]  <= 1'b0;
            I3d79461a85cd6a58bf9f96f6e0d704ac[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iedd7d4ea8d082b40244c04946dfb14a0[5]  <= 1'b0;
            I3d79461a85cd6a58bf9f96f6e0d704ac[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iedd7d4ea8d082b40244c04946dfb14a0[6]  <= 1'b0;
            I3d79461a85cd6a58bf9f96f6e0d704ac[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iedd7d4ea8d082b40244c04946dfb14a0[7]  <= 1'b0;
            I3d79461a85cd6a58bf9f96f6e0d704ac[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iedd7d4ea8d082b40244c04946dfb14a0[8]  <= 1'b0;
            I3d79461a85cd6a58bf9f96f6e0d704ac[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iedd7d4ea8d082b40244c04946dfb14a0[9]  <= 1'b0;
            I3d79461a85cd6a58bf9f96f6e0d704ac[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iedd7d4ea8d082b40244c04946dfb14a0[10]  <= 1'b0;
            I3d79461a85cd6a58bf9f96f6e0d704ac[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iedd7d4ea8d082b40244c04946dfb14a0[11]  <= 1'b0;
            I6e586c5ac59a28b30c377e51287bf04d                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I2fcbccd884710be9c6a34f78d2ae6a18[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I56e1fe0c7a62589c123876f2b4e57a26[0]  <= 1'b0;
            I2fcbccd884710be9c6a34f78d2ae6a18[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I56e1fe0c7a62589c123876f2b4e57a26[1]  <= 1'b0;
            I2fcbccd884710be9c6a34f78d2ae6a18[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I56e1fe0c7a62589c123876f2b4e57a26[2]  <= 1'b0;
            I2fcbccd884710be9c6a34f78d2ae6a18[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I56e1fe0c7a62589c123876f2b4e57a26[3]  <= 1'b0;
            I2fcbccd884710be9c6a34f78d2ae6a18[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I56e1fe0c7a62589c123876f2b4e57a26[4]  <= 1'b0;
            I2fcbccd884710be9c6a34f78d2ae6a18[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I56e1fe0c7a62589c123876f2b4e57a26[5]  <= 1'b0;
            I2fcbccd884710be9c6a34f78d2ae6a18[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I56e1fe0c7a62589c123876f2b4e57a26[6]  <= 1'b0;
            I2fcbccd884710be9c6a34f78d2ae6a18[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I56e1fe0c7a62589c123876f2b4e57a26[7]  <= 1'b0;
            I2fcbccd884710be9c6a34f78d2ae6a18[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I56e1fe0c7a62589c123876f2b4e57a26[8]  <= 1'b0;
            I2fcbccd884710be9c6a34f78d2ae6a18[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I56e1fe0c7a62589c123876f2b4e57a26[9]  <= 1'b0;
            I2fcbccd884710be9c6a34f78d2ae6a18[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I56e1fe0c7a62589c123876f2b4e57a26[10]  <= 1'b0;
            I2fcbccd884710be9c6a34f78d2ae6a18[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I56e1fe0c7a62589c123876f2b4e57a26[11]  <= 1'b0;
            Ib5dc74106d8841d25a793010fdac599a                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I3d3df5d4d89adf508497bac8d75ef0c6[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia8a468877c9f96713c8141df9205f92a[0]  <= 1'b0;
            I3d3df5d4d89adf508497bac8d75ef0c6[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia8a468877c9f96713c8141df9205f92a[1]  <= 1'b0;
            I3d3df5d4d89adf508497bac8d75ef0c6[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia8a468877c9f96713c8141df9205f92a[2]  <= 1'b0;
            I3d3df5d4d89adf508497bac8d75ef0c6[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia8a468877c9f96713c8141df9205f92a[3]  <= 1'b0;
            I3d3df5d4d89adf508497bac8d75ef0c6[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia8a468877c9f96713c8141df9205f92a[4]  <= 1'b0;
            I3d3df5d4d89adf508497bac8d75ef0c6[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia8a468877c9f96713c8141df9205f92a[5]  <= 1'b0;
            I3d3df5d4d89adf508497bac8d75ef0c6[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia8a468877c9f96713c8141df9205f92a[6]  <= 1'b0;
            I3d3df5d4d89adf508497bac8d75ef0c6[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia8a468877c9f96713c8141df9205f92a[7]  <= 1'b0;
            I3d3df5d4d89adf508497bac8d75ef0c6[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia8a468877c9f96713c8141df9205f92a[8]  <= 1'b0;
            I3d3df5d4d89adf508497bac8d75ef0c6[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia8a468877c9f96713c8141df9205f92a[9]  <= 1'b0;
            I3d3df5d4d89adf508497bac8d75ef0c6[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia8a468877c9f96713c8141df9205f92a[10]  <= 1'b0;
            I3d3df5d4d89adf508497bac8d75ef0c6[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia8a468877c9f96713c8141df9205f92a[11]  <= 1'b0;
            I3eaf142d2734d2d0decef084dc037b50                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Iadecdac113e45cd08e095317d07766e5[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ida6059c6e0890f730536f97dfb83770b[0]  <= 1'b0;
            I2d171ad83e27a3745d204849a6f46954                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I2e4a339cb29f80caa8cbd630a0372ae8[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1993c1ed200d7cdf838d23c72a0c1c0b[0]  <= 1'b0;
            I977f1083f5e4f6f8ac38e2c5aecf1b79                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I423e8e9a9f19cf712372622e5c80c732[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I07e04e352df9aa1988ccf05d9cb2d1d7[0]  <= 1'b0;
            I9bcd673a4293e14fd20b48fa20492df7                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I5434db7480d96327d98156af57961745[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic4c0ebcc3711c9844a3aa3875483d2f7[0]  <= 1'b0;
            Icb7422ea46b22b9330c123b40fe343fe                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I20ebcbecf2c13a53be05ff26552b4e72[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I28e344560ba76bb3b76d01d8c53693a9[0]  <= 1'b0;
            Ic414cdba230d7ea73972b0eda1ec6b1b                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I7ba72e4bac9bd64d046733ce50f43769[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0600def6e6caada88ba6dedbb0d322ac[0]  <= 1'b0;
            Ie4e1e00503dba189b0f871c3c0810d76                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I6614526a756edaabd6a25e858b472d14[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iddbf50612c89b5b95a5c9efb5575cae3[0]  <= 1'b0;
            I721c43ab62b42a18c3f5228fc0a73262                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I47b2e8ee0c69e5301365a25d512b1ece[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iadc8f7f87b50bfff53d2d12d82489829[0]  <= 1'b0;
            I1f7cb03cf806b247be1cace4d75de942                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ibb72eb38996b41ce253875df0f620eb7[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I53a658b443200b9f11f1830547b5f42d[0]  <= 1'b0;
            I775cc766b069022bc00220050feee4e4                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I66944cd8c5bc22cd92a5cfcd68cee426[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I170f424df45651abe215ec74d649a9eb[0]  <= 1'b0;
            I08b78f774ed494fa7f119977bd92679e                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I8f2ff78b78e43fe7f6780f19d92ff7b8[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I3c897bfed190017a876c44fd73a7ecea[0]  <= 1'b0;
            Ic7dc7f94af108ca7c8003a2d07e1e168                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ieea0e49da41cdf0d062217a6e6591728[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iaecbbae967be2c62cacf2fa7f9801899[0]  <= 1'b0;
            Ibe1327961152cc2d26b3f19476a6e2c9                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I699c35d4b3c36c35ecaadb87c8b35d9a[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I52f867f1009f2e8d18b50a777942bde3[0]  <= 1'b0;
            I5ba97de444af4e8c9744c3b707502edc                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ie6c95c6ddde379ca7437e78c42a8245e[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I56a39a0c67b1de0a3cab6c61af3eebcf[0]  <= 1'b0;
            I3e4f1314042010b5d7384693b580da7b                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I85e05de515eb28d7172a95ba55da82a2[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I490a65b3f7b30540906262ec5e12717b[0]  <= 1'b0;
            I4a47ce6e21c1a274578397e480c184c9                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I7ed14b994ecbeae0536a721e16c88489[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib3c52fef8251d95e9abc8df0aad45d4e[0]  <= 1'b0;
            Id184731beb200ad6a53ce273b963bb3e                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Iad29b892bf50a3e83e4eb9b7c271292a[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If75725e534dcb00364d73a42769539fb[0]  <= 1'b0;
            I3317f2f6eef9a8ef1fe1ff68b47c5d03                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I35d2bc3f0efd23ded421f195b62a6a33[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9ddc427eef437ecc3ac4a2cf52aad4c3[0]  <= 1'b0;
            Ia6b9fa10c79e6f3847f89b35afb4cc59                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I4aaa94237ac5b28ce1d0db0d4e15ff81[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8999ca1f2fe9d4a30bd38fcb0daad2a4[0]  <= 1'b0;
            I91e98b804ef82eea53c5e8eccfec827f                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I137145b608dfe5138d4bdbea237743bd[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie11cf6677812bb739255b053a9c9cd56[0]  <= 1'b0;
            I5f1e0d0c6b50f70a6f5584124e095501                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I68a784efb51b172af79e3dec88d529e1[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iacc1d5a5c7811f0c9326ef80d1154fbb[0]  <= 1'b0;
            Id61fcc605b4b581f5d42024c2610c8b7                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ic3036adab4495c6a59055dd34a28b2e5[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0efdadfd49c035a49d92243391395bca[0]  <= 1'b0;
            Id64738b7668931553151dbadd5605b71                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I84a699063d2a7944f4a1b72b67ab5b4f[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie34d59bc77e06807937fe6f6860527e9[0]  <= 1'b0;
            I3bdfb451eb96d256da542864d39024df                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I63acf3ed504ad084a12a219790842b4a[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9661cb126908d8550b585e2bad383bd6[0]  <= 1'b0;
            Ia740d8ccd8230b28d078b2ea3e58d6ba                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I23a2a7fb24650eec8812d8671d92bf2b[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic0b832fbcbdb57745fefcc1ac1438808[0]  <= 1'b0;
            I574050722f82569d34bc2cfae1eedaa9                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I6f9156b7b5e13529ec0c34da34cb2b04[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I2afd96714b26f30483c3935c2a68e64f[0]  <= 1'b0;
            Ic8f7ec6ee09fb9ee2467e3cea30a44a3                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I09a4c92baceef72d764c6880fb62c1f7[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id6d4165b752630a1ce7ceb77fdcee477[0]  <= 1'b0;
            I2b77d922a74fdcef0d57debc789bd539                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I13a44a5dfbb198be64c99845122a6e97[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I59baaf1ad22721cde9064b8aad65ac76[0]  <= 1'b0;
            Ia1d8127af4944b23475bd7deac91d60e                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I2b57472e34677b9aafb852a3e421270d[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9094f4e9c5b60add3acee212118a1dfa[0]  <= 1'b0;
            I247abcede9914633c0a33fc402bf58ae                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ic96e056f2208c211122e5008d5fd8ced[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I13168bab2231ed22a3509142f990e408[0]  <= 1'b0;
            I1f413d3e081c6aea012b122fc94f73d5                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ie6b1ee6dfca427a82e4d1016585682d9[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I280145f996e5e249788cacca7caf0095[0]  <= 1'b0;
            I1b812fb764d3b48511c0d15a7efaea29                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ieb0276790e2d912809acc7f3a409ac37[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia9db6d176e9b9579a1aa5f257cd1a9f6[0]  <= 1'b0;
            I88882bd8a9f8718411564221ad85b223                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I9883bdcc250c2eb1f8e691d0f18b3cbc[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0ed43cf9eec83545457c57cfb6181d3c[0]  <= 1'b0;
            I232f24e2798488ee66003f3b8cc294c0                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I28f58fec52ea2df3fa3d8e4a2722468b[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b74f5fc705a0406ff2376cb8ac11db4[0]  <= 1'b0;
            I856284e951773518eb6c4232ea7f3d40                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ibf1bb88a30c8519cf22f684a9bc552e9[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I14f0d3ad4fec9ca492d6b36eb29a5dea[0]  <= 1'b0;
            I82cbeaf5b3e4796b2aaf33dcbd119f4f                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I9d2131bc965972708385d8d79c5b1687[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I3a25c80d9bf7655f4ce70cf29843db43[0]  <= 1'b0;
            Iaa7791bbc193412e5fe25000ceec23d6                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I65dc268c49445ceeef922f9c273df755[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I260dc9154b3a9fe38b0948e807bdb42d[0]  <= 1'b0;
            I44bdc0baed3d51ef54ce2728618ad339                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I7c0af5fba885dca550df150029e9ee36[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic49b2c150e2face8c362e33f2d87f9c4[0]  <= 1'b0;
            Ib6bc7e75ce750a26113cbb8895c2f024                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            If26299fbf3d11a469aa2bc573760fed0[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I714350b3b56a3249aad06d5f59fbb291[0]  <= 1'b0;
            Ib4188380f7e96d5afb99f5045674193d                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I2ba80daf0c2b625370644ab47cef63e9[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia318eb500b8bd71048bde375c1db65a6[0]  <= 1'b0;
            I5bba219c5024301e420e9a5acbdc5845                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I0911e01c831a9e46568122fa6dab2357[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia2c4192b1e4f180402550aebcf1dcd1f[0]  <= 1'b0;
            I1bb52988c9ba03e16b1b69335d3d7e7c                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ic8f0aa27dadc689b1bfb5b284fc13562[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1686a95674ecad0c4e234b8aa6e22dd9[0]  <= 1'b0;
            I1b9990aaeae716f66b0f89fb02be0a74                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I5ad4c6aba210a8b2d343ab17b49c38a3[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5ee21680396395f8338477fa2bb314ec[0]  <= 1'b0;
            Iceec2cf6aba9138648a3340390f39fe9                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I34947a54412d287f3ff730332211dc5a[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I005e89f0a9a9a52aec92752813a70f81[0]  <= 1'b0;
            Iad7842f3d4672f42c1064c28d4c8ec4e                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ia6ac380b9be591fb53c0f36f4d417a7e[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0daca3ad02a67285295cd9fc330d8027[0]  <= 1'b0;
            Ie5a53cf9343fdcdb5788667c45fadc83                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ia5d5342af30d46f66f0e4f41e5170b87[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0d2ddde9edfef483482e6c177a084f6e[0]  <= 1'b0;
            I30e06d190906bc9eb6f1c3156c47f9f1                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ica011579f46e949eda7f8eed2e4d3ada[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I932ad562b582e2c9795f241c82901188[0]  <= 1'b0;
            Ieaaaced47e22029ad2945eac9cc45e6c                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I88b214aeebaffa768ccf7c70423fb0c3[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifee4aa12e36833c935c54ef27b1917da[0]  <= 1'b0;
            I08dc6f8e837b1f6b80bd3fc742290dab                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            If46340645f788fdde3bb8f4d176aae52[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I51e5b79f738795719ac21c6a88711a01[0]  <= 1'b0;
            I8eb6a9c907c5909dad6cda98022d70b8                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ib59f285283d8c3013c20aad73ed9d148[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4e41e628a8af629421544cb4c6f45265[0]  <= 1'b0;
            Ia5067b1b458af82c3c2cd50653099854                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I3229ea9a0c348b17fcaedf6565d6d7cc[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9b2ec7db66661f7c9d85cfb1bc41893b[0]  <= 1'b0;
            I198c6753cf12d423c709d1512e66fa9b                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I3ba17818aa7ea9bbfcebb2a5f405fec1[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0a594a36728c7ac6244c504b8ea9c9af[0]  <= 1'b0;
            Ib600dd8a39fda48d28e1289d44d49a84                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I2ad1769ceb4cf0013f7b032c6e583745[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibd943ebf64fe56a1818d2bb8b9f9f8bd[0]  <= 1'b0;
            Iabf09191227584c76d7fbc634b706d12                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ib35d4bfa08a9364f7f6c8be7feaf15ba[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8c3ba90c84f9375001e727b711dead8d[0]  <= 1'b0;
            I4869ba08cab90a6dcbc454b0001a7a20                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I216edc2024d31f612d05617f6696c6c5[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I387ca23d0e2183522ab041ec48bffef4[0]  <= 1'b0;
            If97974406672507f8c9a1c507c4b6951                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I2be51c29373fe2ddfe456265a54bcc08[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib933575f5224d414f87bc71fa7498534[0]  <= 1'b0;
            I4210341f99ac7cb08245137999739114                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ib3561cb8090e7787ad8c324db3a5456a[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibfe1bddf32fa63ea87c68de7a3af1815[0]  <= 1'b0;
            Ic24f4dbd99c8f4d88c8450d4fef762b8                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I5d701e34c6fea83dccbac286a36fcbbc[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I719c50f9bbc66decebe794fe6ea017dd[0]  <= 1'b0;
            I68dffa1a13eb6ab54615347729c1d6af                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ie479179aee4de4208dda8af63ed9fb66[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I833b0433a33dac70cb215bc8cc9f4863[0]  <= 1'b0;
            I10153d5548b184b9ac2cecdba4ec4b1a                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I0acbd9a7ed1409c7958d6c630a7f96d7[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9769761eb863e3273f9253ace4c69585[0]  <= 1'b0;
            I104b7f0512440cffc0fcce25e477f537                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I390dbe9907497b62162445c90f2f27fc[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1fc63f388d047207a9375842c85e87f7[0]  <= 1'b0;
            I18b6758319272eebbe76e1eee5ae55b2                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I01d386885d97d770ff2ab01da72631a0[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I414c4d389ecc00197f2138eff0b6454e[0]  <= 1'b0;
            I780263b10b98f9bb0eaf66c045d8d37c                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Iedbfdad739e796202d764f909e6ac6b2[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibe387e8fe6f35588e028ba29cda5b912[0]  <= 1'b0;
            I37b772442e55cbcd44ba892a0608d662                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I41ded014d071bd714d053a8aed21cf5a[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I98191a7e6c56aae1b56e3d623004ed75[0]  <= 1'b0;
            I0ac256a6659ff5c6673fd110a8bf578f                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I1f14df209c8c73fe390873ae05063afe[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icd0f5c370462670cd18d30dfc0c81c02[0]  <= 1'b0;
            If134e1d27e736005e5a390e7a2ea1f4b                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I510a362375a9b9c75436ad01388de6db[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I15c59dc8eba10ff8eadfa6078678773b[0]  <= 1'b0;
            I7b37b8f908cd82683832536e02faab0d                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ic2f0b44a83961b8b49f4637ec6750f27[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I3870d672343c002ad9c83c816fd40567[0]  <= 1'b0;
            I08b4bf60c9c7e7229bd1952cc88bc7b3                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Id5cbccb1a2ccacf28b64ece8eec0099e[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic341b9d947f2d3ac57aa41f408214434[0]  <= 1'b0;
            I267d637eb63fef9f4723f7978fad88f0                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I9686b2d0e5248bfb6d3ef9b7c687ed05[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ied40f6b7847158bd08cbd932254dd6ba[0]  <= 1'b0;
            I4fb56a70e5ffa71f58f715da36368e04                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ibe5129eb30f626925a3ab5ed5e239bb3[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6ab04d323306b7290cc89ed66dbd93bf[0]  <= 1'b0;
            I5e9e2acb258baf96ac4b525bba54a462                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I2a656dad40cec86a53e732e78f00c269[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iac4a5fdede87b021e6a8150d3bf34b66[0]  <= 1'b0;
            Ic40f61443a4d8f87769067fc39381cb3                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            If06132c6a0060efdbd695b31c338faf6[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id92b1676e19c5818fa813d06dc9a01f3[0]  <= 1'b0;
            Ieb36710c9a3726f33407436d62639c8d                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I02fd20ab9e4fa12009b63fbe41d647fb[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I93da1192f27c33e21e03b9a2748774ea[0]  <= 1'b0;
            Ic804af393da2e4b9c8ef25d4a3b4e8d5                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ibb97d541a2ed2b0cbad273a09fef5594[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I69a0c79d41af6b6340430b8b337fb0ca[0]  <= 1'b0;
            I52e4c446693c29a42bb3b665f72d382d                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I0905c7e3678f66095194058bb72d22fe[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibd47f48d306ec44d94865a0a81e4f9dc[0]  <= 1'b0;
            Idbf02cf10add496d30fa44bbb18458c6                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I81433ae67b7cb4dee0b2091f3819ea88[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia5707d1275138a5145b2a42190d95183[0]  <= 1'b0;
            Ida095585ad26e215f1c1bf989912da89                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ia6249382442d1dd3062acc63f891465b[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I33bc2f42d997a2963b063326eb210d1c[0]  <= 1'b0;
            I19f1ffa05c7c9a0df5e7014044024c7b                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ie4bd4c14051455f00efdb023c3b58173[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib22e39b701614cd9986061c32adfbc66[0]  <= 1'b0;
            I4d68a2fe778fa93faac38b138138291f                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ie64e67a2316af18c5835c3a32ae9290f[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9b08176fde1cd08c9d7686a659213580[0]  <= 1'b0;
            I54393ada6f76ac82c31f2668e228e29d                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Icaf94b3fea3e29ff77d4793b389c9d14[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1b4e65357a818998d08b83d21584e18c[0]  <= 1'b0;
            If5b9ef84f09680f3593250b13a852c1c                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I334991f6bfe06389e35b7a580982de1f[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibb865ea5891db706b7b54e5c6fa383d0[0]  <= 1'b0;
            Ibb759bc4179e5b7aa759d850c7cfa467                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I6390495458553670944cdbf57bd6ce7b[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I32d42cfd2d516af2e68fc2db4d5dce03[0]  <= 1'b0;
            I05e8b5f8b83f07b609b5ebf272bb2229                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ibafc73f0a3486943914e197a7af4505c[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4d0e8d475a5d2a7da24daca60f23f3d6[0]  <= 1'b0;
            If6ac15373ec1146d38e7aeb71c3ece64                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I2ec83b82756dda6035ddff10dd41fed5[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie3850345b207e59aaaa5c944dab40b90[0]  <= 1'b0;
            I2ab3675e1eede757af80716ba980a4e6                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I5f6abb1000e5416dd4d43fcd052321fb[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4a9a1c932db30dcf04cb105a8d7384f9[0]  <= 1'b0;
            I388c271687ab31b57421ad57192273ed                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Icc865d7264dd89944317be21610dcf9d[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0ef689822226332f5feaf79fcf8f6674[0]  <= 1'b0;
            I6121679cec8caa51dc5ff0d1a61f9821                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I6a301412ef9235f3a609baf10a4200dd[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib5744c2130bb5a9d0ccdd975fdf2ff9c[0]  <= 1'b0;
            Ia0649b990bf5716cfab230127cd5d47f                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I9840f42586460341bb39256726d39ca1[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I039a7ddcb25972501d80c45c938cf683[0]  <= 1'b0;
            I867a0626ca22108b16267d95c0aadf4f                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I0837554bfb175a9ac8a4cb17e091fa9e[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic5f36c15ebad061dfbd5301e02ce2ffe[0]  <= 1'b0;
            I1af54bcb73d7c6b93e55450871207976                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Iacd698956b9ea6f1649063ee612c7e76[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Idf0d9dac06522293f8d7e00a93b6bbb5[0]  <= 1'b0;
            I91883553543d0425e9c6dd726dce3d27                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I68928b2759202e358f75b08e162e6a68[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id557db735a70dbb14504bc3088e8798e[0]  <= 1'b0;
            Ie95405659701278e3f87bf1f823a037b                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I609f881624ec9034823c9f54f4fb9b6d[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I150d31ef31093fdfc5f145d84bb35156[0]  <= 1'b0;
            Ia42392e2104b50c0908aad82738a5ee7                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I075a0a1afc1463e92edb5f7658395424[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I7e40e6f9d82d9b9fc546672e8e8621bb[0]  <= 1'b0;
            I68ad63230a51b9b9e3daffb307ea970d                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Idf1030f0e2aa5e2605bcea5fbe0428f8[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I14133cbbfa6521c5b81477fa1c229cbf[0]  <= 1'b0;
            I7a052d63944ccf42e598efe3a95b88f8                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I1b82e98260c3bdeb5183a3af470e2d4a[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I3728e31a7cf48639ce873d9135dc87fb[0]  <= 1'b0;
            I2b3c6d69f79c8d51e4d1614c62c44fcc                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I75338af3ebc7b7061a499e98a5be1674[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic6be12e390bd3c25c66d9b9e7c0532b8[0]  <= 1'b0;
            Ifcef0e92f50e3920bf1208af5d64c632                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I9f863d33f3c727e13eb52e7563ef9d1e[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icc50e1923274729fe472ca578b68c0f5[0]  <= 1'b0;
            I111340a19625901a3c1b95fd0bd1570e                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I56b8e0a7e6d2229baa9908843c0208ce[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4d98064f544a41b977ba945d2eecdf21[0]  <= 1'b0;
            I11aec4fa85c30f6fe1fd9fa72542ef6c                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I3d04bcd17aa2b98b69dcd671b9666c50[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I12f2a9f1e3e715d7e684ff39dd7942f0[0]  <= 1'b0;
            I80cc333c181c16a96b7bd6501c27c2b3                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Id254880ed38db79c53facbdc0c4a6d1a[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iaa4e3c53a0d55e8f42f60ff40893427e[0]  <= 1'b0;
            Idc6354325a6280ae9890da33c06c33ec                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I988a7c2c284c38fcd6682236dc2d6151[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I26aae317b0b320df86ca4004f64aab88[0]  <= 1'b0;
            Ibb04cf82acc4ac16599ad3ddb0c2ada2                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ida4c48caeba43eccdddd1748824ec551[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9344825cc2e5864f691043a1f94f86a4[0]  <= 1'b0;
            I3ed096dfd8a14f4acb4d53a70cf8aceb                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            If9936b476bb351a9ecbb97e2088cdd6f[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I82988c3879c1de76fe2140c469f6a4c1[0]  <= 1'b0;
            I0fa07f95e96326cb0599c0c3f76e2b48                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I6cbccfdeeb675a8a99d4c394bc8e71cd[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6bdd8334512c7c6a3226ebb4e928a270[0]  <= 1'b0;
            I87d98fbc97d9a78c2e7d6a6280e7a49a                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I79a4a9dfcecca4073c101bdd9b738c7c[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0debec6ace7160558cce7f111dd1bea6[0]  <= 1'b0;
            Ib7ddc4dca877f7cf5697a02c3d1915ba                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ice57a50f53d13e7eaf25af23547b5fb0[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8ee02e65ce9183683f0f3168bfd755c5[0]  <= 1'b0;
            I3612ef280891f6017fad205d0484bde7                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I8ff8106a70daac7c8932e88aeb6d198b[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I80e6d2c9c5f7b6bc6bffa063c4959115[0]  <= 1'b0;
            I561547649aeb5b4c3f10d9506db1f3cf                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I8f9d1ec03357f7f045196050511341a2[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0f21fb041239a7a8895c9506f2754595[0]  <= 1'b0;
            I84cc76c0079b86da7b994844c3ccb875                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ic423bfa7639075130324da59f2cca2fc[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8ce37a8e81b54043276835c11e394df5[0]  <= 1'b0;
            Iec013c508d0c6401d7eb856e7eb60446                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I4eed402353a7fa22fcb11f2adbf6be03[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Idf7d1f78735ce1e9695d99a532a7726e[0]  <= 1'b0;
            Ifd8979aac6b6b24aa560b46b18240e92                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ieb579bed6711928456b296873c5da9cd[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I96a552ed2d18c0ba3fc6cb6d6b6a0f44[0]  <= 1'b0;
            If12394e78dc913b01890b56650856a44                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ifdf316d14ef99080247091609b2c2a8f[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I3c76936e8e3467378210a13645a401d4[0]  <= 1'b0;
            I94d18aa10695f3f22b23246884b72822                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I2a1afeffe5592e35349bfd4384de834e[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic9a1d599fcfd5dd51265e5d0989719b6[0]  <= 1'b0;
            Ic90b38835dd7e760dd54067b196f8470                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I93f88eac6c04d26228b5d7a3b1d00a42[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I60156470e631268c392040d3c5582eca[0]  <= 1'b0;
            If3691ea51f6efe9b165a31964854d2fe                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I8c32ed7572af2a6a41a415ff6c580f3d[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I821126d1516ad7e8191a7b2a3b5e4b47[0]  <= 1'b0;
            Ic2ce582555add38a14f5006d3c87eb15                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I9cc4cd2860ebe1e5d43eb6024ea32dcf[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibe72e9f6d2c3cbbcf98f6b5aa6a4f93b[0]  <= 1'b0;
            I58cc950ee2cbe56b7c5a619be3792511                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I35b73e275ce37c06d10c227595c7c3f6[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1e8b6306d2dfde4a36ee9b9c2caf1c85[0]  <= 1'b0;
            I0d8e329ec5873db96df1ec309445a096                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Iac4ee00e62d47494b2bfe3aff55506ea[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I48ed92480f457fc3cc2ff0dd7d177a10[0]  <= 1'b0;
            I106325488e2ecfdba1cf9e5201e6bc8c                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I6023ec90efcd1ac53ea71eeee1c996e2[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iaed28d88a651f0151501ec4ea6ee3346[0]  <= 1'b0;
            Iff73a0085541a511d3912b64686a82c5                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I6f2b0c5e254aeb7e967f86e914876171[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9d94d9b5414662de841443d7866e66b1[0]  <= 1'b0;
            Icdab59de68f2870504598c9ea18f1d2c                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ie9353d9dd97f3536dfa6bcc2c662bf40[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I870b8a3b11be215a8704ba05568f05e2[0]  <= 1'b0;
            I75604d727e82c977741f90113719183a                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I09fd28ae4656b1282feb899a40b9b233[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia8bbf21e040b326058a9acb7d198a835[0]  <= 1'b0;
            I6f50c4d0d2639857b2dcca300c2d7b04                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Iabbb1734d7e19cd9c7329b30cb26cd3b[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie852f207c8f537621b080ffa0a89bfdc[0]  <= 1'b0;
            I5cd013a2be2e761c10c6a957632517de                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Iacc03e49c3cd6749e4c49e13c8c8593e[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If53029b05bea46d656a6ef72fb6d6642[0]  <= 1'b0;
            Iafeedddd02428bd2610c576e68d4ae25                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I7913101e04088970adf3f1e7429cd06a[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8e8a740d09e000444ba1f4931b5cccf4[0]  <= 1'b0;
            I912d6325e34180e0f668f0f024e63581                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ibddcea3450984eb0b3cc3ca6961fa646[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I46605d823e06af5485e50b256b5c3f22[0]  <= 1'b0;
            Id1e05294dfd02df499ad0c08bb5c191b                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I0a863fcba425a8683ebbb35195ea70a4[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I38344d68127f5c035193bb9030ce4d4d[0]  <= 1'b0;
            Id3bb9b100ee4302473b49ac14615e9b0                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I8138f45ab1b8a10869a2a6078b6c214c[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iba9f33c08db89a7f120cc1e3eaf05dec[0]  <= 1'b0;
            Ief32db1cfc443119b6202b0cc7bf70a2                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ie4c27f8574c8bad0b923796d2544f858[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibde51eb91b3ca50a8a0513c94bd7be15[0]  <= 1'b0;
            Iad7dbe9909b5eed3261adf92d3813acc                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ibea29d15c71d594e4e9cbe6a58ebc550[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifb94196d1653a0166567e170f06ec0db[0]  <= 1'b0;
            Ie7daf0789c35caaadbba06cafabd2b70                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I0b249349485591abcc09c4587efca78d[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9cf7557e2cac4532a77fcb212712db0f[0]  <= 1'b0;
            I2bd1f9b75d9ab94af9ddceb7528935e8                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I6bbe05bfdabac8f312c7800eca53be62[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I3159d7faeee1a904c409bde1967d2c21[0]  <= 1'b0;
            Ic3d9f5c6677758810e4865779ec303e3                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ie28e38c9881297e7ffae5c3aed4dfdd3[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I35dfb5ece5e04504d6e74739ae99c9cc[0]  <= 1'b0;
            I00af04882a25e2832d913a67d4d86d7b                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I1358b8ab0933bd596c33b622d2f9523f[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iabff939ae4acf7d7b038e028c29b6166[0]  <= 1'b0;
            Ic9db631df0a1a9108c10c3e0eca7bf15                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I46ce01ea907e88cafb7d96d22b5fffd6[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia14159444578c6dc88f2d5ea0317774b[0]  <= 1'b0;
            I749f9ed1fb2dddd40ebc28f638e02935                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I64c0e39b2f3c34d724ecf0f511a413c9[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie2306a5c441d621388b73195027fc118[0]  <= 1'b0;
            Ia45b2a24df24bd5e3c95885c8928686c                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I6ffbd03867a92aea248506af197c2e86[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I700a0fbf81e57d4970ce07090ec4f2e2[0]  <= 1'b0;
            I7427464fde340780aba7f9847b4ad564                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ie0a0c3e63be2145dc838faf227a84044[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6007914b3fb3011c3ab2f9a9d7794ab2[0]  <= 1'b0;
            I33fd1ae225e2b881b2b41e0358675e22                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I58265e8a07eede7063d5a80db2412214[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I2096f40fe62e9d6f1ff96f258ffdbe33[0]  <= 1'b0;
            I2e21a35d1cf560936fd19b944a208b6b                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I6734d5f87b795f4a05510778c22b555c[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I93d8b7a24702bacbfc528242991516a9[0]  <= 1'b0;
            I249522a3d42cc75d7a6b9ede1222ee76                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I314ced88cfc50d8b2edf129a6a3bf1a6[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If0863fae91b2ec980ebdb26cfc90ae2e[0]  <= 1'b0;
            I68b4c43d9f40ae4bfd70d2983594392c                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I8cc6f1dc58a26262f18f334b751385ea[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9ec29a319384efd562c2337e1857cb4e[0]  <= 1'b0;
            I63145e0fec15c7e7c0de105f348bfd31                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I18d34c481f17aae6b16b6d0a5aa85357[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia56ecc024eae608d7de1509d75139dc2[0]  <= 1'b0;
            I8af625de86c04016c3424d116fddab5b                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ib54b35abe1088393d275f4f45f7ed966[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iebcd65ea41cd38bfe3c8577277809acd[0]  <= 1'b0;
            I54c9c10527f83b4ee4e1e22f1e4044ed                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ie339493197828e5bd69bc49ca91aeb1d[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I75be12b14694ebcb5aff6e5d3e576315[0]  <= 1'b0;
            I972559e47c7f83bd9000ca1cfc14d8e0                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ic5084e34e9626f2e423283a87ea0d91d[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8e06fe414cd04103baf3882771a63e2c[0]  <= 1'b0;
            Ib97a7f941eb7ce2a867503a04ff86a67                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I3fee16f7ef907bcf1e2f5b2e7ec77866[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0fe8574049166c363c7cc816b1435009[0]  <= 1'b0;
            I5979b55f607c71017537f2b48b40cbea                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Iee529a0d30e79cdc9b33dd3d876a0f23[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id5f435c07240d5fe4a0e48c8f25ad0b7[0]  <= 1'b0;
            I6a56760b621f238843b091279c69897f                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I6c7373fafcfbb14c527e38e0f4440404[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1ae21e0db88f955c4f08f6d52f58974d[0]  <= 1'b0;
            Icec45bf76c241d37c9a50a5cd092da9d                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ided1b79349f8806da8f5c6898cea94bc[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I92efddd59e1ea92902a295c0b8385c68[0]  <= 1'b0;
            I2f6d3f61f2890e584d3063a09587e99b                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Id77e3ee5aded95fe141c26ad08639538[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I56948ad2b2cc245bb1003fd71ae5f899[0]  <= 1'b0;
            I7c396ea2e959d84fd9a6964617cb29c6                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I3c286283659a38021c27b5e5346b59b0[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5fb5081b7a2da89115c0080b0967974d[0]  <= 1'b0;
       end else begin
           if (start_dec || I92354deea988f3beb25bfba90735c6ac) begin
               I748f85f6680918a2e992df339b4b6558  <=
                      (Iea07d1adf9016a29cffd61d183e268d0) +
                      (If92db65b39a83e1c699e4cc6d7f9e57b) +
                      (I8f2986bc015fcc64ac5e5395ac6dd851) +
                      (I355725a804e0df68b4acf96ca98f2448) +
                      (I78212ae965ab2dcb2eed0b060d6b253f) +
                      (I0b56aa7a1b7549c91dddd3a06ecbaacf) +
                      (I71412803cc5229025487255aec62ec4f) +
                      (I32fcb28a27356bc6f403528836ea4c1f) +
                      (Iad354d876cb9fc72fc0143e6f7da9357) +
                      (If6e745bb85abba7282dae1f6f701225e) +
                      (I93bb43c1b89d4c70a57bdc019d64fd22) +
                      (I7a2e554d07bbea291f2cfc18694fca3a) +
                      (I3e59b2419c7dd1553b792d536208514e) +
                      (I46894c6526983bf1ce4b503159131b41) +
                      (I6404d0df952b5bf8292c753e4c6f35d8) +
                      (I8522c402e654d007abffcb0e904af5e6) +
                      (I5ed85845c39337c37791f16e718069b4) +
                      (I89013d61c1ea8da8b1c6071cc21c316f) +
                      (I4102100fa5f1dd299af0190862efcc42) +
                      (I4939f69abb1eac56d5021e06406a93b5) +
                      (Iadbd245bf842aebb456417579a3e6296) +
                      (Ifc8ece44a4e68c3117eda9e65f3084d2) +
                      (({q0_1[0],q0_0[0]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[0],q0_0[0]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ib0f57837099e3fdf1b908d78bcda4a43  <=
                      (I91679dfab57a372eddc7f9b94a231edb) +
                      (I2213c1a2b831f421707a261f5a58b1b1) +
                      (Ic53b875b2ddcba11406eb2ca39354757) +
                      (I634484f00590216c0f74f975c9c83400) +
                      (Ib3b1db2d8b669988c887ed780e439b26) +
                      (I735db8b0ee0ec98e4cce0030b11508da) +
                      (If1607e907e626902ee26d15020a64c21) +
                      (I081b38dbb37d4c14a6a9fd3fefa13daa) +
                      (Ibac5e7b6d4bf5cd6926358318f0c418f) +
                      (Iadfc60386481092ae85cc148a2c40abb) +
                      (Ie0ee5445c56a5f9b41640b57422206de) +
                      (Ie5f8620371236cb11c9e88c16b509ee8) +
                      (I8d7c1fe2e33bbd45379b0325a3c5e989) +
                      (I4fbdc4ee57a3be42b62d9bd43078d6ef) +
                      (I5510b88bfd65811b3200adf4ef975b48) +
                      (Ib57ef2f577cca54713c16717cbbd1ce9) +
                      (I15943aa74e9fbbaebdc0d54eb6a3bffa) +
                      (I6ac24c46319a787daa5c545de8c6eeea) +
                      (I52403a0454e5fa002e79eaab7ea497bd) +
                      (I634f0ce28934600a1a31ab0d8e59b4a9) +
                      (I7103aa739616a39c03e675ea0efb0335) +
                      (I0296d01fd3f9a269a617efd4beea9b8b) +
                      (({q0_1[1],q0_0[1]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[1],q0_0[1]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               If75e99660e3997f53f7b903bc366f47f  <=
                      (I065a81ba25962785215583e7ece27661) +
                      (I631a3300cb6685f47da7781940ec5d27) +
                      (I8bbe1a2ace8f51aa22cca5d9fc66f136) +
                      (I38c3e3e136acb79c8a0ff850bcc55f16) +
                      (I35b2c7e9cdc53a98913e1c16a3a47b37) +
                      (Ib1a2b31d49ae476e2f1fb9acba2d5af0) +
                      (Ic72f41f9bbf470aee3c9b9b8787b31c3) +
                      (I3ea4c33a9419820ed54460eb64134dff) +
                      (Ia0d940e16c8cbd4f7544f5a5cd7d83b2) +
                      (I4a8abfa0896ce414d9b98093ef84455f) +
                      (I680be647bf2a62e0ee9b5d379dc87b4f) +
                      (If4d75f83299a21802b6fbe136913489f) +
                      (Ibddfda6413e3dd2f483c3174ea836b6a) +
                      (I33bddb0adcc2af7b12a83bf843036385) +
                      (I529f92b82248efe2cf64f7da0ec8283c) +
                      (I2f34af0036985cd94ade9cc905bec065) +
                      (Ia1a0d8d7dfd6e877f15cce773f85f5b7) +
                      (I5dd29fd1a73df5662d2b636e7285bad9) +
                      (Ide530e6f4622c8a7b101b6dce9650e42) +
                      (Ibaf00a6780325882067a79f0c4d693d2) +
                      (I16e3559c63ebfed83d6698fc9a9cd93a) +
                      (I9747a02384abb1c2dd1f52b3a5a999cc) +
                      (({q0_1[2],q0_0[2]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[2],q0_0[2]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I3253481bee7dbfc0f3eac94c3252ee4e  <=
                      (Iceb7a1d4c23806b8f5824016779ad129) +
                      (I40ef50004a60ae58aedc49eb5e6797c9) +
                      (I753f92da60980736440aba814a156f1e) +
                      (I4ac79b67a8904b95f7912d24af420585) +
                      (Iad44c932cfa5c249c5e59f8c706173a8) +
                      (I10f14b6433498e3b9e9bf021b60115e8) +
                      (I96008f47b9f134c9c4274cfcfb28e550) +
                      (Id0344146d1a53d418add6d2b185377dd) +
                      (I1eede74f12d37331b399eb7136bc621f) +
                      (I3e4754acc31d99bc71525789bdee0c1a) +
                      (I11c1fc94a3bd6dffa17e1571cc6ae97c) +
                      (I5395ee57418c31e11cf847f0f514ec19) +
                      (Iff125392fa39afebae1637a19c4e23ec) +
                      (Ia6308e16fae5428f4ab6560f5b21479a) +
                      (I5ea02b5349cd4d99ccbcb6b26f0cfdd7) +
                      (I21de4f6194dec9e3c401934db92c25e7) +
                      (I57d0920119f8901bd4dea2d5f8fb5d90) +
                      (I89537301987d6da0dbe6cff3caab3ff4) +
                      (Iaf0bbbe791bb71d0f557dc71caa5fb87) +
                      (Ic7ff9cde71054c1ee9eef81eabdd7061) +
                      (I88c10c47ae424fbdcb852fbf1e94127c) +
                      (Icd2e75e47cab1d539ba9ff1b6e1d7155) +
                      (({q0_1[3],q0_0[3]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[3],q0_0[3]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ia80693da8182ee2c3708b6ec21d397d2  <=
                      (I37e6bc7aff363ed0ed1f84b23c5f3e34) +
                      (I733605337bf6972630c089d32fd7f98f) +
                      (Idcb1d8bbdeaed6768c2a418c3048e6ee) +
                      (Ia89da2f1890524ad3519ab403dd0686c) +
                      (Ie33a780b0221084898c9fc5b237b244a) +
                      (Iabbd1668e0014df518ede5216232834c) +
                      (Ibd89458312687610aa166a9538968851) +
                      (Icbaf92a8e9875bcb19a1d074779a9ea5) +
                      (I80f3c8559da8e97bc5397bb8b621a0bd) +
                      (I7a0eada108891aba06cecab5071232c9) +
                      (Ie21a2c9b22e7bf8425fb5c0f33e5f4f7) +
                      (Iaa5b2807e5cc2403c5787eeb3d10ca6b) +
                      (I6da2b3a481ee71b85f3087b36b399288) +
                      (I11094e852295755925c3c61f1df81643) +
                      (I9c633aa620cca127b0ff8cf882178e76) +
                      (I694d471fd353eb54aae08a2afa7b645a) +
                      (I816704585ad393f685731104ad3ec64f) +
                      (I85d95015a9ce27a18ccbf73bbbcdbd70) +
                      (I992e7c551b4aa818606c3465d33eb798) +
                      (I2ead0e9941e2280309ab53535b1e1ac1) +
                      (I56873feb8418005b5661c7382f2dbeec) +
                      (Ib6ea4a822da2ea32e0abf6cf8a33d295) +
                      (Id1659ccdeaea3e59eb2d3f65a65ebd05) +
                      (({q0_1[4],q0_0[4]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[4],q0_0[4]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I7fa3f2648baacebf9e4b59c179601fa6  <=
                      (Ic2171967791a0329f3e39fc19d0a6bc8) +
                      (I7d5041a6796c00188f74936d283defe6) +
                      (Iba7608ee0a01af103e022bcaf564bf6b) +
                      (Iedbe9d0e48bd36064f59faea51afddb9) +
                      (Ic3871325d57b310c95ca02fcaca529eb) +
                      (I42f9b1f8ef24ad56c10086852678b456) +
                      (I3ed5d0fca86f35b3d4b4a89c6147d0cd) +
                      (Ib0126fb335e32793c400a97c5a4a337c) +
                      (I20590d8fb97ec0b2164ffe17826136a7) +
                      (I3c128efc9f80c9b8334bf7b61de71b43) +
                      (Ic7147944f8835e26b9838fdbdc18ca41) +
                      (I698b1dbc9d8664d1c86c7a763d97b3b7) +
                      (I508bbade361787127e1a2e8687ec884c) +
                      (I2afeb2a7b199c0c6738938f156ae4274) +
                      (I86255756ddd1f88b74e070b19f8c3bfa) +
                      (I7d4924388dc5373ad7936dca76797473) +
                      (Ie317e5ea2ca4ba2060d0f491290af96f) +
                      (I56ea52c50a188ec47e48740839a031c9) +
                      (Id9b9a8fe43992ec0793845715dd2226c) +
                      (I93b69bfb228db4b569a6772179d603be) +
                      (I71afab29cdb962e1f1ca21b61dfb50c6) +
                      (I9905e2686b350e8a6e7f790563a91294) +
                      (I524e78ae6a4204e17ba4532dba047d4b) +
                      (({q0_1[5],q0_0[5]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[5],q0_0[5]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Id7699f8f89380c315303644fdebacb32  <=
                      (I71228fe4188ab1d9796081184a422094) +
                      (Ie19b39200436b0bfca13502ad36c21b9) +
                      (If6657f90c84ca5e2ba08ec705f34be03) +
                      (I60ec7459bbe99fce295406bee1f2af46) +
                      (I29ab844f80c105d247c5c15faa35863c) +
                      (I856fa68463aa5ef1ae53442699d38b33) +
                      (Ic3d00a27f15f8983a120395082854d6b) +
                      (I6b1d01c3cb8fb51e43cdb788b89816be) +
                      (Ib74a56900c1f8b159ad381f61acee801) +
                      (Ia5eba52d169755c507b9e0094e467fab) +
                      (I0899e8fec1a7209cd94757c0b2f87c9a) +
                      (I08ece7cd684e593e02321612b7a88cee) +
                      (I691c84d81c60a462e28e2b2bae3ea845) +
                      (I58dc9cce6384160c0a85c6efb3319cdb) +
                      (I56bf74b5890ec67090f499afdc0a9c88) +
                      (Ibaf2f1f8bda2f6b932dc30f8369c0e1f) +
                      (Id9364a29fd79b52d0442e18dc0227854) +
                      (Ica3a41ace27f7d94377981079952f4f7) +
                      (Ib57795a63d642a73456324bab41384b6) +
                      (Iabf572c97b48c6a7dcc19e56676e3a82) +
                      (Iefd370d0df1a93639af482f78a1e8706) +
                      (I995d2809ffaf0ecda6a004d01cb9c8c4) +
                      (I4e8ebc46bc068c3f9889d970db131112) +
                      (({q0_1[6],q0_0[6]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[6],q0_0[6]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ibf3e1ead3776901898d4b154aeb61267  <=
                      (I7b561638da1b4a45ff59be81243e4471) +
                      (If0a3b88a66a816b25f17ced5d0e8f775) +
                      (I0374ada4fe50717f2158468b7ad205d4) +
                      (I357137b41bb91e0659b1ac6ead9b5c12) +
                      (I5d70bc64cf7b3d3ef4180e082e533237) +
                      (I7d9ad929660cd212387d893266b681da) +
                      (I34be4b353cf75603301372840c2f91c2) +
                      (I14834fc8e6489775359bcecf5a37ff4d) +
                      (I633a74e4dfa841c9fd13dbb6564c8493) +
                      (I157bd468200e63385583b9045758d81e) +
                      (I918c46173eebc5b2a95e041cfd91d958) +
                      (I4f8792c18bd07b23e82bbc44b4ca947f) +
                      (I8d0a1ae4c47edf1f2b99d1175aaa7197) +
                      (I734e601f5f9d568a44a48834559e04db) +
                      (Ie421da1dc5aaea57c50d0c7d9c5a2717) +
                      (Ief5cbddfbfb98fce4812a676849b9a98) +
                      (Id113cab2dd1949d32e3c1c15273185c8) +
                      (Icfe1a689e33b2b9aa9dba692d6d610b9) +
                      (Ia4b671f3360f3ce55db0dc0e4d78ddbe) +
                      (I60cbd4369e7ba9b6532f279e5c59084c) +
                      (Ifb6c65a00d9a2c31d8b1119b949828d8) +
                      (I4a777f0dd62b19dd340ad31517c4e789) +
                      (Ib75747cb32130d44b338ed8c8af8ca11) +
                      (({q0_1[7],q0_0[7]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[7],q0_0[7]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ie486617fc1d6354c7f347692cdbd894d  <=
                      (Ic7e35cf8d5cd230b94c40714f16e2418) +
                      (Ic51bb9184dfd103703cd0c6ad6edff4b) +
                      (I103f1449c78c47396d6a54dc1c810934) +
                      (I56b3a97dc3037f0bb2eed93a9482c813) +
                      (I51e98035b35a35fdc52f5bab8f19c152) +
                      (Ia6a7f9beaceb08d81012f0e72171252f) +
                      (I21b062856ced09cb9131c01b5e166f32) +
                      (I4f1221ce7880729fe584b42ef3afe6b2) +
                      (Ie7f3f1d6cee7f02ae1b17740ed54c049) +
                      (Ib196f5bcf9152703dc32c5101076600a) +
                      (({q0_1[8],q0_0[8]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[8],q0_0[8]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I7ba403c6745e7d026282ad704e065702  <=
                      (Ide9ef5a16d8fe32353c2c2a30e8ee3b0) +
                      (Iee6f2484a381bd42e441ff072ec582e4) +
                      (I53121a39de0bcba91a4d0438be2ae958) +
                      (Iff7950f24f0a6b0073942c37fff49d37) +
                      (Ide86f019e9573706c25bd8b4552396a8) +
                      (I2370042234b0e93bb66e44b97fca3e43) +
                      (If9efe7a1c359ec03014a52870ac13aec) +
                      (I6a6eb62960b616043415406ebfc21346) +
                      (I06c7728ef64be8311f48d10d766d0c44) +
                      (I9fe11f6c8147391aa4a5afd1a4e4f731) +
                      (({q0_1[9],q0_0[9]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[9],q0_0[9]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I93cb3974b8594665b2e7ce5593fde69b  <=
                      (Id50edc56fce48130247fdbc42eeff9ea) +
                      (If3e5161254eb9056914c46263b865c10) +
                      (I58703e8b6d04f8c69ac38f5fcfdc4efc) +
                      (Ie1f41720e296ced1b74cb325b666d88f) +
                      (I5d5701435c96f1078e741921b56e3c65) +
                      (Id96e744d9b10dcddd1ae0115ea57a76a) +
                      (I0c0060fe260afa3cdc72f35ffb6938ff) +
                      (Iaec1f186cb4a65da21d41e637fc628f7) +
                      (I9c15a6a5c0db11ede80ff6d04c9a56d8) +
                      (I8922487573e02d684a3d71448c3828f5) +
                      (({q0_1[10],q0_0[10]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[10],q0_0[10]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Id6a9ab06d58c3a01e1fe04fcf61406fd  <=
                      (I47f17afcd5871fc3ac378316fd3d7ae9) +
                      (Ia9642d79bb50567348083b4435c7d66d) +
                      (I2b2bd845428c49346ef8e94e95b618f8) +
                      (Ib730fdb59198f23d1e590f6d6039e96a) +
                      (I644e83f0a7d432fba38ffb2d99088eca) +
                      (I97f2b15ce0a74e68d5a4438111adcb0a) +
                      (I84c88b631bed5311cb6e99e58941149e) +
                      (I45c5e6710240685bf54b73b0d7a64271) +
                      (I5827bc87b5db1801b7db16e1e61515db) +
                      (I1c85c8f73ef80a6808c6aec0c8eca8ab) +
                      (({q0_1[11],q0_0[11]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[11],q0_0[11]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I261bd53528b82128acabd405389c8d60  <=
                      (Id13c99b7f7500c8195b54627efbc4232) +
                      (I4636821315d702a677dc93113872e647) +
                      (I9c981b0614a29386ca5e8ebc06a17f15) +
                      (I4df3d4dac24877b14e6d361bafc1a800) +
                      (I913d818403024510c55b65b56a38dd89) +
                      (({q0_1[12],q0_0[12]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[12],q0_0[12]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               If7fa833bf1b1438e7a5bc783ee745252  <=
                      (I57015930f5b09a6c6b030ed01dad2177) +
                      (Ib54d55a70605119e37e9898b940ff636) +
                      (If7e146da4f3bd255b8457fd6902005f6) +
                      (Ied00d87af99ae55144fdde41ebfc1357) +
                      (I7774313f1ae5a2de98855aad572b3676) +
                      (({q0_1[13],q0_0[13]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[13],q0_0[13]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ibb103853fc21f8f3d466ca16557ccd3e  <=
                      (I679baea452c3c6d04c53baa88edd8eb3) +
                      (If4132b39ddb92aa02d8d0346fb0e6691) +
                      (Iba70e737d52e6812a67c159520e5192f) +
                      (Ib9ceb8315f0cd848f861bab677c2c694) +
                      (I7846bc2cc11e08d05f7c853c4920d555) +
                      (({q0_1[14],q0_0[14]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[14],q0_0[14]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I37446eb66ccfd268cb418655b8160fe1  <=
                      (I0865623d3350645e63fa6e6c9b78ac57) +
                      (I0262b30a4efa9f1cfb11d1c3940de9e7) +
                      (I7a2e79d42779ad235bca6ce3757cf588) +
                      (I09e9a3cd4c12d204f760758e873a177b) +
                      (I30b0b1d54912c1a41a02a25ab238bb54) +
                      (({q0_1[15],q0_0[15]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[15],q0_0[15]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Id17f6250f8c7f1d7f75fd27f92698da3  <=
                      (I49fb0909ddf66fc0073e6400f1a07844) +
                      (I9938397dc94002481984f5b560fadc58) +
                      (I4378d139db4b710e3587aa72df22b70d) +
                      (Ifa43d74fa91b7b9884969f575ef9ca8e) +
                      (I7c19a79f441ecbb73685db5a505e7479) +
                      (({q0_1[16],q0_0[16]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[16],q0_0[16]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I9957b02e8d0d888e6950eb553d9084d7  <=
                      (If2af8106efc1f7dd02c074af68278b3d) +
                      (I89a3f8d5f760d1a650f85814cbfdc017) +
                      (Ifae345c79662c3df3dff0fe68ad68746) +
                      (I88a61cf72347d695489909d0819332ab) +
                      (I9aaa036a6158d11c235bdc8406d79f4c) +
                      (({q0_1[17],q0_0[17]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[17],q0_0[17]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ic71258b745437bc8463fb4f847c55e27  <=
                      (Ie8df350430970b5f1229cda772440f85) +
                      (I7d77ac9b64b2e8cae21c6e36947e3ca2) +
                      (Ic1faed76fca5a9ceb7db26c2f43623d9) +
                      (I3ca2b9b77ed8d78a10aff42a07a53b07) +
                      (I1f00849ea055a7893df386aed162a7b6) +
                      (({q0_1[18],q0_0[18]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[18],q0_0[18]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I24bb5c315eacf0f4e8c86f6582389e39  <=
                      (Iaf8a19fde3de660c3fa925593bebbe0c) +
                      (Icd1da43a4d95230e79dbd35a7ae41066) +
                      (Ice9079fb6e08d629f8c0c9ce332c8f11) +
                      (I15fafe2baba4d2f28037023a81ce0a81) +
                      (If4d5b48882e9e628cf51ad2ac2f38c22) +
                      (({q0_1[19],q0_0[19]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[19],q0_0[19]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I607f203694ff76930cfee4103cb73c30  <=
                      (Id0eef1adba01447c14a6f005782dd9a2) +
                      (I1d1a7c5928982c278d068ebd262254da) +
                      (I6354a0e638340378124e4df7f3d145b8) +
                      (I0236c912c6d684bf4862b725be9d5951) +
                      (I6f3be51d69b2b64a04e55b8946d5dd56) +
                      (Icde3e6dbcf985682041f30903ad95572) +
                      (I46ee30b46020d91707689f3468f00e26) +
                      (I2605f078c1a9006c93855a9a2b0cf6b9) +
                      (I4d226dd2f0bfcdbea6a2e6a6613c1b64) +
                      (I5c942076b173cf527e1be2ddb8560e84) +
                      (Ic95191bccb18e26c10e56be395ca6b1a) +
                      (Ia284f974dd8a526f31eb81ed71a06e94) +
                      (Icc93450a007cee4c0a42717ed7600528) +
                      (I9ec9f389d0489908d497487e44c6edcd) +
                      (({q0_1[20],q0_0[20]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[20],q0_0[20]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ica8e4c56ebb37e189ca8e6b3daafdb80  <=
                      (If8a527cc7f06a9963a80a880d225d34c) +
                      (I39ff4663007dbc89b403f3b08a69bb6c) +
                      (I9590eb28a81c730b83b92ef7653e71a1) +
                      (I2ba1acca919bddcc22a41a28d43a4e3e) +
                      (I62d8efd4227cb3dc88aa08b6585fafc8) +
                      (I749e987266a20840bb8a4b1a2a2fc5b0) +
                      (I7607af5d98e8070e3d15cee23cdf877e) +
                      (I2e11a697d7f17ac30302eadb500de72d) +
                      (Ia0886ce792e062e22d0c224158cdfb7d) +
                      (I6b3cd79aa87235ff174c0299b855dd3d) +
                      (Ie4ae993ddb776bdffec843db0def2f5c) +
                      (I3ed2da9b53daac0852a06ad1acfad21b) +
                      (Idefa29d4d4e2a6e9147f84893520096f) +
                      (Id1fbbe0594dae272856566522633bb3d) +
                      (({q0_1[21],q0_0[21]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[21],q0_0[21]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I7089386c94261e0febf3b4f7dc1aec30  <=
                      (I8070a3b7d8b1a7ae90c1a2d27aed09aa) +
                      (Ie88285ce2b9c71de02ebd62e8f44ca72) +
                      (Ica1997c6c569c1d1f45224fbaa4e6b59) +
                      (Iaf08bcaaeb15bb0c971432f7f8b16d0a) +
                      (Idcb37cfc357cc088c775409fb9225b51) +
                      (Ic419255414995e7168afb97b051fa64f) +
                      (Iee6da3120d73373627b25ab7c0dedd28) +
                      (I56fc99a22960232b305d6e683c66fcc7) +
                      (I0a9a09b0ab43d2a0f1d1d01e13f0333c) +
                      (Ibc73d07e0c97a6fcae791e04106cb082) +
                      (I224bbdf94ac86c5c376d1db4f4d4e060) +
                      (I43f2b69c6b427de3095c44d4166b77cd) +
                      (I1e50c90010a3df1a8ce1cff811cc7a0c) +
                      (Ie1817cbf3a80dae435a5571dfbd2f5ad) +
                      (({q0_1[22],q0_0[22]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[22],q0_0[22]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ia1e4f20f32f7371cb0078d6e80fe8b7e  <=
                      (I0052d562fb3182890c8828e52d437b11) +
                      (I1eedecb1d8ff505c75be7787199afada) +
                      (I7ef544597a185b1de63b4ffc4a1d44c2) +
                      (Iadeedf3870f0b1eae98d0f7dbbeff04a) +
                      (I70ae07db9b44d530be220f06401d3d3d) +
                      (I7992ea31927b4f0e268462a3b0f18c5d) +
                      (Iadf927d18644a232ad1f1eba7db82934) +
                      (I2a9c673cdd7ded79e09ada38c0f47e6f) +
                      (Ia86740e870d8063f0266b68ad6d7481d) +
                      (I6627bcdbaa8afb115123777abd45435b) +
                      (I96fe3eb633eff6958ac575b997460bb9) +
                      (Iefdcb71f2903b11f5cb0b8857f7a1727) +
                      (I2eb90278aaa54b9c8212b3b4af7c3617) +
                      (I43493f70f0336453d77caf7f27503daa) +
                      (({q0_1[23],q0_0[23]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[23],q0_0[23]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I790cbca796af58b1726d0a4680cc164f  <=
                      (I26a7fe395eb583258c1ac58aaaa3234a) +
                      (I21668ff77cf75570cae97f575cbcf644) +
                      (Ie48be9e6b6fd63baa104d0a6a4561a1a) +
                      (I05370777439b01811fe7f750d2f724f4) +
                      (Icdcd83341f6b5c404f91ec7e97d0550c) +
                      (Ibba4e82d1510ddc16eb4ef64893cec02) +
                      (Ifb00ae47340bc99669c71da34cccc59e) +
                      (({q0_1[24],q0_0[24]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[24],q0_0[24]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I0a93f095f9efb1542116a295c0db9c8b  <=
                      (I75a4cf2948bebc58e12bb039ed273ff2) +
                      (I5a9fdec7d7ff99fe33ad6cd8afd9e059) +
                      (I47b1695a74e4d27389b97543415dcc67) +
                      (Ieb38fa62119a5a77c060d6634e051298) +
                      (I3459d98131faef5a5040a03847890b55) +
                      (Ie9b9221b2122087cd5f309570b6d31ca) +
                      (Id4451722e8e2393d627dcd0175dc9903) +
                      (({q0_1[25],q0_0[25]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[25],q0_0[25]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I989ba39f188a44475a83e65a4960d2af  <=
                      (Ic10356f9069e3651b9c045c906e63512) +
                      (Ic3a431f39c678b7175ed30fde1fa6424) +
                      (Ib01cfd833a63500e03333f263805db3d) +
                      (I0b7b4c0a8503c751229edfe0237cc903) +
                      (Iace01234164c8a9f7c98eeb83268745b) +
                      (Iace8b3b3a4c16763132b5aaa6b24212d) +
                      (I80a89644e278e96b1cd1c4b7f764dc34) +
                      (({q0_1[26],q0_0[26]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[26],q0_0[26]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I9bcc1d9b3dd258fa7b6042f0185d48cb  <=
                      (Ia92d2276a8a23521ad1b88df7c27bc2e) +
                      (I39bbec42c442d1e8c818f46ad9c096a8) +
                      (I88f1b5c12759a5efb2d2ded8483c9ed2) +
                      (Iaf4ae293c576af16f5f43a8b86c1aa3d) +
                      (I68b575fcbc5321d4d26a22bcdbb506f6) +
                      (Idf600b93ee1018ecf969ed7944b6bc7b) +
                      (I1cd93172cf5996bc870063aa642188a2) +
                      (({q0_1[27],q0_0[27]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[27],q0_0[27]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I9ba14715d9f33ef45681ad52f5be9593  <=
                      (I4af080cb4e5cc525db95e5f401019e8c) +
                      (I6fc8044eb226a14ff1a786ddc96d2414) +
                      (I27fd0073dbcdee599fbe85cf48806efc) +
                      (Iaee6d725a8b2653eeac6d5acb91f8f36) +
                      (I4afdeba4fc2a12a6cbe3567a519367fc) +
                      (Ib42816335dd8475dcc78662c4c0786c1) +
                      (I343c9efe71164c01e9c7d599e032864a) +
                      (I108c269ceec4adcff9afeda01101b838) +
                      (I761983331fb6e3c6c437b3f1660f0b6b) +
                      (I70d32affde22f9dcb2d77430fca39069) +
                      (Ic08e85346f61da036a15345a13ac12f0) +
                      (If5dfdadb3868ed5a495007362f7db648) +
                      (Ia1ee5579358b564de06c08ca418a9bf4) +
                      (({q0_1[28],q0_0[28]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[28],q0_0[28]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I396a897f79b519f4fa02af39d0274f64  <=
                      (I9bb81dda8102b829441be46460eb8900) +
                      (I8eef6ca0a61a21882ea28b3d63735228) +
                      (I438522d92cce6f7010246424746ca255) +
                      (I92496f68b44a94565af28a2c28d6fbae) +
                      (I66528f43f614f0edb715564eba3c77c1) +
                      (I8cab9fba615b94fd4bb6934325be8ab8) +
                      (I92d9fec22d36b1baac8bd78abfc1bbd5) +
                      (I4eadce87f47df6d8f0e4acd057de5a09) +
                      (I73203143fe37933c16fff873c1abf512) +
                      (Ibed2a63af723a7abf96dacf1951e5266) +
                      (Id667c80003b5541de9f84d3b8709c828) +
                      (I02cbb4255db2b21ea32140f9e9ddb36b) +
                      (I65354f2069de0c25bbe7cd50fbe892aa) +
                      (({q0_1[29],q0_0[29]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[29],q0_0[29]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I197c0cd576e16ee2197a28c86397f801  <=
                      (Ic279867ebf3055980f3d813d5dc8dec6) +
                      (I5c05da8a222ad5effb9815cbf3ec25f3) +
                      (Ib8bf21f32c0e8b9cfa42a53807bfe3a3) +
                      (I7208256bb198bfce1be71390b01bc028) +
                      (I49f2a06ceb3a59773c65b19f54ff362b) +
                      (I86e495dc894d2aace15c1aff89798bf7) +
                      (I0d53bb5344cabe5fa5ce3ecf7122a260) +
                      (Ib2f5f5fc77ea8b529f2471c54388f2d1) +
                      (Idcada1bfb3c0d1f2a09aab58a2071a57) +
                      (I814b62120953991f9da055f118967e05) +
                      (I123a212546a8ac394051425db4924812) +
                      (Ie95f1a7e0effcec0aa423dc803056a13) +
                      (I106deaff50b8480eac31ddbae2ec7c61) +
                      (({q0_1[30],q0_0[30]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[30],q0_0[30]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I094a178e55425f27ac1ff6195217396b  <=
                      (I68528be9951f5b8805411711cd11ea59) +
                      (I0f034a8f077b0ab231727b6298e366d8) +
                      (If9c12f8662333fb54a45cfa1bc5da487) +
                      (Ie1681d905517daafcc7584725cd6014c) +
                      (I2ff3edcdb6158f1e3c9a555aeefc0850) +
                      (I43b380be6df7df0d354223d0a0d6d6b6) +
                      (I23eb1dc4d1c992f804dd04a2d823c778) +
                      (I7f90f96c0260560ad5e6dc7448b2670a) +
                      (I07b417cdcc99eaea3413f563e26ddc73) +
                      (I2f3ab9654e515a54e22e73d6c130ccc3) +
                      (Iebdc41368d57498a04fa73e30b10a966) +
                      (I5b4305bef5b4350c1d7ae143667afddd) +
                      (I2795d21d343b83a69146314a2407cfa2) +
                      (({q0_1[31],q0_0[31]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[31],q0_0[31]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I3177408f7d08b431be99297fb10586e6  <=
                      (Ic6386d7d8813731d612e24b715740275) +
                      (I4c366a57920ff090a98a2cb8b9caa00b) +
                      (I14cf5d43fc9864820a8a25efcc5c6d86) +
                      (I33b99994abbb5ecf8eed4de39033e4f8) +
                      (I7c3291f0250d13ca94802b0b071a95c6) +
                      (I2c926fd9d306e9ae13364e07c4b0395b) +
                      (({q0_1[32],q0_0[32]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[32],q0_0[32]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Id4948c876d48bdbf317d32f135e645b4  <=
                      (Ib23edc35fa5bbfe0415fcf0861a22d9b) +
                      (I3e0e682047f7cc36142e668828cbff1e) +
                      (I99fb9030e8361e57818c07511479a9b8) +
                      (Ic87c3d7762a18772972552162e1d1a8c) +
                      (I7e393e6c1d1bc44daaab120d55f5dd59) +
                      (I448f126fd3932d5065abbe7bb2d92c56) +
                      (({q0_1[33],q0_0[33]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[33],q0_0[33]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ice5ff01d4fb4583898498651a0ac0171  <=
                      (Ifc8c6df8904b97674f2970ebc95b523c) +
                      (Icd0622a90782b9c451950e7ab0399567) +
                      (I6493b3c087d4685a6b3f98c73dc2ff49) +
                      (I20c2057240417146df144b518b43d052) +
                      (Ied029d0bdea3bf134744c99426fa72dc) +
                      (Icb82c9ff4cb58159a1c3115c6fdd5f8c) +
                      (({q0_1[34],q0_0[34]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[34],q0_0[34]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I0fb33a5ced3d15622c9aefa188052e24  <=
                      (Ia3450e134e4086c35acbdee1e6042396) +
                      (I5a0f27df5158309f32f0df31e8ae3ae3) +
                      (I17d9e19854cef197fd3267618617efc3) +
                      (I2993acb61f1abe529f8a60c94a438550) +
                      (Ic8be2c94235fb40f78da33179ce4873a) +
                      (Ib3367565e4456da15e7c2315dccdb5e4) +
                      (({q0_1[35],q0_0[35]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[35],q0_0[35]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I0074e1c3ca0ff903a9201ac5fe7ca841  <=
                      (I15a1671def323cd294591564ae6ef8b1) +
                      (Ic512effb493a06ece58a2af155135004) +
                      (I2c72248cbe49ec0a0febac2437b8a6dc) +
                      (I964e17c41a134c080e9c43412a514f3f) +
                      (I94f1724740defe5bb7e40041d0e266a0) +
                      (Ic19486b6ab0373b9c0ad8f7597782d8f) +
                      (I31243de90dc2a1656ca9d5e03bdd78da) +
                      (I242a30bdc8699d8ff550b25dd53d6c59) +
                      (({q0_1[36],q0_0[36]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[36],q0_0[36]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               If65f587e987a51c093e8dd4df532e26c  <=
                      (I9d15f76bb68b214057566cba4b511214) +
                      (I9cc16a00912e7dfc05fb505a9db23cd8) +
                      (Iacf9640cbf486411d6ceb8fe1a2fd5c9) +
                      (I9015033ab0caf3fa41dae4de43f24a82) +
                      (Ia630e59cbce82a570ae3890a6c0221e5) +
                      (I4904ab14b19fa1b6befc218bc7be3842) +
                      (I282d2eb4e74e034694e33273b9cb19d5) +
                      (I3f33901c407a87e10d86c13c83dd52eb) +
                      (({q0_1[37],q0_0[37]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[37],q0_0[37]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I33d7e77d08590f0dfb1867e741dd8b6b  <=
                      (I43f41bf07836cee48069e9890c1de2a0) +
                      (Id88480a0a350bb5fcf01ed5fff0bbd4c) +
                      (I1d9b9ff357667a362f0442f19986f451) +
                      (Ice73589836da9028def6efb24a04dbbd) +
                      (Idb72c046c5996fbbd80b706666ffbd92) +
                      (Ie5757e7b1647ab7d43cdbcf98cbb77fc) +
                      (I6072331f838d82329a07a4ffa340c7b6) +
                      (Idf6875955525d80dc660ce956f4a84e7) +
                      (({q0_1[38],q0_0[38]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[38],q0_0[38]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I678c22563e0273403b046df4261f21cf  <=
                      (Ia96955d9c0a8a587e0afab37c8415d8c) +
                      (Ifec374bce7f5507438f550df22d61a01) +
                      (Ief67e897e57b96e2ec200e82bbc7caeb) +
                      (Ide604e9bbe35cb55892a4602e18b2527) +
                      (I262f2390e77ec486ccd3a6ed05816e2d) +
                      (I280e20c20c0b4f26278b3de9b2ff84e4) +
                      (Ib3a0307176d424a4733720416d71069d) +
                      (I76060709de3ea188748849f043c59ac0) +
                      (({q0_1[39],q0_0[39]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[39],q0_0[39]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Icca700c12ae2e8155ca6b41e692e8a8c  <=
                      (I8be20605d26d218911e80a883a90d085) +
                      (Ieafa9d74d4a61d28ac4a913db460bf33) +
                      (I6fd1b4395af175eff85b3bfeef4c329b) +
                      (I39e6d3fb468aa40ea73535e81556ea65) +
                      (Iae449b74e50e0907feae9e60f2329426) +
                      (Iebf769a6bdaf214c1006c55c608d4eda) +
                      (Ia030c08757123aae947f86ab8bfb6d94) +
                      (I8c35c5b343b552c22000e194c517ca12) +
                      (Ibf80bb564263ea85bd886a8617f09bb2) +
                      (({q0_1[40],q0_0[40]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[40],q0_0[40]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I5ed74e81d2497681af5a0ca13fe23088  <=
                      (Ib8dfd9b8badef282ca00a4f793c3c868) +
                      (I596ad7e132f272cb196b74faa8c75aa4) +
                      (Idc629414f6d0236ce0714cfaae23f065) +
                      (I157fdf8775206858c08682db3039b084) +
                      (Iacbb4daf5ce5c7eb1a2afe30d0cb5382) +
                      (I4e08021c0235fafb60200aab97827a8f) +
                      (I730634ea15ac94d241f3ad2d6393a227) +
                      (Iee367c535d9c39f872d2ec043e7e7b33) +
                      (I68bb1f26f878862f288c1f57049cf58b) +
                      (({q0_1[41],q0_0[41]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[41],q0_0[41]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ic7fa6b8cdfcf7d83d4e101d9c8b7b34f  <=
                      (Ia9b5d9ede006c56a6d83905529c77b7b) +
                      (I1487170cb1f3370ad45efc801cefc8ab) +
                      (Id88568dd34fbee42c9cb8cc15ac5c31d) +
                      (Ia30539545e66c4cfc16828140149180a) +
                      (Icbfbb37bad6344005dd233b3605a784f) +
                      (I91a6408a11fab36a8ba3dbd3f895a803) +
                      (I47b878f27c30f79a37e97e022307e9e9) +
                      (Ie76b0739aec66f8860870e66e87a6445) +
                      (I50383e3d7c172eedfa00aa50a9faac4c) +
                      (({q0_1[42],q0_0[42]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[42],q0_0[42]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I26010e26e22d8a2ea831e86fae34a24e  <=
                      (Ifeaa99e03bda8ded058f98387de3d49d) +
                      (I4255ac1af4367c321567c4e46b06ab25) +
                      (Ia445bdc7def7d8c1eec31ab892c25c41) +
                      (Ic3b4752136ac08e343933ccc3a4ec47c) +
                      (Ica6707efd6d44ba6bbb87c0593a3d828) +
                      (I739267bcc50c54b8a685cb3c6afc5cc1) +
                      (I9160d11439c5140c0109b5190eb82e6b) +
                      (I6ff7b86cd7f63f9243646f1be10b2577) +
                      (I165653ab165cfafe2b74cd441331f9e1) +
                      (({q0_1[43],q0_0[43]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[43],q0_0[43]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I578efe5c2c504f12c8f2466a7f734215  <=
                      (I08a8cd6965c23af6650568b654831b20) +
                      (I9b6a674dbcbfcf65f1ae0deb8fc3566d) +
                      (Ie3a336de822ac7baf8486b1618ef1126) +
                      (I5fc3c26d6c5aa893dfd5caa0f677233a) +
                      (Ie22b94121b58f17af14c75bfb27f96dd) +
                      (I0d9f8c99194d9d6e187b4ad02fcce8b4) +
                      (I71e101962e766a4d1484b3235359a4b5) +
                      (If2539da6722562bbf31786fd0036666a) +
                      (I22c8ccd4a9018ad1c129aa058bf579d8) +
                      (I83330fef69470d2f5def8e6d7d9c50d2) +
                      (I0539d598bbe3d50940329a282c801328) +
                      (I202f88fdc946494d55fc8831c2e8a34c) +
                      (I3ee10f6a7785a236db317515fdd23a2d) +
                      (I453fdf4fbb5af5bd28a20d7643da9eb2) +
                      (Ic4a6c02880a9aead7353332708e3f388) +
                      (I7fb3b66cb48521f8715f66bf5642cdb2) +
                      (({q0_1[44],q0_0[44]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[44],q0_0[44]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ida86d05f907d23ff9fed06927c2ec9d9  <=
                      (I2fd872df07f50688486c0d602cfc5549) +
                      (Iccefa45795486757515d95e5908b306a) +
                      (Ib1357cb20f471f1670ac2448f964f8eb) +
                      (Iab953a8974a1eb619dc0f074c003b5f9) +
                      (I6e37582849c2c98fd15ad92d22c222da) +
                      (If004de0cac6e5f7701a1fce48c6936d5) +
                      (Ic1efa395cc1fd2c5a1d1559fb169a5a0) +
                      (I8e96c69e7d872be23229353808c34953) +
                      (Ib6aded6c73a8cc3cb964b0ae895b859e) +
                      (I939368b76d98b43826c68c7f468a5632) +
                      (I544f6263f16cd5e0b7cf28c511a8f6e3) +
                      (I484545c4d2c869d79eb17f51e11070a3) +
                      (I39289e6385a9bc378a9b8dd440249a7f) +
                      (Ie9cce5746a83479a567bbaeac6dbf497) +
                      (Ic044d7419cc43736d278c2df33b4a3cc) +
                      (I6714551e8885ef5e4490673fe1b2dad1) +
                      (({q0_1[45],q0_0[45]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[45],q0_0[45]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I9d9f8c7a23d9750ec44e706bf763df76  <=
                      (Ie9ab3c88ac62369e3d92d110165a94a8) +
                      (If38feb4f76f761dce6145731ad235d7f) +
                      (I6359856a1843d8c8b65dc478bccb3acd) +
                      (If6f3d91c3c7a43622b9a522492cd83d3) +
                      (Id023a6298e65da1f4da3831f5136afc2) +
                      (I6b24690f394792edb0d82b3b9e110851) +
                      (I5b55c285f7e3e78447fee68532ab9f7f) +
                      (I32701d9e4b96853c53f0ab651a6a4ba2) +
                      (I82f266e5792cdb6e7ebd264e246161f5) +
                      (Ibfacfe5b83819afe7fbd4bffa2d6d4e2) +
                      (Ib8e68a77ad8b9e7cf415bee17645c3f9) +
                      (I644ee0055a55f54ab3544bb532e39c61) +
                      (Ic5467e42aa377c6ffd8f70673808774f) +
                      (Ic57eb4a034247a4c952d8224ea9f2bac) +
                      (Ia642db613c0ec1ca4e69afde7a14a839) +
                      (I432aa7cb844286c442356954f8814260) +
                      (({q0_1[46],q0_0[46]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[46],q0_0[46]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I0b41b002a32b8e9e2fe68e819f228fb7  <=
                      (If520c1cd27f9d4bc52d0d029f693b660) +
                      (Ie87075ac979410cc11099a356966b8a2) +
                      (I6fab46b1766878b26b53f352fee98223) +
                      (Ieaf14683f40374c4531326d228cb43c3) +
                      (I5149125aaaad943d891df6a3c2be93a0) +
                      (I770dff588ee1f52f58bea1921cb23383) +
                      (I8f0a90e761111a613d2488285534a500) +
                      (I765a8825e42180a6c63f7b33703bb483) +
                      (I512cc8f6519aa08aee18225b56d47c9f) +
                      (If08370fd0e8af818c6db20f43e74034d) +
                      (I0ff382edfc8051459657ffa3899f5f73) +
                      (I9d2864024148337277523ef7fa2e1600) +
                      (I1c85a2d1df6749a194072eb731506bfe) +
                      (I3e3ce8b4ead150a6eae2e5c701c7b598) +
                      (I45bc13ae0e0554a79c62cd9c6aa8f2a5) +
                      (I92678f5b52c9c55556ff7f17f0f607b7) +
                      (({q0_1[47],q0_0[47]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[47],q0_0[47]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I0e872d4c07169cac84549178fa144274  <=
                      (Ib4bdc9069d0c08655f5e87f705943eda) +
                      (Idbf9094c94c931f16fba468b9dd59a25) +
                      (I1c3c4ce44610e04c5eef2fcbc2ea5114) +
                      (Ie84be0ae8311d906eff08f7f5b214943) +
                      (Ic90b98708faa8c8b75d4bd9a52c292f7) +
                      (I8eba6f14f42701d22859fbea94bd1871) +
                      (I6d83efa9f988328f487e9232bf2633a2) +
                      (Ic23e01562c8a753fd70c343297be288a) +
                      (I5669856f88f5e2c98f64df696db76414) +
                      (({q0_1[48],q0_0[48]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[48],q0_0[48]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I6f4ef0f404ae046519b8436171d51e09  <=
                      (Ic3a608b850709286ea0ad2f67425d9ac) +
                      (I5267fa34449e6eebe891017fc32d0749) +
                      (I599d01cfe6e54d8e45d64446c446818d) +
                      (I8f94dbafaac589ac9f14b56d4556ff96) +
                      (I754563caea429d3d0e22df5d193b84eb) +
                      (If7f373506cac70f8ba1222db135c27e8) +
                      (I69f563e7b7ad483893ac9c4684349769) +
                      (Ia0a02781c674fe5d769206448d475245) +
                      (I1b7a401bc11741e6f011fb9895b5c797) +
                      (({q0_1[49],q0_0[49]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[49],q0_0[49]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I4d04e66ad9103a685fbe088b74517452  <=
                      (Ieb528d666fdb708279184bb59eac25d9) +
                      (Ic3ff7ce12c836bf0693252b9a7a7cfe8) +
                      (I19bba6a58ad3ef959b33701f82761984) +
                      (I8acc93b34974c1e708b0e1591f7b2d3d) +
                      (Ib60d4ac0fcadcdfce5a14fb92f58423f) +
                      (I039f05d5be891a37e04556f1eae674d2) +
                      (Id0f75e19b94541ed5c5c352d13390d2d) +
                      (Ife1190f76c2e251704c2960c23330a48) +
                      (Id3e0c98bff2636e216b4d3a0ffd51054) +
                      (({q0_1[50],q0_0[50]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[50],q0_0[50]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I988e525020c1e43d238fad41dab4e6ea  <=
                      (If4d3b31b87c0f723241d35ce7e854eba) +
                      (I72369dedfe36cb22269033cc305b730c) +
                      (Iec71fe7fcebccf1ae0d10a5d187fcc44) +
                      (Ie11da10808c4ca84f399535df6261307) +
                      (I280fa9d114e227cd649bf0e55e845651) +
                      (I94c4e11670b4233fa072517a8f19c901) +
                      (I4dca2dd40a7127ce44f83b430a34c738) +
                      (I1a24e98165afa62bd14986911a36fb6e) +
                      (Ife1164cad7cda4aa9a08d94dfe86add6) +
                      (({q0_1[51],q0_0[51]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[51],q0_0[51]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I90d92887cb2526a2956d5e8c9fad760c  <=
                      (I8d8d95ff26f33f69a182b32ccde23905) +
                      (I2508854bcbab37bd09c9465c377c06aa) +
                      (I140078292f7209eccacd53a8bab18016) +
                      (I141fb1cbe09f9abe282cffd4de815d25) +
                      (If79d1d378f7c6fd29fc3335ec5f5c51d) +
                      (I4a41999cea9357a85c73a0af509eeac9) +
                      (I8e517c401d62dbb10dcc96ab536f6afb) +
                      (I8ad3627f171eadcc960a688ac0afcbc0) +
                      (I85c4d3d6c8408c6f38741257ed177ca6) +
                      (Id66c47fd69c175a4393e975a269cf053) +
                      (I37dca40506d61bdeab1255ed4892ca20) +
                      (I340c98b886123c541a1b8d9fc8a6d48c) +
                      (({q0_1[52],q0_0[52]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[52],q0_0[52]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I00fe3792cde1eeab36e576fd6634c4fa  <=
                      (I2dc64c3b06588542b027f997437bee63) +
                      (Id92a37c091100e9df08e24498ecb4022) +
                      (I74a4b9365391fd20c34588002ad40547) +
                      (I461195b7ae78743e09ee50486ad6ebe5) +
                      (I356d747600182675699a2d2634d4c5ce) +
                      (I87d6a5d30c3e4202cf51f33c7a770c51) +
                      (I960768a84aec9d5b8bc7c1c523024a25) +
                      (I09b5273bb15d48a7fd78559930fa6d1c) +
                      (I5814a85c45fd0f7be21ed325235fe4b7) +
                      (Ib06b60cf9933dd8952206c5f3ccced8e) +
                      (I67347c413b5efd8ff9e0d5bc7ab2a047) +
                      (I72b1bb104bf2843f161448baf7aab44b) +
                      (({q0_1[53],q0_0[53]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[53],q0_0[53]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I6e586c5ac59a28b30c377e51287bf04d  <=
                      (Ib23d889edb5a6d9f27de977d3b1a2616) +
                      (Ifaff9dd032cf96487be819c59b03000a) +
                      (I028ce03be0618b816e0ecdf43d4cd6e6) +
                      (I6ae2523095237282533e0b5f1c26b488) +
                      (I5aba6218461e8d571be03a3ef041ebaa) +
                      (I6ca8a1fa2c72b1c61d11dc7d1ba5f37b) +
                      (I3ec5819176ad4b0895a9118d90ab22b5) +
                      (I49b64469d298012dbb131d879bff38d6) +
                      (I95361d5f524ccb9feb42811af5c482e2) +
                      (I9c4b34b5fb1d59c132bcaeb6258675df) +
                      (I613d4b1e3b9e812b785c9cf14fefdfe6) +
                      (I848ed394bd4f0b199d11c0ff458394a7) +
                      (({q0_1[54],q0_0[54]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[54],q0_0[54]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ib5dc74106d8841d25a793010fdac599a  <=
                      (Ie65a0634454381e24bb3223a333e3ad0) +
                      (Iad166146f7df5e8068fc6efe4d3e4141) +
                      (I63e45abd4d27219bddcef06108b72021) +
                      (Id1bacd13718f7c29c26b63c239d04dd8) +
                      (Ia3104c69fb4f7abfb5efa3874169a7ad) +
                      (Ie1b7257c99831ec5864f65958ecf14fb) +
                      (I4accbad1b451ed2b622e15ef9ae16d13) +
                      (I5ce8b2f633011e89356243a1a71edeb6) +
                      (I3e5139f24e3d082eb31b0e61ea9fa1aa) +
                      (I61cc8a0f49e393721a62a776e4793deb) +
                      (Ie631e40caade823a196370fc3358f042) +
                      (I4c971e714427664c59c6371e14781bae) +
                      (({q0_1[55],q0_0[55]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[55],q0_0[55]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I3eaf142d2734d2d0decef084dc037b50  <=
                      (I36ca732e811d67cd742d24fd4cae887b) +
                      (({q0_1[56],q0_0[56]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[56],q0_0[56]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I2d171ad83e27a3745d204849a6f46954  <=
                      (I354fdd241d5d07f0d8380fe8924e0a8c) +
                      (({q0_1[57],q0_0[57]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[57],q0_0[57]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I977f1083f5e4f6f8ac38e2c5aecf1b79  <=
                      (Id38b705f5d2863a020a475ffffc8afd6) +
                      (({q0_1[58],q0_0[58]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[58],q0_0[58]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I9bcd673a4293e14fd20b48fa20492df7  <=
                      (Id6e5d67e7bb7c4b999459374ea80459a) +
                      (({q0_1[59],q0_0[59]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[59],q0_0[59]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Icb7422ea46b22b9330c123b40fe343fe  <=
                      (I05341013abd4206eb66fcddfd63bfe26) +
                      (({q0_1[60],q0_0[60]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[60],q0_0[60]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ic414cdba230d7ea73972b0eda1ec6b1b  <=
                      (I15da71a21f5842cb65b543d9bc3e267b) +
                      (({q0_1[61],q0_0[61]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[61],q0_0[61]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ie4e1e00503dba189b0f871c3c0810d76  <=
                      (Iccf255fb3422c558465e45226068a16d) +
                      (({q0_1[62],q0_0[62]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[62],q0_0[62]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I721c43ab62b42a18c3f5228fc0a73262  <=
                      (I1c2674b2e6b269ed539827412c5199a5) +
                      (({q0_1[63],q0_0[63]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[63],q0_0[63]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I1f7cb03cf806b247be1cace4d75de942  <=
                      (I6a3f405bb4a0c4448d9b9d3dd95d036c) +
                      (({q0_1[64],q0_0[64]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[64],q0_0[64]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I775cc766b069022bc00220050feee4e4  <=
                      (Ib528bb7a64cce4f694081d151fa6fa86) +
                      (({q0_1[65],q0_0[65]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[65],q0_0[65]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I08b78f774ed494fa7f119977bd92679e  <=
                      (Iaa40bd3abf668a21e0f87c7bda7b3f69) +
                      (({q0_1[66],q0_0[66]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[66],q0_0[66]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ic7dc7f94af108ca7c8003a2d07e1e168  <=
                      (I919d36a7f6ad42c4bbc23222beb73106) +
                      (({q0_1[67],q0_0[67]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[67],q0_0[67]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ibe1327961152cc2d26b3f19476a6e2c9  <=
                      (I648d2a279dd1f587b1e45eeb35f2fa90) +
                      (({q0_1[68],q0_0[68]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[68],q0_0[68]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I5ba97de444af4e8c9744c3b707502edc  <=
                      (I194a64bef92ecf6714141eaa5d41c9d4) +
                      (({q0_1[69],q0_0[69]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[69],q0_0[69]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I3e4f1314042010b5d7384693b580da7b  <=
                      (Id332e7f482524adeac7f7cdafcf5ca46) +
                      (({q0_1[70],q0_0[70]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[70],q0_0[70]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I4a47ce6e21c1a274578397e480c184c9  <=
                      (I226383d68f89db716cfd8d08b837865a) +
                      (({q0_1[71],q0_0[71]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[71],q0_0[71]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Id184731beb200ad6a53ce273b963bb3e  <=
                      (I2bdf5d319ba9089a4da34b108f5c5ae5) +
                      (({q0_1[72],q0_0[72]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[72],q0_0[72]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I3317f2f6eef9a8ef1fe1ff68b47c5d03  <=
                      (Ia91800792941ec7cc60415c3f844e4ed) +
                      (({q0_1[73],q0_0[73]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[73],q0_0[73]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ia6b9fa10c79e6f3847f89b35afb4cc59  <=
                      (Id7c507d96098ee7a955af8a48ee5d72a) +
                      (({q0_1[74],q0_0[74]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[74],q0_0[74]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I91e98b804ef82eea53c5e8eccfec827f  <=
                      (Ie15e4c1bcdb0e18085d4b320ac6a925c) +
                      (({q0_1[75],q0_0[75]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[75],q0_0[75]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I5f1e0d0c6b50f70a6f5584124e095501  <=
                      (I5485d9edcafc6202f6e5f0969979802f) +
                      (({q0_1[76],q0_0[76]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[76],q0_0[76]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Id61fcc605b4b581f5d42024c2610c8b7  <=
                      (I7fe364f9f537cbef782e7007848a1c10) +
                      (({q0_1[77],q0_0[77]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[77],q0_0[77]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Id64738b7668931553151dbadd5605b71  <=
                      (I52dcf5bace9cadcf8a895aaa6a8c1da8) +
                      (({q0_1[78],q0_0[78]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[78],q0_0[78]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I3bdfb451eb96d256da542864d39024df  <=
                      (I13a9eec6175e695ab8bc4516cf57d6ec) +
                      (({q0_1[79],q0_0[79]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[79],q0_0[79]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ia740d8ccd8230b28d078b2ea3e58d6ba  <=
                      (Iee73a7c685a4cee03f33d3ef379b1c8a) +
                      (({q0_1[80],q0_0[80]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[80],q0_0[80]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I574050722f82569d34bc2cfae1eedaa9  <=
                      (I740dc91716e3906ad078e2c7cc3c925a) +
                      (({q0_1[81],q0_0[81]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[81],q0_0[81]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ic8f7ec6ee09fb9ee2467e3cea30a44a3  <=
                      (I514d2dc697e9b39ba027c418a6df6cb9) +
                      (({q0_1[82],q0_0[82]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[82],q0_0[82]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I2b77d922a74fdcef0d57debc789bd539  <=
                      (I782726e317a2aada9e755bcbc4b0d3fa) +
                      (({q0_1[83],q0_0[83]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[83],q0_0[83]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ia1d8127af4944b23475bd7deac91d60e  <=
                      (I11eb26cf0f0b3a334e8f7317bf8d9eb0) +
                      (({q0_1[84],q0_0[84]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[84],q0_0[84]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I247abcede9914633c0a33fc402bf58ae  <=
                      (I26cb63ba20245b2c332b09e25c4409aa) +
                      (({q0_1[85],q0_0[85]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[85],q0_0[85]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I1f413d3e081c6aea012b122fc94f73d5  <=
                      (Idd7691d31f8d0c09ee988116d574ec59) +
                      (({q0_1[86],q0_0[86]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[86],q0_0[86]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I1b812fb764d3b48511c0d15a7efaea29  <=
                      (Iecc02842a2d2b9b9e8187f2d39e62e05) +
                      (({q0_1[87],q0_0[87]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[87],q0_0[87]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I88882bd8a9f8718411564221ad85b223  <=
                      (I5551342f1751fc64f32744a46b9649be) +
                      (({q0_1[88],q0_0[88]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[88],q0_0[88]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I232f24e2798488ee66003f3b8cc294c0  <=
                      (Iff7c29299f005c1cd5a16b64601e727e) +
                      (({q0_1[89],q0_0[89]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[89],q0_0[89]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I856284e951773518eb6c4232ea7f3d40  <=
                      (I17a5446e942bcc1dc2c96930e0a87a70) +
                      (({q0_1[90],q0_0[90]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[90],q0_0[90]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I82cbeaf5b3e4796b2aaf33dcbd119f4f  <=
                      (I719b67f84e07e90dfd29a8cd5d94cf39) +
                      (({q0_1[91],q0_0[91]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[91],q0_0[91]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Iaa7791bbc193412e5fe25000ceec23d6  <=
                      (I2c835dfb3596b8bf057a7cc21122c81f) +
                      (({q0_1[92],q0_0[92]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[92],q0_0[92]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I44bdc0baed3d51ef54ce2728618ad339  <=
                      (Ib71b3d357c98dcdfae5c777ca3082275) +
                      (({q0_1[93],q0_0[93]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[93],q0_0[93]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ib6bc7e75ce750a26113cbb8895c2f024  <=
                      (I086bf19f620c8a8f6888e775cb1ed7f4) +
                      (({q0_1[94],q0_0[94]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[94],q0_0[94]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ib4188380f7e96d5afb99f5045674193d  <=
                      (I802c554d5b04af6b949677819a4966ed) +
                      (({q0_1[95],q0_0[95]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[95],q0_0[95]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I5bba219c5024301e420e9a5acbdc5845  <=
                      (Iceefb06cb3715e1b41e6f7d89420e5ba) +
                      (({q0_1[96],q0_0[96]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[96],q0_0[96]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I1bb52988c9ba03e16b1b69335d3d7e7c  <=
                      (I56948bc48c0220893d68004615a6ebaa) +
                      (({q0_1[97],q0_0[97]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[97],q0_0[97]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I1b9990aaeae716f66b0f89fb02be0a74  <=
                      (Iec1368f034655d61354ab5b5e94d7d89) +
                      (({q0_1[98],q0_0[98]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[98],q0_0[98]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Iceec2cf6aba9138648a3340390f39fe9  <=
                      (I1e43c0aeeb8a2461d208eba24967af30) +
                      (({q0_1[99],q0_0[99]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[99],q0_0[99]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Iad7842f3d4672f42c1064c28d4c8ec4e  <=
                      (Ia6eb85b127cf9c1a437611556296b967) +
                      (({q0_1[100],q0_0[100]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[100],q0_0[100]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ie5a53cf9343fdcdb5788667c45fadc83  <=
                      (Ieba89aa901e61218074af53a2484a74b) +
                      (({q0_1[101],q0_0[101]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[101],q0_0[101]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I30e06d190906bc9eb6f1c3156c47f9f1  <=
                      (I8b3b875c6c07bd97ba598a5139156fa4) +
                      (({q0_1[102],q0_0[102]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[102],q0_0[102]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ieaaaced47e22029ad2945eac9cc45e6c  <=
                      (I7b33ddad346077928620344542b9481e) +
                      (({q0_1[103],q0_0[103]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[103],q0_0[103]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I08dc6f8e837b1f6b80bd3fc742290dab  <=
                      (I11d967a5c5d14c88b5587d4cfed1d05f) +
                      (({q0_1[104],q0_0[104]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[104],q0_0[104]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I8eb6a9c907c5909dad6cda98022d70b8  <=
                      (I27458d76b3ac6520fb379405c6b2956f) +
                      (({q0_1[105],q0_0[105]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[105],q0_0[105]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ia5067b1b458af82c3c2cd50653099854  <=
                      (I2525111a2fb5f10d64bbd16e148653b8) +
                      (({q0_1[106],q0_0[106]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[106],q0_0[106]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I198c6753cf12d423c709d1512e66fa9b  <=
                      (I7b7cbcd1c6d2a2eeaaff474536a69eed) +
                      (({q0_1[107],q0_0[107]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[107],q0_0[107]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ib600dd8a39fda48d28e1289d44d49a84  <=
                      (Id2a7f0781d18dccc7c4e0b383b7cddfa) +
                      (({q0_1[108],q0_0[108]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[108],q0_0[108]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Iabf09191227584c76d7fbc634b706d12  <=
                      (If8bc141d98ebe1be7fa81cde5c65868e) +
                      (({q0_1[109],q0_0[109]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[109],q0_0[109]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I4869ba08cab90a6dcbc454b0001a7a20  <=
                      (I8645e1326c66f5efef4b9c923599d1a3) +
                      (({q0_1[110],q0_0[110]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[110],q0_0[110]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               If97974406672507f8c9a1c507c4b6951  <=
                      (I0426ef66185128dd1ef4dbb68dcda585) +
                      (({q0_1[111],q0_0[111]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[111],q0_0[111]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I4210341f99ac7cb08245137999739114  <=
                      (Iddd954df5bae9b4240e0512f746669a9) +
                      (({q0_1[112],q0_0[112]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[112],q0_0[112]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ic24f4dbd99c8f4d88c8450d4fef762b8  <=
                      (I29e940970d87e8e09b26ab1b0b8f2286) +
                      (({q0_1[113],q0_0[113]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[113],q0_0[113]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I68dffa1a13eb6ab54615347729c1d6af  <=
                      (I488f6d9676aa85a55d030bf12e8997a7) +
                      (({q0_1[114],q0_0[114]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[114],q0_0[114]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I10153d5548b184b9ac2cecdba4ec4b1a  <=
                      (I99d761b75ade1fb2e8afbb1a77752609) +
                      (({q0_1[115],q0_0[115]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[115],q0_0[115]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I104b7f0512440cffc0fcce25e477f537  <=
                      (Iac4e3d20178049f9c59abf374752dccc) +
                      (({q0_1[116],q0_0[116]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[116],q0_0[116]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I18b6758319272eebbe76e1eee5ae55b2  <=
                      (I618d33f26badabfa578908903a613bce) +
                      (({q0_1[117],q0_0[117]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[117],q0_0[117]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I780263b10b98f9bb0eaf66c045d8d37c  <=
                      (I822d7973afe090b2764335f1b72dfd0e) +
                      (({q0_1[118],q0_0[118]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[118],q0_0[118]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I37b772442e55cbcd44ba892a0608d662  <=
                      (I12c1035353e553b3b6a13bb174ce6020) +
                      (({q0_1[119],q0_0[119]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[119],q0_0[119]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I0ac256a6659ff5c6673fd110a8bf578f  <=
                      (Ia6d61947d36fc128c689808c82db80f6) +
                      (({q0_1[120],q0_0[120]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[120],q0_0[120]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               If134e1d27e736005e5a390e7a2ea1f4b  <=
                      (Ie9b042f686381739b9ff219041f1e0ce) +
                      (({q0_1[121],q0_0[121]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[121],q0_0[121]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I7b37b8f908cd82683832536e02faab0d  <=
                      (I0c4268c01aed70ce4fc71531bf4bb862) +
                      (({q0_1[122],q0_0[122]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[122],q0_0[122]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I08b4bf60c9c7e7229bd1952cc88bc7b3  <=
                      (Ia34e42f8de91fa4861b0c6cac5dcfc29) +
                      (({q0_1[123],q0_0[123]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[123],q0_0[123]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I267d637eb63fef9f4723f7978fad88f0  <=
                      (Ib7c5850b4f7cc77be2048d114a2128d9) +
                      (({q0_1[124],q0_0[124]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[124],q0_0[124]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I4fb56a70e5ffa71f58f715da36368e04  <=
                      (I32bb50faa2b246b2d3b462a79be597c5) +
                      (({q0_1[125],q0_0[125]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[125],q0_0[125]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I5e9e2acb258baf96ac4b525bba54a462  <=
                      (Idc6d40a49f05c5422758cee50f787eb1) +
                      (({q0_1[126],q0_0[126]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[126],q0_0[126]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ic40f61443a4d8f87769067fc39381cb3  <=
                      (Ide1d7dc22a4b271ef764df14ac22366a) +
                      (({q0_1[127],q0_0[127]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[127],q0_0[127]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ieb36710c9a3726f33407436d62639c8d  <=
                      (I7ace6778ac86b3e05939a3fcc716136f) +
                      (({q0_1[128],q0_0[128]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[128],q0_0[128]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ic804af393da2e4b9c8ef25d4a3b4e8d5  <=
                      (I044e01e8d2df46e03f00a0af2beb0bf5) +
                      (({q0_1[129],q0_0[129]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[129],q0_0[129]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I52e4c446693c29a42bb3b665f72d382d  <=
                      (I45a7ddcda2662e36b7617dfe64514346) +
                      (({q0_1[130],q0_0[130]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[130],q0_0[130]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Idbf02cf10add496d30fa44bbb18458c6  <=
                      (Idada779a1ac7b844867571d77054b657) +
                      (({q0_1[131],q0_0[131]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[131],q0_0[131]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ida095585ad26e215f1c1bf989912da89  <=
                      (Ieeba01b18a244ab8c0ac263c138fabcc) +
                      (({q0_1[132],q0_0[132]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[132],q0_0[132]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I19f1ffa05c7c9a0df5e7014044024c7b  <=
                      (Ie4c9797a955778694dd8615219cb51e7) +
                      (({q0_1[133],q0_0[133]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[133],q0_0[133]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I4d68a2fe778fa93faac38b138138291f  <=
                      (I28a5ed4c239e64c76bb6e566b50cfd23) +
                      (({q0_1[134],q0_0[134]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[134],q0_0[134]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I54393ada6f76ac82c31f2668e228e29d  <=
                      (I79a705ee1e414fe4a5fb14e9b3ce9597) +
                      (({q0_1[135],q0_0[135]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[135],q0_0[135]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               If5b9ef84f09680f3593250b13a852c1c  <=
                      (I04f90a907f10a7fa1ae3591b48094d5c) +
                      (({q0_1[136],q0_0[136]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[136],q0_0[136]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ibb759bc4179e5b7aa759d850c7cfa467  <=
                      (I31d25b1b49e65216e90b39aa27acd6be) +
                      (({q0_1[137],q0_0[137]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[137],q0_0[137]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I05e8b5f8b83f07b609b5ebf272bb2229  <=
                      (I1f6540c5f037d861dee2c0091cba01ec) +
                      (({q0_1[138],q0_0[138]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[138],q0_0[138]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               If6ac15373ec1146d38e7aeb71c3ece64  <=
                      (I9632bb500b7faaaaeb649d74c21cbe8c) +
                      (({q0_1[139],q0_0[139]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[139],q0_0[139]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I2ab3675e1eede757af80716ba980a4e6  <=
                      (Idd0217a35c3adc8abc7bb581a5df7a2d) +
                      (({q0_1[140],q0_0[140]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[140],q0_0[140]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I388c271687ab31b57421ad57192273ed  <=
                      (Ic05b46168884322644db4e331d37d759) +
                      (({q0_1[141],q0_0[141]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[141],q0_0[141]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I6121679cec8caa51dc5ff0d1a61f9821  <=
                      (I53c88dc237bb2cd02d50fd7f0a168a48) +
                      (({q0_1[142],q0_0[142]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[142],q0_0[142]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ia0649b990bf5716cfab230127cd5d47f  <=
                      (I7450d4ab3ef0227e93a02bfd620d047b) +
                      (({q0_1[143],q0_0[143]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[143],q0_0[143]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I867a0626ca22108b16267d95c0aadf4f  <=
                      (I2b16e5b4e279bb29c3c675b72083e5fe) +
                      (({q0_1[144],q0_0[144]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[144],q0_0[144]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I1af54bcb73d7c6b93e55450871207976  <=
                      (I70c92e8ada46476d15ef4b3c620d2601) +
                      (({q0_1[145],q0_0[145]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[145],q0_0[145]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I91883553543d0425e9c6dd726dce3d27  <=
                      (Ib193b07804d6d5f111b06bda487bfa5f) +
                      (({q0_1[146],q0_0[146]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[146],q0_0[146]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ie95405659701278e3f87bf1f823a037b  <=
                      (I885433b0ab16c6d87abe45af13c9e529) +
                      (({q0_1[147],q0_0[147]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[147],q0_0[147]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ia42392e2104b50c0908aad82738a5ee7  <=
                      (I198c055930cb89d0390c336eda8fed4f) +
                      (({q0_1[148],q0_0[148]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[148],q0_0[148]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I68ad63230a51b9b9e3daffb307ea970d  <=
                      (I688a2c72e69b217d2673e8da75146a83) +
                      (({q0_1[149],q0_0[149]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[149],q0_0[149]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I7a052d63944ccf42e598efe3a95b88f8  <=
                      (I3b6fde4ed14cd68af1468ae1d4cc1a22) +
                      (({q0_1[150],q0_0[150]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[150],q0_0[150]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I2b3c6d69f79c8d51e4d1614c62c44fcc  <=
                      (I5d3df1e7563630311f56143ee6d97a8e) +
                      (({q0_1[151],q0_0[151]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[151],q0_0[151]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ifcef0e92f50e3920bf1208af5d64c632  <=
                      (I90a7ea789d3bf7f9126c786474a56da0) +
                      (({q0_1[152],q0_0[152]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[152],q0_0[152]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I111340a19625901a3c1b95fd0bd1570e  <=
                      (I5029424c9d9fe923eeb858b1e62cd758) +
                      (({q0_1[153],q0_0[153]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[153],q0_0[153]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I11aec4fa85c30f6fe1fd9fa72542ef6c  <=
                      (I1e805c70d50c2765b4a03ad2982dc421) +
                      (({q0_1[154],q0_0[154]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[154],q0_0[154]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I80cc333c181c16a96b7bd6501c27c2b3  <=
                      (Iba58175a7fd5c5da650222193caff0b3) +
                      (({q0_1[155],q0_0[155]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[155],q0_0[155]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Idc6354325a6280ae9890da33c06c33ec  <=
                      (I7401a0501ba69c5559fbf00c77e58dc5) +
                      (({q0_1[156],q0_0[156]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[156],q0_0[156]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ibb04cf82acc4ac16599ad3ddb0c2ada2  <=
                      (Idd9f7ea657ea9cdcb45a7e4b573b9d50) +
                      (({q0_1[157],q0_0[157]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[157],q0_0[157]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I3ed096dfd8a14f4acb4d53a70cf8aceb  <=
                      (I53f275395dd6be17961a5edc3e8da7f2) +
                      (({q0_1[158],q0_0[158]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[158],q0_0[158]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I0fa07f95e96326cb0599c0c3f76e2b48  <=
                      (Icab010d78cd66b02e089c74f04bf4e75) +
                      (({q0_1[159],q0_0[159]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[159],q0_0[159]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I87d98fbc97d9a78c2e7d6a6280e7a49a  <=
                      (I376a48b7e0195a5aacc76a0ad8bd14b2) +
                      (({q0_1[160],q0_0[160]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[160],q0_0[160]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ib7ddc4dca877f7cf5697a02c3d1915ba  <=
                      (I241622b0367dde514f96ece55c8c3964) +
                      (({q0_1[161],q0_0[161]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[161],q0_0[161]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I3612ef280891f6017fad205d0484bde7  <=
                      (If94a1abfb972f63629d07e64dc23863c) +
                      (({q0_1[162],q0_0[162]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[162],q0_0[162]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I561547649aeb5b4c3f10d9506db1f3cf  <=
                      (I07b9b1f4fa01b16cc69356057d3b6154) +
                      (({q0_1[163],q0_0[163]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[163],q0_0[163]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I84cc76c0079b86da7b994844c3ccb875  <=
                      (I2288a6ad3b748b716249f4adc42d52c4) +
                      (({q0_1[164],q0_0[164]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[164],q0_0[164]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Iec013c508d0c6401d7eb856e7eb60446  <=
                      (I022df337bcc05ac5648b8ae2e42f3a76) +
                      (({q0_1[165],q0_0[165]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[165],q0_0[165]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ifd8979aac6b6b24aa560b46b18240e92  <=
                      (I60d9a7f95fb8623753002ecaf9a4efcc) +
                      (({q0_1[166],q0_0[166]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[166],q0_0[166]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               If12394e78dc913b01890b56650856a44  <=
                      (I23a74ea5e7174d95e6d16a5e85ac236b) +
                      (({q0_1[167],q0_0[167]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[167],q0_0[167]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I94d18aa10695f3f22b23246884b72822  <=
                      (Ie697d28d757df82b3901564bda43251c) +
                      (({q0_1[168],q0_0[168]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[168],q0_0[168]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ic90b38835dd7e760dd54067b196f8470  <=
                      (I8572aedc94f7243ce5eacb332c81eae2) +
                      (({q0_1[169],q0_0[169]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[169],q0_0[169]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               If3691ea51f6efe9b165a31964854d2fe  <=
                      (I6734123aaf6320da75638b212812732f) +
                      (({q0_1[170],q0_0[170]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[170],q0_0[170]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ic2ce582555add38a14f5006d3c87eb15  <=
                      (I7f6dc6f0f403c58f9aaaa70c2383a666) +
                      (({q0_1[171],q0_0[171]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[171],q0_0[171]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I58cc950ee2cbe56b7c5a619be3792511  <=
                      (I66391978843c39b6acbdb4847a01050a) +
                      (({q0_1[172],q0_0[172]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[172],q0_0[172]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I0d8e329ec5873db96df1ec309445a096  <=
                      (I4f756e4125c8af5c412944b273e01cb0) +
                      (({q0_1[173],q0_0[173]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[173],q0_0[173]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I106325488e2ecfdba1cf9e5201e6bc8c  <=
                      (Id2c9f7ac95de07148c54803f69347f56) +
                      (({q0_1[174],q0_0[174]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[174],q0_0[174]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Iff73a0085541a511d3912b64686a82c5  <=
                      (I5061e13a179d27e1ba5f89ce8ee0fd4a) +
                      (({q0_1[175],q0_0[175]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[175],q0_0[175]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Icdab59de68f2870504598c9ea18f1d2c  <=
                      (I0f7c32fc1548fb49b8041f55c157498a) +
                      (({q0_1[176],q0_0[176]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[176],q0_0[176]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I75604d727e82c977741f90113719183a  <=
                      (I89ffab735ee30423c82e079ed98216c5) +
                      (({q0_1[177],q0_0[177]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[177],q0_0[177]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I6f50c4d0d2639857b2dcca300c2d7b04  <=
                      (I9494921d8487ee0b314f75cf0380fd2f) +
                      (({q0_1[178],q0_0[178]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[178],q0_0[178]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I5cd013a2be2e761c10c6a957632517de  <=
                      (If2b3e7d1541cbd8ffc2b4cfc3ad13a57) +
                      (({q0_1[179],q0_0[179]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[179],q0_0[179]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Iafeedddd02428bd2610c576e68d4ae25  <=
                      (Idf3d79da44f2d686f5bd43c3c1427430) +
                      (({q0_1[180],q0_0[180]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[180],q0_0[180]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I912d6325e34180e0f668f0f024e63581  <=
                      (If8125ad3c9e7f0a2b84106064d320996) +
                      (({q0_1[181],q0_0[181]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[181],q0_0[181]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Id1e05294dfd02df499ad0c08bb5c191b  <=
                      (Ic9018b88fa91fb638bbab0613795ae13) +
                      (({q0_1[182],q0_0[182]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[182],q0_0[182]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Id3bb9b100ee4302473b49ac14615e9b0  <=
                      (Iad4ea0196eb32f9a152c9e6fe5059e46) +
                      (({q0_1[183],q0_0[183]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[183],q0_0[183]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ief32db1cfc443119b6202b0cc7bf70a2  <=
                      (Ia8ff29ed728e7f2ae4213f00328b495d) +
                      (({q0_1[184],q0_0[184]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[184],q0_0[184]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Iad7dbe9909b5eed3261adf92d3813acc  <=
                      (I70717726200ec02929f679ef05496455) +
                      (({q0_1[185],q0_0[185]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[185],q0_0[185]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ie7daf0789c35caaadbba06cafabd2b70  <=
                      (Iaf1e4c7dae6ad89567836877c08f57d2) +
                      (({q0_1[186],q0_0[186]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[186],q0_0[186]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I2bd1f9b75d9ab94af9ddceb7528935e8  <=
                      (Icd09aa81e9b43528af73e23b2f0f80cb) +
                      (({q0_1[187],q0_0[187]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[187],q0_0[187]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ic3d9f5c6677758810e4865779ec303e3  <=
                      (I6ebb2b94f0f80425f8401ae823d92a1d) +
                      (({q0_1[188],q0_0[188]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[188],q0_0[188]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I00af04882a25e2832d913a67d4d86d7b  <=
                      (I4a2c3204a6a9936d4a215b46c0ffd045) +
                      (({q0_1[189],q0_0[189]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[189],q0_0[189]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ic9db631df0a1a9108c10c3e0eca7bf15  <=
                      (Ib02c0694762c4815448b2c8d3df767c2) +
                      (({q0_1[190],q0_0[190]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[190],q0_0[190]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I749f9ed1fb2dddd40ebc28f638e02935  <=
                      (I98cee6efbbe565d3a4de16703189782f) +
                      (({q0_1[191],q0_0[191]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[191],q0_0[191]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ia45b2a24df24bd5e3c95885c8928686c  <=
                      (Ibf981c01a9d44cbea3c6d8ead92bc2ab) +
                      (({q0_1[192],q0_0[192]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[192],q0_0[192]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I7427464fde340780aba7f9847b4ad564  <=
                      (I864c33e8ea204d20a9baef4584f22d4e) +
                      (({q0_1[193],q0_0[193]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[193],q0_0[193]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I33fd1ae225e2b881b2b41e0358675e22  <=
                      (I6ad3228e0e2e1f19648d73e83ba5a229) +
                      (({q0_1[194],q0_0[194]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[194],q0_0[194]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I2e21a35d1cf560936fd19b944a208b6b  <=
                      (Ie099210a99a4899c53baf39559592690) +
                      (({q0_1[195],q0_0[195]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[195],q0_0[195]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I249522a3d42cc75d7a6b9ede1222ee76  <=
                      (Ieeec71d9df4613555fade2ced7b3baf1) +
                      (({q0_1[196],q0_0[196]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[196],q0_0[196]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I68b4c43d9f40ae4bfd70d2983594392c  <=
                      (I4931884e3544af182bcda9061091a42d) +
                      (({q0_1[197],q0_0[197]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[197],q0_0[197]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I63145e0fec15c7e7c0de105f348bfd31  <=
                      (Ib3fb10da528d450251764a9b9ede0dba) +
                      (({q0_1[198],q0_0[198]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[198],q0_0[198]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I8af625de86c04016c3424d116fddab5b  <=
                      (Icdc9e676957b2223d60c413331fa982f) +
                      (({q0_1[199],q0_0[199]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[199],q0_0[199]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I54c9c10527f83b4ee4e1e22f1e4044ed  <=
                      (I381f6051282c062ccf53866830344cd4) +
                      (({q0_1[200],q0_0[200]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[200],q0_0[200]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I972559e47c7f83bd9000ca1cfc14d8e0  <=
                      (Icfc21935c007fbbceb2a67ebe1a68a0b) +
                      (({q0_1[201],q0_0[201]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[201],q0_0[201]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ib97a7f941eb7ce2a867503a04ff86a67  <=
                      (I120d597a80158374726e064fb0f099fb) +
                      (({q0_1[202],q0_0[202]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[202],q0_0[202]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I5979b55f607c71017537f2b48b40cbea  <=
                      (I2520aa556aadf851f58f0b1820498730) +
                      (({q0_1[203],q0_0[203]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[203],q0_0[203]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I6a56760b621f238843b091279c69897f  <=
                      (I6203f49a08107f7185ebadeecf2c16b0) +
                      (({q0_1[204],q0_0[204]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[204],q0_0[204]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Icec45bf76c241d37c9a50a5cd092da9d  <=
                      (Ia706fb593b63cebbee0321c154cb859b) +
                      (({q0_1[205],q0_0[205]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[205],q0_0[205]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I2f6d3f61f2890e584d3063a09587e99b  <=
                      (Ia4b5f2b07556629673fc6576bc49a5dc) +
                      (({q0_1[206],q0_0[206]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[206],q0_0[206]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I7c396ea2e959d84fd9a6964617cb29c6  <=
                      (Ic532c6b85b156f821e0742f47239a65c) +
                      (({q0_1[207],q0_0[207]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[207],q0_0[207]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"

                 if ({q0_1[0],q0_0[0]} != 1 ) begin
                 end
                 if ({q0_1[1],q0_0[1]} != 1 ) begin
                 end
                 if ({q0_1[2],q0_0[2]} != 0 ) begin
                 end
                 if ({q0_1[3],q0_0[3]} != 0 ) begin
                 end
                 if ({q0_1[4],q0_0[4]} != 0 ) begin
                 end
                 if ({q0_1[5],q0_0[5]} != 0 ) begin
                 end
                 if ({q0_1[6],q0_0[6]} != 0 ) begin
                 end
                 if ({q0_1[7],q0_0[7]} != 1 ) begin
                 end
                 if ({q0_1[8],q0_0[8]} != 0 ) begin
                 end
                 if ({q0_1[9],q0_0[9]} != 1 ) begin
                 end
                 if ({q0_1[10],q0_0[10]} != 1 ) begin
                 end
                 if ({q0_1[11],q0_0[11]} != 1 ) begin
                 end
                 if ({q0_1[12],q0_0[12]} != 0 ) begin
                 end
                 if ({q0_1[13],q0_0[13]} != 0 ) begin
                 end
                 if ({q0_1[14],q0_0[14]} != 1 ) begin
                 end
                 if ({q0_1[15],q0_0[15]} != 1 ) begin
                 end
                 if ({q0_1[16],q0_0[16]} != 0 ) begin
                 end
                 if ({q0_1[17],q0_0[17]} != 0 ) begin
                 end
                 if ({q0_1[18],q0_0[18]} != 1 ) begin
                 end
                 if ({q0_1[19],q0_0[19]} != 0 ) begin
                 end
                 if ({q0_1[20],q0_0[20]} != 1 ) begin
                 end
                 if ({q0_1[21],q0_0[21]} != 1 ) begin
                 end
                 if ({q0_1[22],q0_0[22]} != 1 ) begin
                 end
                 if ({q0_1[23],q0_0[23]} != 0 ) begin
                 end
                 if ({q0_1[24],q0_0[24]} != 1 ) begin
                 end
                 if ({q0_1[25],q0_0[25]} != 1 ) begin
                 end
                 if ({q0_1[26],q0_0[26]} != 1 ) begin
                 end
                 if ({q0_1[27],q0_0[27]} != 0 ) begin
                 end
                 if ({q0_1[28],q0_0[28]} != 0 ) begin
                 end
                 if ({q0_1[29],q0_0[29]} != 1 ) begin
                 end
                 if ({q0_1[30],q0_0[30]} != 1 ) begin
                 end
                 if ({q0_1[31],q0_0[31]} != 1 ) begin
                 end
                 if ({q0_1[32],q0_0[32]} != 0 ) begin
                 end
                 if ({q0_1[33],q0_0[33]} != 0 ) begin
                 end
                 if ({q0_1[34],q0_0[34]} != 1 ) begin
                 end
                 if ({q0_1[35],q0_0[35]} != 0 ) begin
                 end
                 if ({q0_1[36],q0_0[36]} != 0 ) begin
                 end
                 if ({q0_1[37],q0_0[37]} != 0 ) begin
                 end
                 if ({q0_1[38],q0_0[38]} != 0 ) begin
                 end
                 if ({q0_1[39],q0_0[39]} != 0 ) begin
                 end
                 if ({q0_1[40],q0_0[40]} != 1 ) begin
                 end
                 if ({q0_1[41],q0_0[41]} != 0 ) begin
                 end
                 if ({q0_1[42],q0_0[42]} != 0 ) begin
                 end
                 if ({q0_1[43],q0_0[43]} != 0 ) begin
                 end
                 if ({q0_1[44],q0_0[44]} != 1 ) begin
                 end
                 if ({q0_1[45],q0_0[45]} != 1 ) begin
                 end
                 if ({q0_1[46],q0_0[46]} != 1 ) begin
                 end
                 if ({q0_1[47],q0_0[47]} != 0 ) begin
                 end
                 if ({q0_1[48],q0_0[48]} != 0 ) begin
                 end
                 if ({q0_1[49],q0_0[49]} != 1 ) begin
                 end
                 if ({q0_1[50],q0_0[50]} != 0 ) begin
                 end
                 if ({q0_1[51],q0_0[51]} != 0 ) begin
                 end
                 if ({q0_1[52],q0_0[52]} != 1 ) begin
                 end
                 if ({q0_1[53],q0_0[53]} != 1 ) begin
                 end
                 if ({q0_1[54],q0_0[54]} != 0 ) begin
                 end
                 if ({q0_1[55],q0_0[55]} != 1 ) begin
                 end
                 if ({q0_1[56],q0_0[56]} != 1 ) begin
                 end
                 if ({q0_1[57],q0_0[57]} != 0 ) begin
                 end
                 if ({q0_1[58],q0_0[58]} != 0 ) begin
                 end
                 if ({q0_1[59],q0_0[59]} != 1 ) begin
                 end
                 if ({q0_1[60],q0_0[60]} != 0 ) begin
                 end
                 if ({q0_1[61],q0_0[61]} != 0 ) begin
                 end
                 if ({q0_1[62],q0_0[62]} != 1 ) begin
                 end
                 if ({q0_1[63],q0_0[63]} != 0 ) begin
                 end
                 if ({q0_1[64],q0_0[64]} != 1 ) begin
                 end
                 if ({q0_1[65],q0_0[65]} != 1 ) begin
                 end
                 if ({q0_1[66],q0_0[66]} != 1 ) begin
                 end
                 if ({q0_1[67],q0_0[67]} != 1 ) begin
                 end
                 if ({q0_1[68],q0_0[68]} != 1 ) begin
                 end
                 if ({q0_1[69],q0_0[69]} != 1 ) begin
                 end
                 if ({q0_1[70],q0_0[70]} != 1 ) begin
                 end
                 if ({q0_1[71],q0_0[71]} != 1 ) begin
                 end
                 if ({q0_1[72],q0_0[72]} != 0 ) begin
                 end
                 if ({q0_1[73],q0_0[73]} != 0 ) begin
                 end
                 if ({q0_1[74],q0_0[74]} != 0 ) begin
                 end
                 if ({q0_1[75],q0_0[75]} != 0 ) begin
                 end
                 if ({q0_1[76],q0_0[76]} != 0 ) begin
                 end
                 if ({q0_1[77],q0_0[77]} != 0 ) begin
                 end
                 if ({q0_1[78],q0_0[78]} != 1 ) begin
                 end
                 if ({q0_1[79],q0_0[79]} != 0 ) begin
                 end
                 if ({q0_1[80],q0_0[80]} != 0 ) begin
                 end
                 if ({q0_1[81],q0_0[81]} != 1 ) begin
                 end
                 if ({q0_1[82],q0_0[82]} != 1 ) begin
                 end
                 if ({q0_1[83],q0_0[83]} != 0 ) begin
                 end
                 if ({q0_1[84],q0_0[84]} != 0 ) begin
                 end
                 if ({q0_1[85],q0_0[85]} != 0 ) begin
                 end
                 if ({q0_1[86],q0_0[86]} != 0 ) begin
                 end
                 if ({q0_1[87],q0_0[87]} != 0 ) begin
                 end
                 if ({q0_1[88],q0_0[88]} != 1 ) begin
                 end
                 if ({q0_1[89],q0_0[89]} != 1 ) begin
                 end
                 if ({q0_1[90],q0_0[90]} != 0 ) begin
                 end
                 if ({q0_1[91],q0_0[91]} != 1 ) begin
                 end
                 if ({q0_1[92],q0_0[92]} != 0 ) begin
                 end
                 if ({q0_1[93],q0_0[93]} != 0 ) begin
                 end
                 if ({q0_1[94],q0_0[94]} != 0 ) begin
                 end
                 if ({q0_1[95],q0_0[95]} != 0 ) begin
                 end
                 if ({q0_1[96],q0_0[96]} != 0 ) begin
                 end
                 if ({q0_1[97],q0_0[97]} != 1 ) begin
                 end
                 if ({q0_1[98],q0_0[98]} != 0 ) begin
                 end
                 if ({q0_1[99],q0_0[99]} != 0 ) begin
                 end
                 if ({q0_1[100],q0_0[100]} != 0 ) begin
                 end
                 if ({q0_1[101],q0_0[101]} != 1 ) begin
                 end
                 if ({q0_1[102],q0_0[102]} != 1 ) begin
                 end
                 if ({q0_1[103],q0_0[103]} != 1 ) begin
                 end
                 if ({q0_1[104],q0_0[104]} != 1 ) begin
                 end
                 if ({q0_1[105],q0_0[105]} != 1 ) begin
                 end
                 if ({q0_1[106],q0_0[106]} != 1 ) begin
                 end
                 if ({q0_1[107],q0_0[107]} != 1 ) begin
                 end
                 if ({q0_1[108],q0_0[108]} != 0 ) begin
                 end
                 if ({q0_1[109],q0_0[109]} != 0 ) begin
                 end
                 if ({q0_1[110],q0_0[110]} != 0 ) begin
                 end
                 if ({q0_1[111],q0_0[111]} != 1 ) begin
                 end
                 if ({q0_1[112],q0_0[112]} != 0 ) begin
                 end
                 if ({q0_1[113],q0_0[113]} != 1 ) begin
                 end
                 if ({q0_1[114],q0_0[114]} != 0 ) begin
                 end
                 if ({q0_1[115],q0_0[115]} != 0 ) begin
                 end
                 if ({q0_1[116],q0_0[116]} != 0 ) begin
                 end
                 if ({q0_1[117],q0_0[117]} != 1 ) begin
                 end
                 if ({q0_1[118],q0_0[118]} != 1 ) begin
                 end
                 if ({q0_1[119],q0_0[119]} != 0 ) begin
                 end
                 if ({q0_1[120],q0_0[120]} != 1 ) begin
                 end
                 if ({q0_1[121],q0_0[121]} != 0 ) begin
                 end
                 if ({q0_1[122],q0_0[122]} != 0 ) begin
                 end
                 if ({q0_1[123],q0_0[123]} != 1 ) begin
                 end
                 if ({q0_1[124],q0_0[124]} != 0 ) begin
                 end
                 if ({q0_1[125],q0_0[125]} != 0 ) begin
                 end
                 if ({q0_1[126],q0_0[126]} != 1 ) begin
                 end
                 if ({q0_1[127],q0_0[127]} != 0 ) begin
                 end
                 if ({q0_1[128],q0_0[128]} != 1 ) begin
                 end
                 if ({q0_1[129],q0_0[129]} != 0 ) begin
                 end
                 if ({q0_1[130],q0_0[130]} != 0 ) begin
                 end
                 if ({q0_1[131],q0_0[131]} != 0 ) begin
                 end
                 if ({q0_1[132],q0_0[132]} != 0 ) begin
                 end
                 if ({q0_1[133],q0_0[133]} != 1 ) begin
                 end
                 if ({q0_1[134],q0_0[134]} != 1 ) begin
                 end
                 if ({q0_1[135],q0_0[135]} != 1 ) begin
                 end
                 if ({q0_1[136],q0_0[136]} != 1 ) begin
                 end
                 if ({q0_1[137],q0_0[137]} != 0 ) begin
                 end
                 if ({q0_1[138],q0_0[138]} != 0 ) begin
                 end
                 if ({q0_1[139],q0_0[139]} != 1 ) begin
                 end
                 if ({q0_1[140],q0_0[140]} != 1 ) begin
                 end
                 if ({q0_1[141],q0_0[141]} != 1 ) begin
                 end
                 if ({q0_1[142],q0_0[142]} != 0 ) begin
                 end
                 if ({q0_1[143],q0_0[143]} != 0 ) begin
                 end
                 if ({q0_1[144],q0_0[144]} != 1 ) begin
                 end
                 if ({q0_1[145],q0_0[145]} != 1 ) begin
                 end
                 if ({q0_1[146],q0_0[146]} != 0 ) begin
                 end
                 if ({q0_1[147],q0_0[147]} != 1 ) begin
                 end
                 if ({q0_1[148],q0_0[148]} != 1 ) begin
                 end
                 if ({q0_1[149],q0_0[149]} != 1 ) begin
                 end
                 if ({q0_1[150],q0_0[150]} != 1 ) begin
                 end
                 if ({q0_1[151],q0_0[151]} != 0 ) begin
                 end
                 if ({q0_1[152],q0_0[152]} != 1 ) begin
                 end
                 if ({q0_1[153],q0_0[153]} != 0 ) begin
                 end
                 if ({q0_1[154],q0_0[154]} != 0 ) begin
                 end
                 if ({q0_1[155],q0_0[155]} != 0 ) begin
                 end
                 if ({q0_1[156],q0_0[156]} != 0 ) begin
                 end
                 if ({q0_1[157],q0_0[157]} != 1 ) begin
                 end
                 if ({q0_1[158],q0_0[158]} != 0 ) begin
                 end
                 if ({q0_1[159],q0_0[159]} != 1 ) begin
                 end
                 if ({q0_1[160],q0_0[160]} != 1 ) begin
                 end
                 if ({q0_1[161],q0_0[161]} != 1 ) begin
                 end
                 if ({q0_1[162],q0_0[162]} != 0 ) begin
                 end
                 if ({q0_1[163],q0_0[163]} != 1 ) begin
                 end
                 if ({q0_1[164],q0_0[164]} != 0 ) begin
                 end
                 if ({q0_1[165],q0_0[165]} != 1 ) begin
                 end
                 if ({q0_1[166],q0_0[166]} != 1 ) begin
                 end
                 if ({q0_1[167],q0_0[167]} != 0 ) begin
                 end
                 if ({q0_1[168],q0_0[168]} != 0 ) begin
                 end
                 if ({q0_1[169],q0_0[169]} != 1 ) begin
                 end
                 if ({q0_1[170],q0_0[170]} != 1 ) begin
                 end
                 if ({q0_1[171],q0_0[171]} != 0 ) begin
                 end
                 if ({q0_1[172],q0_0[172]} != 1 ) begin
                 end
                 if ({q0_1[173],q0_0[173]} != 1 ) begin
                 end
                 if ({q0_1[174],q0_0[174]} != 0 ) begin
                 end
                 if ({q0_1[175],q0_0[175]} != 0 ) begin
                 end
                 if ({q0_1[176],q0_0[176]} != 1 ) begin
                 end
                 if ({q0_1[177],q0_0[177]} != 0 ) begin
                 end
                 if ({q0_1[178],q0_0[178]} != 1 ) begin
                 end
                 if ({q0_1[179],q0_0[179]} != 1 ) begin
                 end
                 if ({q0_1[180],q0_0[180]} != 0 ) begin
                 end
                 if ({q0_1[181],q0_0[181]} != 0 ) begin
                 end
                 if ({q0_1[182],q0_0[182]} != 1 ) begin
                 end
                 if ({q0_1[183],q0_0[183]} != 1 ) begin
                 end
                 if ({q0_1[184],q0_0[184]} != 1 ) begin
                 end
                 if ({q0_1[185],q0_0[185]} != 1 ) begin
                 end
                 if ({q0_1[186],q0_0[186]} != 0 ) begin
                 end
                 if ({q0_1[187],q0_0[187]} != 0 ) begin
                 end
                 if ({q0_1[188],q0_0[188]} != 0 ) begin
                 end
                 if ({q0_1[189],q0_0[189]} != 0 ) begin
                 end
                 if ({q0_1[190],q0_0[190]} != 0 ) begin
                 end
                 if ({q0_1[191],q0_0[191]} != 0 ) begin
                 end
                 if ({q0_1[192],q0_0[192]} != 1 ) begin
                 end
                 if ({q0_1[193],q0_0[193]} != 0 ) begin
                 end
                 if ({q0_1[194],q0_0[194]} != 1 ) begin
                 end
                 if ({q0_1[195],q0_0[195]} != 1 ) begin
                 end
                 if ({q0_1[196],q0_0[196]} != 0 ) begin
                 end
                 if ({q0_1[197],q0_0[197]} != 1 ) begin
                 end
                 if ({q0_1[198],q0_0[198]} != 0 ) begin
                 end
                 if ({q0_1[199],q0_0[199]} != 0 ) begin
                 end
                 if ({q0_1[200],q0_0[200]} != 0 ) begin
                 end
                 if ({q0_1[201],q0_0[201]} != 1 ) begin
                 end
                 if ({q0_1[202],q0_0[202]} != 1 ) begin
                 end
                 if ({q0_1[203],q0_0[203]} != 0 ) begin
                 end
                 if ({q0_1[204],q0_0[204]} != 0 ) begin
                 end
                 if ({q0_1[205],q0_0[205]} != 0 ) begin
                 end
                 if ({q0_1[206],q0_0[206]} != 1 ) begin
                 end
                 if ({q0_1[207],q0_0[207]} != 0 ) begin
                 end


           end

           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I95878a848ec38c4f334bc1915576e6d6[0]        <=  I583b1bfc712ec29d08acc68c27675882[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I583b1bfc712ec29d08acc68c27675882[0] + 1 :
                                             I583b1bfc712ec29d08acc68c27675882[0] ;
            Ib58043c04b5c4c86c1c67e57cc66dcf7[0]  <=  I583b1bfc712ec29d08acc68c27675882[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I95878a848ec38c4f334bc1915576e6d6[1]        <=  I583b1bfc712ec29d08acc68c27675882[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I583b1bfc712ec29d08acc68c27675882[1] + 1 :
                                             I583b1bfc712ec29d08acc68c27675882[1] ;
            Ib58043c04b5c4c86c1c67e57cc66dcf7[1]  <=  I583b1bfc712ec29d08acc68c27675882[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I95878a848ec38c4f334bc1915576e6d6[2]        <=  I583b1bfc712ec29d08acc68c27675882[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I583b1bfc712ec29d08acc68c27675882[2] + 1 :
                                             I583b1bfc712ec29d08acc68c27675882[2] ;
            Ib58043c04b5c4c86c1c67e57cc66dcf7[2]  <=  I583b1bfc712ec29d08acc68c27675882[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I95878a848ec38c4f334bc1915576e6d6[3]        <=  I583b1bfc712ec29d08acc68c27675882[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I583b1bfc712ec29d08acc68c27675882[3] + 1 :
                                             I583b1bfc712ec29d08acc68c27675882[3] ;
            Ib58043c04b5c4c86c1c67e57cc66dcf7[3]  <=  I583b1bfc712ec29d08acc68c27675882[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I95878a848ec38c4f334bc1915576e6d6[4]        <=  I583b1bfc712ec29d08acc68c27675882[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I583b1bfc712ec29d08acc68c27675882[4] + 1 :
                                             I583b1bfc712ec29d08acc68c27675882[4] ;
            Ib58043c04b5c4c86c1c67e57cc66dcf7[4]  <=  I583b1bfc712ec29d08acc68c27675882[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I95878a848ec38c4f334bc1915576e6d6[5]        <=  I583b1bfc712ec29d08acc68c27675882[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I583b1bfc712ec29d08acc68c27675882[5] + 1 :
                                             I583b1bfc712ec29d08acc68c27675882[5] ;
            Ib58043c04b5c4c86c1c67e57cc66dcf7[5]  <=  I583b1bfc712ec29d08acc68c27675882[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I95878a848ec38c4f334bc1915576e6d6[6]        <=  I583b1bfc712ec29d08acc68c27675882[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I583b1bfc712ec29d08acc68c27675882[6] + 1 :
                                             I583b1bfc712ec29d08acc68c27675882[6] ;
            Ib58043c04b5c4c86c1c67e57cc66dcf7[6]  <=  I583b1bfc712ec29d08acc68c27675882[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I95878a848ec38c4f334bc1915576e6d6[7]        <=  I583b1bfc712ec29d08acc68c27675882[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I583b1bfc712ec29d08acc68c27675882[7] + 1 :
                                             I583b1bfc712ec29d08acc68c27675882[7] ;
            Ib58043c04b5c4c86c1c67e57cc66dcf7[7]  <=  I583b1bfc712ec29d08acc68c27675882[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I95878a848ec38c4f334bc1915576e6d6[8]        <=  I583b1bfc712ec29d08acc68c27675882[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I583b1bfc712ec29d08acc68c27675882[8] + 1 :
                                             I583b1bfc712ec29d08acc68c27675882[8] ;
            Ib58043c04b5c4c86c1c67e57cc66dcf7[8]  <=  I583b1bfc712ec29d08acc68c27675882[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I95878a848ec38c4f334bc1915576e6d6[9]        <=  I583b1bfc712ec29d08acc68c27675882[9][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I583b1bfc712ec29d08acc68c27675882[9] + 1 :
                                             I583b1bfc712ec29d08acc68c27675882[9] ;
            Ib58043c04b5c4c86c1c67e57cc66dcf7[9]  <=  I583b1bfc712ec29d08acc68c27675882[9][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I95878a848ec38c4f334bc1915576e6d6[10]        <=  I583b1bfc712ec29d08acc68c27675882[10][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I583b1bfc712ec29d08acc68c27675882[10] + 1 :
                                             I583b1bfc712ec29d08acc68c27675882[10] ;
            Ib58043c04b5c4c86c1c67e57cc66dcf7[10]  <=  I583b1bfc712ec29d08acc68c27675882[10][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I95878a848ec38c4f334bc1915576e6d6[11]        <=  I583b1bfc712ec29d08acc68c27675882[11][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I583b1bfc712ec29d08acc68c27675882[11] + 1 :
                                             I583b1bfc712ec29d08acc68c27675882[11] ;
            Ib58043c04b5c4c86c1c67e57cc66dcf7[11]  <=  I583b1bfc712ec29d08acc68c27675882[11][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I95878a848ec38c4f334bc1915576e6d6[12]        <=  I583b1bfc712ec29d08acc68c27675882[12][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I583b1bfc712ec29d08acc68c27675882[12] + 1 :
                                             I583b1bfc712ec29d08acc68c27675882[12] ;
            Ib58043c04b5c4c86c1c67e57cc66dcf7[12]  <=  I583b1bfc712ec29d08acc68c27675882[12][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I95878a848ec38c4f334bc1915576e6d6[13]        <=  I583b1bfc712ec29d08acc68c27675882[13][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I583b1bfc712ec29d08acc68c27675882[13] + 1 :
                                             I583b1bfc712ec29d08acc68c27675882[13] ;
            Ib58043c04b5c4c86c1c67e57cc66dcf7[13]  <=  I583b1bfc712ec29d08acc68c27675882[13][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I95878a848ec38c4f334bc1915576e6d6[14]        <=  I583b1bfc712ec29d08acc68c27675882[14][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I583b1bfc712ec29d08acc68c27675882[14] + 1 :
                                             I583b1bfc712ec29d08acc68c27675882[14] ;
            Ib58043c04b5c4c86c1c67e57cc66dcf7[14]  <=  I583b1bfc712ec29d08acc68c27675882[14][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I95878a848ec38c4f334bc1915576e6d6[15]        <=  I583b1bfc712ec29d08acc68c27675882[15][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I583b1bfc712ec29d08acc68c27675882[15] + 1 :
                                             I583b1bfc712ec29d08acc68c27675882[15] ;
            Ib58043c04b5c4c86c1c67e57cc66dcf7[15]  <=  I583b1bfc712ec29d08acc68c27675882[15][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I95878a848ec38c4f334bc1915576e6d6[16]        <=  I583b1bfc712ec29d08acc68c27675882[16][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I583b1bfc712ec29d08acc68c27675882[16] + 1 :
                                             I583b1bfc712ec29d08acc68c27675882[16] ;
            Ib58043c04b5c4c86c1c67e57cc66dcf7[16]  <=  I583b1bfc712ec29d08acc68c27675882[16][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I95878a848ec38c4f334bc1915576e6d6[17]        <=  I583b1bfc712ec29d08acc68c27675882[17][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I583b1bfc712ec29d08acc68c27675882[17] + 1 :
                                             I583b1bfc712ec29d08acc68c27675882[17] ;
            Ib58043c04b5c4c86c1c67e57cc66dcf7[17]  <=  I583b1bfc712ec29d08acc68c27675882[17][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I95878a848ec38c4f334bc1915576e6d6[18]        <=  I583b1bfc712ec29d08acc68c27675882[18][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I583b1bfc712ec29d08acc68c27675882[18] + 1 :
                                             I583b1bfc712ec29d08acc68c27675882[18] ;
            Ib58043c04b5c4c86c1c67e57cc66dcf7[18]  <=  I583b1bfc712ec29d08acc68c27675882[18][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I95878a848ec38c4f334bc1915576e6d6[19]        <=  I583b1bfc712ec29d08acc68c27675882[19][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I583b1bfc712ec29d08acc68c27675882[19] + 1 :
                                             I583b1bfc712ec29d08acc68c27675882[19] ;
            Ib58043c04b5c4c86c1c67e57cc66dcf7[19]  <=  I583b1bfc712ec29d08acc68c27675882[19][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I95878a848ec38c4f334bc1915576e6d6[20]        <=  I583b1bfc712ec29d08acc68c27675882[20][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I583b1bfc712ec29d08acc68c27675882[20] + 1 :
                                             I583b1bfc712ec29d08acc68c27675882[20] ;
            Ib58043c04b5c4c86c1c67e57cc66dcf7[20]  <=  I583b1bfc712ec29d08acc68c27675882[20][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I95878a848ec38c4f334bc1915576e6d6[21]        <=  I583b1bfc712ec29d08acc68c27675882[21][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I583b1bfc712ec29d08acc68c27675882[21] + 1 :
                                             I583b1bfc712ec29d08acc68c27675882[21] ;
            Ib58043c04b5c4c86c1c67e57cc66dcf7[21]  <=  I583b1bfc712ec29d08acc68c27675882[21][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3eb1902edf9266038f39c281d134c26c[0]        <=  Ifba287889bea3585954fef5efdf5bb24[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ifba287889bea3585954fef5efdf5bb24[0] + 1 :
                                             Ifba287889bea3585954fef5efdf5bb24[0] ;
            Ibc0871b3c992fd278815fdbefcd2bac0[0]  <=  Ifba287889bea3585954fef5efdf5bb24[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3eb1902edf9266038f39c281d134c26c[1]        <=  Ifba287889bea3585954fef5efdf5bb24[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ifba287889bea3585954fef5efdf5bb24[1] + 1 :
                                             Ifba287889bea3585954fef5efdf5bb24[1] ;
            Ibc0871b3c992fd278815fdbefcd2bac0[1]  <=  Ifba287889bea3585954fef5efdf5bb24[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3eb1902edf9266038f39c281d134c26c[2]        <=  Ifba287889bea3585954fef5efdf5bb24[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ifba287889bea3585954fef5efdf5bb24[2] + 1 :
                                             Ifba287889bea3585954fef5efdf5bb24[2] ;
            Ibc0871b3c992fd278815fdbefcd2bac0[2]  <=  Ifba287889bea3585954fef5efdf5bb24[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3eb1902edf9266038f39c281d134c26c[3]        <=  Ifba287889bea3585954fef5efdf5bb24[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ifba287889bea3585954fef5efdf5bb24[3] + 1 :
                                             Ifba287889bea3585954fef5efdf5bb24[3] ;
            Ibc0871b3c992fd278815fdbefcd2bac0[3]  <=  Ifba287889bea3585954fef5efdf5bb24[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3eb1902edf9266038f39c281d134c26c[4]        <=  Ifba287889bea3585954fef5efdf5bb24[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ifba287889bea3585954fef5efdf5bb24[4] + 1 :
                                             Ifba287889bea3585954fef5efdf5bb24[4] ;
            Ibc0871b3c992fd278815fdbefcd2bac0[4]  <=  Ifba287889bea3585954fef5efdf5bb24[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3eb1902edf9266038f39c281d134c26c[5]        <=  Ifba287889bea3585954fef5efdf5bb24[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ifba287889bea3585954fef5efdf5bb24[5] + 1 :
                                             Ifba287889bea3585954fef5efdf5bb24[5] ;
            Ibc0871b3c992fd278815fdbefcd2bac0[5]  <=  Ifba287889bea3585954fef5efdf5bb24[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3eb1902edf9266038f39c281d134c26c[6]        <=  Ifba287889bea3585954fef5efdf5bb24[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ifba287889bea3585954fef5efdf5bb24[6] + 1 :
                                             Ifba287889bea3585954fef5efdf5bb24[6] ;
            Ibc0871b3c992fd278815fdbefcd2bac0[6]  <=  Ifba287889bea3585954fef5efdf5bb24[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3eb1902edf9266038f39c281d134c26c[7]        <=  Ifba287889bea3585954fef5efdf5bb24[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ifba287889bea3585954fef5efdf5bb24[7] + 1 :
                                             Ifba287889bea3585954fef5efdf5bb24[7] ;
            Ibc0871b3c992fd278815fdbefcd2bac0[7]  <=  Ifba287889bea3585954fef5efdf5bb24[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3eb1902edf9266038f39c281d134c26c[8]        <=  Ifba287889bea3585954fef5efdf5bb24[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ifba287889bea3585954fef5efdf5bb24[8] + 1 :
                                             Ifba287889bea3585954fef5efdf5bb24[8] ;
            Ibc0871b3c992fd278815fdbefcd2bac0[8]  <=  Ifba287889bea3585954fef5efdf5bb24[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3eb1902edf9266038f39c281d134c26c[9]        <=  Ifba287889bea3585954fef5efdf5bb24[9][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ifba287889bea3585954fef5efdf5bb24[9] + 1 :
                                             Ifba287889bea3585954fef5efdf5bb24[9] ;
            Ibc0871b3c992fd278815fdbefcd2bac0[9]  <=  Ifba287889bea3585954fef5efdf5bb24[9][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3eb1902edf9266038f39c281d134c26c[10]        <=  Ifba287889bea3585954fef5efdf5bb24[10][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ifba287889bea3585954fef5efdf5bb24[10] + 1 :
                                             Ifba287889bea3585954fef5efdf5bb24[10] ;
            Ibc0871b3c992fd278815fdbefcd2bac0[10]  <=  Ifba287889bea3585954fef5efdf5bb24[10][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3eb1902edf9266038f39c281d134c26c[11]        <=  Ifba287889bea3585954fef5efdf5bb24[11][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ifba287889bea3585954fef5efdf5bb24[11] + 1 :
                                             Ifba287889bea3585954fef5efdf5bb24[11] ;
            Ibc0871b3c992fd278815fdbefcd2bac0[11]  <=  Ifba287889bea3585954fef5efdf5bb24[11][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3eb1902edf9266038f39c281d134c26c[12]        <=  Ifba287889bea3585954fef5efdf5bb24[12][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ifba287889bea3585954fef5efdf5bb24[12] + 1 :
                                             Ifba287889bea3585954fef5efdf5bb24[12] ;
            Ibc0871b3c992fd278815fdbefcd2bac0[12]  <=  Ifba287889bea3585954fef5efdf5bb24[12][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3eb1902edf9266038f39c281d134c26c[13]        <=  Ifba287889bea3585954fef5efdf5bb24[13][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ifba287889bea3585954fef5efdf5bb24[13] + 1 :
                                             Ifba287889bea3585954fef5efdf5bb24[13] ;
            Ibc0871b3c992fd278815fdbefcd2bac0[13]  <=  Ifba287889bea3585954fef5efdf5bb24[13][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3eb1902edf9266038f39c281d134c26c[14]        <=  Ifba287889bea3585954fef5efdf5bb24[14][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ifba287889bea3585954fef5efdf5bb24[14] + 1 :
                                             Ifba287889bea3585954fef5efdf5bb24[14] ;
            Ibc0871b3c992fd278815fdbefcd2bac0[14]  <=  Ifba287889bea3585954fef5efdf5bb24[14][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3eb1902edf9266038f39c281d134c26c[15]        <=  Ifba287889bea3585954fef5efdf5bb24[15][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ifba287889bea3585954fef5efdf5bb24[15] + 1 :
                                             Ifba287889bea3585954fef5efdf5bb24[15] ;
            Ibc0871b3c992fd278815fdbefcd2bac0[15]  <=  Ifba287889bea3585954fef5efdf5bb24[15][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3eb1902edf9266038f39c281d134c26c[16]        <=  Ifba287889bea3585954fef5efdf5bb24[16][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ifba287889bea3585954fef5efdf5bb24[16] + 1 :
                                             Ifba287889bea3585954fef5efdf5bb24[16] ;
            Ibc0871b3c992fd278815fdbefcd2bac0[16]  <=  Ifba287889bea3585954fef5efdf5bb24[16][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3eb1902edf9266038f39c281d134c26c[17]        <=  Ifba287889bea3585954fef5efdf5bb24[17][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ifba287889bea3585954fef5efdf5bb24[17] + 1 :
                                             Ifba287889bea3585954fef5efdf5bb24[17] ;
            Ibc0871b3c992fd278815fdbefcd2bac0[17]  <=  Ifba287889bea3585954fef5efdf5bb24[17][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3eb1902edf9266038f39c281d134c26c[18]        <=  Ifba287889bea3585954fef5efdf5bb24[18][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ifba287889bea3585954fef5efdf5bb24[18] + 1 :
                                             Ifba287889bea3585954fef5efdf5bb24[18] ;
            Ibc0871b3c992fd278815fdbefcd2bac0[18]  <=  Ifba287889bea3585954fef5efdf5bb24[18][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3eb1902edf9266038f39c281d134c26c[19]        <=  Ifba287889bea3585954fef5efdf5bb24[19][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ifba287889bea3585954fef5efdf5bb24[19] + 1 :
                                             Ifba287889bea3585954fef5efdf5bb24[19] ;
            Ibc0871b3c992fd278815fdbefcd2bac0[19]  <=  Ifba287889bea3585954fef5efdf5bb24[19][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3eb1902edf9266038f39c281d134c26c[20]        <=  Ifba287889bea3585954fef5efdf5bb24[20][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ifba287889bea3585954fef5efdf5bb24[20] + 1 :
                                             Ifba287889bea3585954fef5efdf5bb24[20] ;
            Ibc0871b3c992fd278815fdbefcd2bac0[20]  <=  Ifba287889bea3585954fef5efdf5bb24[20][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3eb1902edf9266038f39c281d134c26c[21]        <=  Ifba287889bea3585954fef5efdf5bb24[21][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ifba287889bea3585954fef5efdf5bb24[21] + 1 :
                                             Ifba287889bea3585954fef5efdf5bb24[21] ;
            Ibc0871b3c992fd278815fdbefcd2bac0[21]  <=  Ifba287889bea3585954fef5efdf5bb24[21][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie791b43e8d5c9d1669743ea4d6e3139c[0]        <=  I8e5ae9e6fa38cea8e5d320fe582c0729[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8e5ae9e6fa38cea8e5d320fe582c0729[0] + 1 :
                                             I8e5ae9e6fa38cea8e5d320fe582c0729[0] ;
            I8695e1e94cbfcbe4b9eae315b042529e[0]  <=  I8e5ae9e6fa38cea8e5d320fe582c0729[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie791b43e8d5c9d1669743ea4d6e3139c[1]        <=  I8e5ae9e6fa38cea8e5d320fe582c0729[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8e5ae9e6fa38cea8e5d320fe582c0729[1] + 1 :
                                             I8e5ae9e6fa38cea8e5d320fe582c0729[1] ;
            I8695e1e94cbfcbe4b9eae315b042529e[1]  <=  I8e5ae9e6fa38cea8e5d320fe582c0729[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie791b43e8d5c9d1669743ea4d6e3139c[2]        <=  I8e5ae9e6fa38cea8e5d320fe582c0729[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8e5ae9e6fa38cea8e5d320fe582c0729[2] + 1 :
                                             I8e5ae9e6fa38cea8e5d320fe582c0729[2] ;
            I8695e1e94cbfcbe4b9eae315b042529e[2]  <=  I8e5ae9e6fa38cea8e5d320fe582c0729[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie791b43e8d5c9d1669743ea4d6e3139c[3]        <=  I8e5ae9e6fa38cea8e5d320fe582c0729[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8e5ae9e6fa38cea8e5d320fe582c0729[3] + 1 :
                                             I8e5ae9e6fa38cea8e5d320fe582c0729[3] ;
            I8695e1e94cbfcbe4b9eae315b042529e[3]  <=  I8e5ae9e6fa38cea8e5d320fe582c0729[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie791b43e8d5c9d1669743ea4d6e3139c[4]        <=  I8e5ae9e6fa38cea8e5d320fe582c0729[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8e5ae9e6fa38cea8e5d320fe582c0729[4] + 1 :
                                             I8e5ae9e6fa38cea8e5d320fe582c0729[4] ;
            I8695e1e94cbfcbe4b9eae315b042529e[4]  <=  I8e5ae9e6fa38cea8e5d320fe582c0729[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie791b43e8d5c9d1669743ea4d6e3139c[5]        <=  I8e5ae9e6fa38cea8e5d320fe582c0729[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8e5ae9e6fa38cea8e5d320fe582c0729[5] + 1 :
                                             I8e5ae9e6fa38cea8e5d320fe582c0729[5] ;
            I8695e1e94cbfcbe4b9eae315b042529e[5]  <=  I8e5ae9e6fa38cea8e5d320fe582c0729[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie791b43e8d5c9d1669743ea4d6e3139c[6]        <=  I8e5ae9e6fa38cea8e5d320fe582c0729[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8e5ae9e6fa38cea8e5d320fe582c0729[6] + 1 :
                                             I8e5ae9e6fa38cea8e5d320fe582c0729[6] ;
            I8695e1e94cbfcbe4b9eae315b042529e[6]  <=  I8e5ae9e6fa38cea8e5d320fe582c0729[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie791b43e8d5c9d1669743ea4d6e3139c[7]        <=  I8e5ae9e6fa38cea8e5d320fe582c0729[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8e5ae9e6fa38cea8e5d320fe582c0729[7] + 1 :
                                             I8e5ae9e6fa38cea8e5d320fe582c0729[7] ;
            I8695e1e94cbfcbe4b9eae315b042529e[7]  <=  I8e5ae9e6fa38cea8e5d320fe582c0729[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie791b43e8d5c9d1669743ea4d6e3139c[8]        <=  I8e5ae9e6fa38cea8e5d320fe582c0729[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8e5ae9e6fa38cea8e5d320fe582c0729[8] + 1 :
                                             I8e5ae9e6fa38cea8e5d320fe582c0729[8] ;
            I8695e1e94cbfcbe4b9eae315b042529e[8]  <=  I8e5ae9e6fa38cea8e5d320fe582c0729[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie791b43e8d5c9d1669743ea4d6e3139c[9]        <=  I8e5ae9e6fa38cea8e5d320fe582c0729[9][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8e5ae9e6fa38cea8e5d320fe582c0729[9] + 1 :
                                             I8e5ae9e6fa38cea8e5d320fe582c0729[9] ;
            I8695e1e94cbfcbe4b9eae315b042529e[9]  <=  I8e5ae9e6fa38cea8e5d320fe582c0729[9][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie791b43e8d5c9d1669743ea4d6e3139c[10]        <=  I8e5ae9e6fa38cea8e5d320fe582c0729[10][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8e5ae9e6fa38cea8e5d320fe582c0729[10] + 1 :
                                             I8e5ae9e6fa38cea8e5d320fe582c0729[10] ;
            I8695e1e94cbfcbe4b9eae315b042529e[10]  <=  I8e5ae9e6fa38cea8e5d320fe582c0729[10][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie791b43e8d5c9d1669743ea4d6e3139c[11]        <=  I8e5ae9e6fa38cea8e5d320fe582c0729[11][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8e5ae9e6fa38cea8e5d320fe582c0729[11] + 1 :
                                             I8e5ae9e6fa38cea8e5d320fe582c0729[11] ;
            I8695e1e94cbfcbe4b9eae315b042529e[11]  <=  I8e5ae9e6fa38cea8e5d320fe582c0729[11][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie791b43e8d5c9d1669743ea4d6e3139c[12]        <=  I8e5ae9e6fa38cea8e5d320fe582c0729[12][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8e5ae9e6fa38cea8e5d320fe582c0729[12] + 1 :
                                             I8e5ae9e6fa38cea8e5d320fe582c0729[12] ;
            I8695e1e94cbfcbe4b9eae315b042529e[12]  <=  I8e5ae9e6fa38cea8e5d320fe582c0729[12][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie791b43e8d5c9d1669743ea4d6e3139c[13]        <=  I8e5ae9e6fa38cea8e5d320fe582c0729[13][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8e5ae9e6fa38cea8e5d320fe582c0729[13] + 1 :
                                             I8e5ae9e6fa38cea8e5d320fe582c0729[13] ;
            I8695e1e94cbfcbe4b9eae315b042529e[13]  <=  I8e5ae9e6fa38cea8e5d320fe582c0729[13][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie791b43e8d5c9d1669743ea4d6e3139c[14]        <=  I8e5ae9e6fa38cea8e5d320fe582c0729[14][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8e5ae9e6fa38cea8e5d320fe582c0729[14] + 1 :
                                             I8e5ae9e6fa38cea8e5d320fe582c0729[14] ;
            I8695e1e94cbfcbe4b9eae315b042529e[14]  <=  I8e5ae9e6fa38cea8e5d320fe582c0729[14][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie791b43e8d5c9d1669743ea4d6e3139c[15]        <=  I8e5ae9e6fa38cea8e5d320fe582c0729[15][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8e5ae9e6fa38cea8e5d320fe582c0729[15] + 1 :
                                             I8e5ae9e6fa38cea8e5d320fe582c0729[15] ;
            I8695e1e94cbfcbe4b9eae315b042529e[15]  <=  I8e5ae9e6fa38cea8e5d320fe582c0729[15][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie791b43e8d5c9d1669743ea4d6e3139c[16]        <=  I8e5ae9e6fa38cea8e5d320fe582c0729[16][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8e5ae9e6fa38cea8e5d320fe582c0729[16] + 1 :
                                             I8e5ae9e6fa38cea8e5d320fe582c0729[16] ;
            I8695e1e94cbfcbe4b9eae315b042529e[16]  <=  I8e5ae9e6fa38cea8e5d320fe582c0729[16][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie791b43e8d5c9d1669743ea4d6e3139c[17]        <=  I8e5ae9e6fa38cea8e5d320fe582c0729[17][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8e5ae9e6fa38cea8e5d320fe582c0729[17] + 1 :
                                             I8e5ae9e6fa38cea8e5d320fe582c0729[17] ;
            I8695e1e94cbfcbe4b9eae315b042529e[17]  <=  I8e5ae9e6fa38cea8e5d320fe582c0729[17][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie791b43e8d5c9d1669743ea4d6e3139c[18]        <=  I8e5ae9e6fa38cea8e5d320fe582c0729[18][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8e5ae9e6fa38cea8e5d320fe582c0729[18] + 1 :
                                             I8e5ae9e6fa38cea8e5d320fe582c0729[18] ;
            I8695e1e94cbfcbe4b9eae315b042529e[18]  <=  I8e5ae9e6fa38cea8e5d320fe582c0729[18][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie791b43e8d5c9d1669743ea4d6e3139c[19]        <=  I8e5ae9e6fa38cea8e5d320fe582c0729[19][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8e5ae9e6fa38cea8e5d320fe582c0729[19] + 1 :
                                             I8e5ae9e6fa38cea8e5d320fe582c0729[19] ;
            I8695e1e94cbfcbe4b9eae315b042529e[19]  <=  I8e5ae9e6fa38cea8e5d320fe582c0729[19][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie791b43e8d5c9d1669743ea4d6e3139c[20]        <=  I8e5ae9e6fa38cea8e5d320fe582c0729[20][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8e5ae9e6fa38cea8e5d320fe582c0729[20] + 1 :
                                             I8e5ae9e6fa38cea8e5d320fe582c0729[20] ;
            I8695e1e94cbfcbe4b9eae315b042529e[20]  <=  I8e5ae9e6fa38cea8e5d320fe582c0729[20][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie791b43e8d5c9d1669743ea4d6e3139c[21]        <=  I8e5ae9e6fa38cea8e5d320fe582c0729[21][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8e5ae9e6fa38cea8e5d320fe582c0729[21] + 1 :
                                             I8e5ae9e6fa38cea8e5d320fe582c0729[21] ;
            I8695e1e94cbfcbe4b9eae315b042529e[21]  <=  I8e5ae9e6fa38cea8e5d320fe582c0729[21][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5b892f00b2642ca102f7755ab512d067[0]        <=  I67315420a608e257df8cfb520ef9f0a1[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I67315420a608e257df8cfb520ef9f0a1[0] + 1 :
                                             I67315420a608e257df8cfb520ef9f0a1[0] ;
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[0]  <=  I67315420a608e257df8cfb520ef9f0a1[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5b892f00b2642ca102f7755ab512d067[1]        <=  I67315420a608e257df8cfb520ef9f0a1[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I67315420a608e257df8cfb520ef9f0a1[1] + 1 :
                                             I67315420a608e257df8cfb520ef9f0a1[1] ;
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[1]  <=  I67315420a608e257df8cfb520ef9f0a1[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5b892f00b2642ca102f7755ab512d067[2]        <=  I67315420a608e257df8cfb520ef9f0a1[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I67315420a608e257df8cfb520ef9f0a1[2] + 1 :
                                             I67315420a608e257df8cfb520ef9f0a1[2] ;
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[2]  <=  I67315420a608e257df8cfb520ef9f0a1[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5b892f00b2642ca102f7755ab512d067[3]        <=  I67315420a608e257df8cfb520ef9f0a1[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I67315420a608e257df8cfb520ef9f0a1[3] + 1 :
                                             I67315420a608e257df8cfb520ef9f0a1[3] ;
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[3]  <=  I67315420a608e257df8cfb520ef9f0a1[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5b892f00b2642ca102f7755ab512d067[4]        <=  I67315420a608e257df8cfb520ef9f0a1[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I67315420a608e257df8cfb520ef9f0a1[4] + 1 :
                                             I67315420a608e257df8cfb520ef9f0a1[4] ;
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[4]  <=  I67315420a608e257df8cfb520ef9f0a1[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5b892f00b2642ca102f7755ab512d067[5]        <=  I67315420a608e257df8cfb520ef9f0a1[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I67315420a608e257df8cfb520ef9f0a1[5] + 1 :
                                             I67315420a608e257df8cfb520ef9f0a1[5] ;
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[5]  <=  I67315420a608e257df8cfb520ef9f0a1[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5b892f00b2642ca102f7755ab512d067[6]        <=  I67315420a608e257df8cfb520ef9f0a1[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I67315420a608e257df8cfb520ef9f0a1[6] + 1 :
                                             I67315420a608e257df8cfb520ef9f0a1[6] ;
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[6]  <=  I67315420a608e257df8cfb520ef9f0a1[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5b892f00b2642ca102f7755ab512d067[7]        <=  I67315420a608e257df8cfb520ef9f0a1[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I67315420a608e257df8cfb520ef9f0a1[7] + 1 :
                                             I67315420a608e257df8cfb520ef9f0a1[7] ;
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[7]  <=  I67315420a608e257df8cfb520ef9f0a1[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5b892f00b2642ca102f7755ab512d067[8]        <=  I67315420a608e257df8cfb520ef9f0a1[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I67315420a608e257df8cfb520ef9f0a1[8] + 1 :
                                             I67315420a608e257df8cfb520ef9f0a1[8] ;
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[8]  <=  I67315420a608e257df8cfb520ef9f0a1[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5b892f00b2642ca102f7755ab512d067[9]        <=  I67315420a608e257df8cfb520ef9f0a1[9][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I67315420a608e257df8cfb520ef9f0a1[9] + 1 :
                                             I67315420a608e257df8cfb520ef9f0a1[9] ;
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[9]  <=  I67315420a608e257df8cfb520ef9f0a1[9][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5b892f00b2642ca102f7755ab512d067[10]        <=  I67315420a608e257df8cfb520ef9f0a1[10][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I67315420a608e257df8cfb520ef9f0a1[10] + 1 :
                                             I67315420a608e257df8cfb520ef9f0a1[10] ;
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[10]  <=  I67315420a608e257df8cfb520ef9f0a1[10][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5b892f00b2642ca102f7755ab512d067[11]        <=  I67315420a608e257df8cfb520ef9f0a1[11][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I67315420a608e257df8cfb520ef9f0a1[11] + 1 :
                                             I67315420a608e257df8cfb520ef9f0a1[11] ;
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[11]  <=  I67315420a608e257df8cfb520ef9f0a1[11][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5b892f00b2642ca102f7755ab512d067[12]        <=  I67315420a608e257df8cfb520ef9f0a1[12][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I67315420a608e257df8cfb520ef9f0a1[12] + 1 :
                                             I67315420a608e257df8cfb520ef9f0a1[12] ;
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[12]  <=  I67315420a608e257df8cfb520ef9f0a1[12][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5b892f00b2642ca102f7755ab512d067[13]        <=  I67315420a608e257df8cfb520ef9f0a1[13][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I67315420a608e257df8cfb520ef9f0a1[13] + 1 :
                                             I67315420a608e257df8cfb520ef9f0a1[13] ;
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[13]  <=  I67315420a608e257df8cfb520ef9f0a1[13][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5b892f00b2642ca102f7755ab512d067[14]        <=  I67315420a608e257df8cfb520ef9f0a1[14][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I67315420a608e257df8cfb520ef9f0a1[14] + 1 :
                                             I67315420a608e257df8cfb520ef9f0a1[14] ;
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[14]  <=  I67315420a608e257df8cfb520ef9f0a1[14][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5b892f00b2642ca102f7755ab512d067[15]        <=  I67315420a608e257df8cfb520ef9f0a1[15][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I67315420a608e257df8cfb520ef9f0a1[15] + 1 :
                                             I67315420a608e257df8cfb520ef9f0a1[15] ;
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[15]  <=  I67315420a608e257df8cfb520ef9f0a1[15][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5b892f00b2642ca102f7755ab512d067[16]        <=  I67315420a608e257df8cfb520ef9f0a1[16][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I67315420a608e257df8cfb520ef9f0a1[16] + 1 :
                                             I67315420a608e257df8cfb520ef9f0a1[16] ;
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[16]  <=  I67315420a608e257df8cfb520ef9f0a1[16][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5b892f00b2642ca102f7755ab512d067[17]        <=  I67315420a608e257df8cfb520ef9f0a1[17][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I67315420a608e257df8cfb520ef9f0a1[17] + 1 :
                                             I67315420a608e257df8cfb520ef9f0a1[17] ;
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[17]  <=  I67315420a608e257df8cfb520ef9f0a1[17][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5b892f00b2642ca102f7755ab512d067[18]        <=  I67315420a608e257df8cfb520ef9f0a1[18][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I67315420a608e257df8cfb520ef9f0a1[18] + 1 :
                                             I67315420a608e257df8cfb520ef9f0a1[18] ;
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[18]  <=  I67315420a608e257df8cfb520ef9f0a1[18][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5b892f00b2642ca102f7755ab512d067[19]        <=  I67315420a608e257df8cfb520ef9f0a1[19][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I67315420a608e257df8cfb520ef9f0a1[19] + 1 :
                                             I67315420a608e257df8cfb520ef9f0a1[19] ;
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[19]  <=  I67315420a608e257df8cfb520ef9f0a1[19][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5b892f00b2642ca102f7755ab512d067[20]        <=  I67315420a608e257df8cfb520ef9f0a1[20][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I67315420a608e257df8cfb520ef9f0a1[20] + 1 :
                                             I67315420a608e257df8cfb520ef9f0a1[20] ;
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[20]  <=  I67315420a608e257df8cfb520ef9f0a1[20][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5b892f00b2642ca102f7755ab512d067[21]        <=  I67315420a608e257df8cfb520ef9f0a1[21][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I67315420a608e257df8cfb520ef9f0a1[21] + 1 :
                                             I67315420a608e257df8cfb520ef9f0a1[21] ;
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[21]  <=  I67315420a608e257df8cfb520ef9f0a1[21][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8f906015dba99b4a73dcf767cbd948ee[0]        <=  Ic80a23c7b47f2236087fd7818d8d7c7f[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic80a23c7b47f2236087fd7818d8d7c7f[0] + 1 :
                                             Ic80a23c7b47f2236087fd7818d8d7c7f[0] ;
            I61f0c04673dfb262ef6912eb2df39120[0]  <=  Ic80a23c7b47f2236087fd7818d8d7c7f[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8f906015dba99b4a73dcf767cbd948ee[1]        <=  Ic80a23c7b47f2236087fd7818d8d7c7f[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic80a23c7b47f2236087fd7818d8d7c7f[1] + 1 :
                                             Ic80a23c7b47f2236087fd7818d8d7c7f[1] ;
            I61f0c04673dfb262ef6912eb2df39120[1]  <=  Ic80a23c7b47f2236087fd7818d8d7c7f[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8f906015dba99b4a73dcf767cbd948ee[2]        <=  Ic80a23c7b47f2236087fd7818d8d7c7f[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic80a23c7b47f2236087fd7818d8d7c7f[2] + 1 :
                                             Ic80a23c7b47f2236087fd7818d8d7c7f[2] ;
            I61f0c04673dfb262ef6912eb2df39120[2]  <=  Ic80a23c7b47f2236087fd7818d8d7c7f[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8f906015dba99b4a73dcf767cbd948ee[3]        <=  Ic80a23c7b47f2236087fd7818d8d7c7f[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic80a23c7b47f2236087fd7818d8d7c7f[3] + 1 :
                                             Ic80a23c7b47f2236087fd7818d8d7c7f[3] ;
            I61f0c04673dfb262ef6912eb2df39120[3]  <=  Ic80a23c7b47f2236087fd7818d8d7c7f[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8f906015dba99b4a73dcf767cbd948ee[4]        <=  Ic80a23c7b47f2236087fd7818d8d7c7f[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic80a23c7b47f2236087fd7818d8d7c7f[4] + 1 :
                                             Ic80a23c7b47f2236087fd7818d8d7c7f[4] ;
            I61f0c04673dfb262ef6912eb2df39120[4]  <=  Ic80a23c7b47f2236087fd7818d8d7c7f[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8f906015dba99b4a73dcf767cbd948ee[5]        <=  Ic80a23c7b47f2236087fd7818d8d7c7f[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic80a23c7b47f2236087fd7818d8d7c7f[5] + 1 :
                                             Ic80a23c7b47f2236087fd7818d8d7c7f[5] ;
            I61f0c04673dfb262ef6912eb2df39120[5]  <=  Ic80a23c7b47f2236087fd7818d8d7c7f[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8f906015dba99b4a73dcf767cbd948ee[6]        <=  Ic80a23c7b47f2236087fd7818d8d7c7f[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic80a23c7b47f2236087fd7818d8d7c7f[6] + 1 :
                                             Ic80a23c7b47f2236087fd7818d8d7c7f[6] ;
            I61f0c04673dfb262ef6912eb2df39120[6]  <=  Ic80a23c7b47f2236087fd7818d8d7c7f[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8f906015dba99b4a73dcf767cbd948ee[7]        <=  Ic80a23c7b47f2236087fd7818d8d7c7f[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic80a23c7b47f2236087fd7818d8d7c7f[7] + 1 :
                                             Ic80a23c7b47f2236087fd7818d8d7c7f[7] ;
            I61f0c04673dfb262ef6912eb2df39120[7]  <=  Ic80a23c7b47f2236087fd7818d8d7c7f[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8f906015dba99b4a73dcf767cbd948ee[8]        <=  Ic80a23c7b47f2236087fd7818d8d7c7f[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic80a23c7b47f2236087fd7818d8d7c7f[8] + 1 :
                                             Ic80a23c7b47f2236087fd7818d8d7c7f[8] ;
            I61f0c04673dfb262ef6912eb2df39120[8]  <=  Ic80a23c7b47f2236087fd7818d8d7c7f[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8f906015dba99b4a73dcf767cbd948ee[9]        <=  Ic80a23c7b47f2236087fd7818d8d7c7f[9][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic80a23c7b47f2236087fd7818d8d7c7f[9] + 1 :
                                             Ic80a23c7b47f2236087fd7818d8d7c7f[9] ;
            I61f0c04673dfb262ef6912eb2df39120[9]  <=  Ic80a23c7b47f2236087fd7818d8d7c7f[9][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8f906015dba99b4a73dcf767cbd948ee[10]        <=  Ic80a23c7b47f2236087fd7818d8d7c7f[10][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic80a23c7b47f2236087fd7818d8d7c7f[10] + 1 :
                                             Ic80a23c7b47f2236087fd7818d8d7c7f[10] ;
            I61f0c04673dfb262ef6912eb2df39120[10]  <=  Ic80a23c7b47f2236087fd7818d8d7c7f[10][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8f906015dba99b4a73dcf767cbd948ee[11]        <=  Ic80a23c7b47f2236087fd7818d8d7c7f[11][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic80a23c7b47f2236087fd7818d8d7c7f[11] + 1 :
                                             Ic80a23c7b47f2236087fd7818d8d7c7f[11] ;
            I61f0c04673dfb262ef6912eb2df39120[11]  <=  Ic80a23c7b47f2236087fd7818d8d7c7f[11][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8f906015dba99b4a73dcf767cbd948ee[12]        <=  Ic80a23c7b47f2236087fd7818d8d7c7f[12][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic80a23c7b47f2236087fd7818d8d7c7f[12] + 1 :
                                             Ic80a23c7b47f2236087fd7818d8d7c7f[12] ;
            I61f0c04673dfb262ef6912eb2df39120[12]  <=  Ic80a23c7b47f2236087fd7818d8d7c7f[12][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8f906015dba99b4a73dcf767cbd948ee[13]        <=  Ic80a23c7b47f2236087fd7818d8d7c7f[13][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic80a23c7b47f2236087fd7818d8d7c7f[13] + 1 :
                                             Ic80a23c7b47f2236087fd7818d8d7c7f[13] ;
            I61f0c04673dfb262ef6912eb2df39120[13]  <=  Ic80a23c7b47f2236087fd7818d8d7c7f[13][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8f906015dba99b4a73dcf767cbd948ee[14]        <=  Ic80a23c7b47f2236087fd7818d8d7c7f[14][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic80a23c7b47f2236087fd7818d8d7c7f[14] + 1 :
                                             Ic80a23c7b47f2236087fd7818d8d7c7f[14] ;
            I61f0c04673dfb262ef6912eb2df39120[14]  <=  Ic80a23c7b47f2236087fd7818d8d7c7f[14][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8f906015dba99b4a73dcf767cbd948ee[15]        <=  Ic80a23c7b47f2236087fd7818d8d7c7f[15][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic80a23c7b47f2236087fd7818d8d7c7f[15] + 1 :
                                             Ic80a23c7b47f2236087fd7818d8d7c7f[15] ;
            I61f0c04673dfb262ef6912eb2df39120[15]  <=  Ic80a23c7b47f2236087fd7818d8d7c7f[15][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8f906015dba99b4a73dcf767cbd948ee[16]        <=  Ic80a23c7b47f2236087fd7818d8d7c7f[16][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic80a23c7b47f2236087fd7818d8d7c7f[16] + 1 :
                                             Ic80a23c7b47f2236087fd7818d8d7c7f[16] ;
            I61f0c04673dfb262ef6912eb2df39120[16]  <=  Ic80a23c7b47f2236087fd7818d8d7c7f[16][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8f906015dba99b4a73dcf767cbd948ee[17]        <=  Ic80a23c7b47f2236087fd7818d8d7c7f[17][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic80a23c7b47f2236087fd7818d8d7c7f[17] + 1 :
                                             Ic80a23c7b47f2236087fd7818d8d7c7f[17] ;
            I61f0c04673dfb262ef6912eb2df39120[17]  <=  Ic80a23c7b47f2236087fd7818d8d7c7f[17][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8f906015dba99b4a73dcf767cbd948ee[18]        <=  Ic80a23c7b47f2236087fd7818d8d7c7f[18][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic80a23c7b47f2236087fd7818d8d7c7f[18] + 1 :
                                             Ic80a23c7b47f2236087fd7818d8d7c7f[18] ;
            I61f0c04673dfb262ef6912eb2df39120[18]  <=  Ic80a23c7b47f2236087fd7818d8d7c7f[18][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8f906015dba99b4a73dcf767cbd948ee[19]        <=  Ic80a23c7b47f2236087fd7818d8d7c7f[19][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic80a23c7b47f2236087fd7818d8d7c7f[19] + 1 :
                                             Ic80a23c7b47f2236087fd7818d8d7c7f[19] ;
            I61f0c04673dfb262ef6912eb2df39120[19]  <=  Ic80a23c7b47f2236087fd7818d8d7c7f[19][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8f906015dba99b4a73dcf767cbd948ee[20]        <=  Ic80a23c7b47f2236087fd7818d8d7c7f[20][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic80a23c7b47f2236087fd7818d8d7c7f[20] + 1 :
                                             Ic80a23c7b47f2236087fd7818d8d7c7f[20] ;
            I61f0c04673dfb262ef6912eb2df39120[20]  <=  Ic80a23c7b47f2236087fd7818d8d7c7f[20][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8f906015dba99b4a73dcf767cbd948ee[21]        <=  Ic80a23c7b47f2236087fd7818d8d7c7f[21][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic80a23c7b47f2236087fd7818d8d7c7f[21] + 1 :
                                             Ic80a23c7b47f2236087fd7818d8d7c7f[21] ;
            I61f0c04673dfb262ef6912eb2df39120[21]  <=  Ic80a23c7b47f2236087fd7818d8d7c7f[21][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8f906015dba99b4a73dcf767cbd948ee[22]        <=  Ic80a23c7b47f2236087fd7818d8d7c7f[22][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic80a23c7b47f2236087fd7818d8d7c7f[22] + 1 :
                                             Ic80a23c7b47f2236087fd7818d8d7c7f[22] ;
            I61f0c04673dfb262ef6912eb2df39120[22]  <=  Ic80a23c7b47f2236087fd7818d8d7c7f[22][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9ab4bbe4191d0f284defcdce6b885054[0]        <=  Ie53d62e3ef9caf35092d7a63be1f565f[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie53d62e3ef9caf35092d7a63be1f565f[0] + 1 :
                                             Ie53d62e3ef9caf35092d7a63be1f565f[0] ;
            Ibeb5edab51cd6aedad9c2ecedaded6f5[0]  <=  Ie53d62e3ef9caf35092d7a63be1f565f[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9ab4bbe4191d0f284defcdce6b885054[1]        <=  Ie53d62e3ef9caf35092d7a63be1f565f[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie53d62e3ef9caf35092d7a63be1f565f[1] + 1 :
                                             Ie53d62e3ef9caf35092d7a63be1f565f[1] ;
            Ibeb5edab51cd6aedad9c2ecedaded6f5[1]  <=  Ie53d62e3ef9caf35092d7a63be1f565f[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9ab4bbe4191d0f284defcdce6b885054[2]        <=  Ie53d62e3ef9caf35092d7a63be1f565f[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie53d62e3ef9caf35092d7a63be1f565f[2] + 1 :
                                             Ie53d62e3ef9caf35092d7a63be1f565f[2] ;
            Ibeb5edab51cd6aedad9c2ecedaded6f5[2]  <=  Ie53d62e3ef9caf35092d7a63be1f565f[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9ab4bbe4191d0f284defcdce6b885054[3]        <=  Ie53d62e3ef9caf35092d7a63be1f565f[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie53d62e3ef9caf35092d7a63be1f565f[3] + 1 :
                                             Ie53d62e3ef9caf35092d7a63be1f565f[3] ;
            Ibeb5edab51cd6aedad9c2ecedaded6f5[3]  <=  Ie53d62e3ef9caf35092d7a63be1f565f[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9ab4bbe4191d0f284defcdce6b885054[4]        <=  Ie53d62e3ef9caf35092d7a63be1f565f[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie53d62e3ef9caf35092d7a63be1f565f[4] + 1 :
                                             Ie53d62e3ef9caf35092d7a63be1f565f[4] ;
            Ibeb5edab51cd6aedad9c2ecedaded6f5[4]  <=  Ie53d62e3ef9caf35092d7a63be1f565f[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9ab4bbe4191d0f284defcdce6b885054[5]        <=  Ie53d62e3ef9caf35092d7a63be1f565f[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie53d62e3ef9caf35092d7a63be1f565f[5] + 1 :
                                             Ie53d62e3ef9caf35092d7a63be1f565f[5] ;
            Ibeb5edab51cd6aedad9c2ecedaded6f5[5]  <=  Ie53d62e3ef9caf35092d7a63be1f565f[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9ab4bbe4191d0f284defcdce6b885054[6]        <=  Ie53d62e3ef9caf35092d7a63be1f565f[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie53d62e3ef9caf35092d7a63be1f565f[6] + 1 :
                                             Ie53d62e3ef9caf35092d7a63be1f565f[6] ;
            Ibeb5edab51cd6aedad9c2ecedaded6f5[6]  <=  Ie53d62e3ef9caf35092d7a63be1f565f[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9ab4bbe4191d0f284defcdce6b885054[7]        <=  Ie53d62e3ef9caf35092d7a63be1f565f[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie53d62e3ef9caf35092d7a63be1f565f[7] + 1 :
                                             Ie53d62e3ef9caf35092d7a63be1f565f[7] ;
            Ibeb5edab51cd6aedad9c2ecedaded6f5[7]  <=  Ie53d62e3ef9caf35092d7a63be1f565f[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9ab4bbe4191d0f284defcdce6b885054[8]        <=  Ie53d62e3ef9caf35092d7a63be1f565f[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie53d62e3ef9caf35092d7a63be1f565f[8] + 1 :
                                             Ie53d62e3ef9caf35092d7a63be1f565f[8] ;
            Ibeb5edab51cd6aedad9c2ecedaded6f5[8]  <=  Ie53d62e3ef9caf35092d7a63be1f565f[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9ab4bbe4191d0f284defcdce6b885054[9]        <=  Ie53d62e3ef9caf35092d7a63be1f565f[9][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie53d62e3ef9caf35092d7a63be1f565f[9] + 1 :
                                             Ie53d62e3ef9caf35092d7a63be1f565f[9] ;
            Ibeb5edab51cd6aedad9c2ecedaded6f5[9]  <=  Ie53d62e3ef9caf35092d7a63be1f565f[9][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9ab4bbe4191d0f284defcdce6b885054[10]        <=  Ie53d62e3ef9caf35092d7a63be1f565f[10][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie53d62e3ef9caf35092d7a63be1f565f[10] + 1 :
                                             Ie53d62e3ef9caf35092d7a63be1f565f[10] ;
            Ibeb5edab51cd6aedad9c2ecedaded6f5[10]  <=  Ie53d62e3ef9caf35092d7a63be1f565f[10][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9ab4bbe4191d0f284defcdce6b885054[11]        <=  Ie53d62e3ef9caf35092d7a63be1f565f[11][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie53d62e3ef9caf35092d7a63be1f565f[11] + 1 :
                                             Ie53d62e3ef9caf35092d7a63be1f565f[11] ;
            Ibeb5edab51cd6aedad9c2ecedaded6f5[11]  <=  Ie53d62e3ef9caf35092d7a63be1f565f[11][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9ab4bbe4191d0f284defcdce6b885054[12]        <=  Ie53d62e3ef9caf35092d7a63be1f565f[12][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie53d62e3ef9caf35092d7a63be1f565f[12] + 1 :
                                             Ie53d62e3ef9caf35092d7a63be1f565f[12] ;
            Ibeb5edab51cd6aedad9c2ecedaded6f5[12]  <=  Ie53d62e3ef9caf35092d7a63be1f565f[12][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9ab4bbe4191d0f284defcdce6b885054[13]        <=  Ie53d62e3ef9caf35092d7a63be1f565f[13][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie53d62e3ef9caf35092d7a63be1f565f[13] + 1 :
                                             Ie53d62e3ef9caf35092d7a63be1f565f[13] ;
            Ibeb5edab51cd6aedad9c2ecedaded6f5[13]  <=  Ie53d62e3ef9caf35092d7a63be1f565f[13][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9ab4bbe4191d0f284defcdce6b885054[14]        <=  Ie53d62e3ef9caf35092d7a63be1f565f[14][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie53d62e3ef9caf35092d7a63be1f565f[14] + 1 :
                                             Ie53d62e3ef9caf35092d7a63be1f565f[14] ;
            Ibeb5edab51cd6aedad9c2ecedaded6f5[14]  <=  Ie53d62e3ef9caf35092d7a63be1f565f[14][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9ab4bbe4191d0f284defcdce6b885054[15]        <=  Ie53d62e3ef9caf35092d7a63be1f565f[15][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie53d62e3ef9caf35092d7a63be1f565f[15] + 1 :
                                             Ie53d62e3ef9caf35092d7a63be1f565f[15] ;
            Ibeb5edab51cd6aedad9c2ecedaded6f5[15]  <=  Ie53d62e3ef9caf35092d7a63be1f565f[15][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9ab4bbe4191d0f284defcdce6b885054[16]        <=  Ie53d62e3ef9caf35092d7a63be1f565f[16][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie53d62e3ef9caf35092d7a63be1f565f[16] + 1 :
                                             Ie53d62e3ef9caf35092d7a63be1f565f[16] ;
            Ibeb5edab51cd6aedad9c2ecedaded6f5[16]  <=  Ie53d62e3ef9caf35092d7a63be1f565f[16][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9ab4bbe4191d0f284defcdce6b885054[17]        <=  Ie53d62e3ef9caf35092d7a63be1f565f[17][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie53d62e3ef9caf35092d7a63be1f565f[17] + 1 :
                                             Ie53d62e3ef9caf35092d7a63be1f565f[17] ;
            Ibeb5edab51cd6aedad9c2ecedaded6f5[17]  <=  Ie53d62e3ef9caf35092d7a63be1f565f[17][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9ab4bbe4191d0f284defcdce6b885054[18]        <=  Ie53d62e3ef9caf35092d7a63be1f565f[18][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie53d62e3ef9caf35092d7a63be1f565f[18] + 1 :
                                             Ie53d62e3ef9caf35092d7a63be1f565f[18] ;
            Ibeb5edab51cd6aedad9c2ecedaded6f5[18]  <=  Ie53d62e3ef9caf35092d7a63be1f565f[18][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9ab4bbe4191d0f284defcdce6b885054[19]        <=  Ie53d62e3ef9caf35092d7a63be1f565f[19][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie53d62e3ef9caf35092d7a63be1f565f[19] + 1 :
                                             Ie53d62e3ef9caf35092d7a63be1f565f[19] ;
            Ibeb5edab51cd6aedad9c2ecedaded6f5[19]  <=  Ie53d62e3ef9caf35092d7a63be1f565f[19][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9ab4bbe4191d0f284defcdce6b885054[20]        <=  Ie53d62e3ef9caf35092d7a63be1f565f[20][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie53d62e3ef9caf35092d7a63be1f565f[20] + 1 :
                                             Ie53d62e3ef9caf35092d7a63be1f565f[20] ;
            Ibeb5edab51cd6aedad9c2ecedaded6f5[20]  <=  Ie53d62e3ef9caf35092d7a63be1f565f[20][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9ab4bbe4191d0f284defcdce6b885054[21]        <=  Ie53d62e3ef9caf35092d7a63be1f565f[21][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie53d62e3ef9caf35092d7a63be1f565f[21] + 1 :
                                             Ie53d62e3ef9caf35092d7a63be1f565f[21] ;
            Ibeb5edab51cd6aedad9c2ecedaded6f5[21]  <=  Ie53d62e3ef9caf35092d7a63be1f565f[21][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9ab4bbe4191d0f284defcdce6b885054[22]        <=  Ie53d62e3ef9caf35092d7a63be1f565f[22][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie53d62e3ef9caf35092d7a63be1f565f[22] + 1 :
                                             Ie53d62e3ef9caf35092d7a63be1f565f[22] ;
            Ibeb5edab51cd6aedad9c2ecedaded6f5[22]  <=  Ie53d62e3ef9caf35092d7a63be1f565f[22][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[0]        <=  Ia73bc9712b861f909d0e3683ec91ea1c[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia73bc9712b861f909d0e3683ec91ea1c[0] + 1 :
                                             Ia73bc9712b861f909d0e3683ec91ea1c[0] ;
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[0]  <=  Ia73bc9712b861f909d0e3683ec91ea1c[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[1]        <=  Ia73bc9712b861f909d0e3683ec91ea1c[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia73bc9712b861f909d0e3683ec91ea1c[1] + 1 :
                                             Ia73bc9712b861f909d0e3683ec91ea1c[1] ;
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[1]  <=  Ia73bc9712b861f909d0e3683ec91ea1c[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[2]        <=  Ia73bc9712b861f909d0e3683ec91ea1c[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia73bc9712b861f909d0e3683ec91ea1c[2] + 1 :
                                             Ia73bc9712b861f909d0e3683ec91ea1c[2] ;
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[2]  <=  Ia73bc9712b861f909d0e3683ec91ea1c[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[3]        <=  Ia73bc9712b861f909d0e3683ec91ea1c[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia73bc9712b861f909d0e3683ec91ea1c[3] + 1 :
                                             Ia73bc9712b861f909d0e3683ec91ea1c[3] ;
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[3]  <=  Ia73bc9712b861f909d0e3683ec91ea1c[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[4]        <=  Ia73bc9712b861f909d0e3683ec91ea1c[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia73bc9712b861f909d0e3683ec91ea1c[4] + 1 :
                                             Ia73bc9712b861f909d0e3683ec91ea1c[4] ;
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[4]  <=  Ia73bc9712b861f909d0e3683ec91ea1c[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[5]        <=  Ia73bc9712b861f909d0e3683ec91ea1c[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia73bc9712b861f909d0e3683ec91ea1c[5] + 1 :
                                             Ia73bc9712b861f909d0e3683ec91ea1c[5] ;
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[5]  <=  Ia73bc9712b861f909d0e3683ec91ea1c[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[6]        <=  Ia73bc9712b861f909d0e3683ec91ea1c[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia73bc9712b861f909d0e3683ec91ea1c[6] + 1 :
                                             Ia73bc9712b861f909d0e3683ec91ea1c[6] ;
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[6]  <=  Ia73bc9712b861f909d0e3683ec91ea1c[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[7]        <=  Ia73bc9712b861f909d0e3683ec91ea1c[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia73bc9712b861f909d0e3683ec91ea1c[7] + 1 :
                                             Ia73bc9712b861f909d0e3683ec91ea1c[7] ;
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[7]  <=  Ia73bc9712b861f909d0e3683ec91ea1c[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[8]        <=  Ia73bc9712b861f909d0e3683ec91ea1c[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia73bc9712b861f909d0e3683ec91ea1c[8] + 1 :
                                             Ia73bc9712b861f909d0e3683ec91ea1c[8] ;
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[8]  <=  Ia73bc9712b861f909d0e3683ec91ea1c[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[9]        <=  Ia73bc9712b861f909d0e3683ec91ea1c[9][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia73bc9712b861f909d0e3683ec91ea1c[9] + 1 :
                                             Ia73bc9712b861f909d0e3683ec91ea1c[9] ;
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[9]  <=  Ia73bc9712b861f909d0e3683ec91ea1c[9][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[10]        <=  Ia73bc9712b861f909d0e3683ec91ea1c[10][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia73bc9712b861f909d0e3683ec91ea1c[10] + 1 :
                                             Ia73bc9712b861f909d0e3683ec91ea1c[10] ;
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[10]  <=  Ia73bc9712b861f909d0e3683ec91ea1c[10][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[11]        <=  Ia73bc9712b861f909d0e3683ec91ea1c[11][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia73bc9712b861f909d0e3683ec91ea1c[11] + 1 :
                                             Ia73bc9712b861f909d0e3683ec91ea1c[11] ;
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[11]  <=  Ia73bc9712b861f909d0e3683ec91ea1c[11][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[12]        <=  Ia73bc9712b861f909d0e3683ec91ea1c[12][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia73bc9712b861f909d0e3683ec91ea1c[12] + 1 :
                                             Ia73bc9712b861f909d0e3683ec91ea1c[12] ;
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[12]  <=  Ia73bc9712b861f909d0e3683ec91ea1c[12][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[13]        <=  Ia73bc9712b861f909d0e3683ec91ea1c[13][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia73bc9712b861f909d0e3683ec91ea1c[13] + 1 :
                                             Ia73bc9712b861f909d0e3683ec91ea1c[13] ;
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[13]  <=  Ia73bc9712b861f909d0e3683ec91ea1c[13][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[14]        <=  Ia73bc9712b861f909d0e3683ec91ea1c[14][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia73bc9712b861f909d0e3683ec91ea1c[14] + 1 :
                                             Ia73bc9712b861f909d0e3683ec91ea1c[14] ;
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[14]  <=  Ia73bc9712b861f909d0e3683ec91ea1c[14][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[15]        <=  Ia73bc9712b861f909d0e3683ec91ea1c[15][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia73bc9712b861f909d0e3683ec91ea1c[15] + 1 :
                                             Ia73bc9712b861f909d0e3683ec91ea1c[15] ;
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[15]  <=  Ia73bc9712b861f909d0e3683ec91ea1c[15][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[16]        <=  Ia73bc9712b861f909d0e3683ec91ea1c[16][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia73bc9712b861f909d0e3683ec91ea1c[16] + 1 :
                                             Ia73bc9712b861f909d0e3683ec91ea1c[16] ;
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[16]  <=  Ia73bc9712b861f909d0e3683ec91ea1c[16][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[17]        <=  Ia73bc9712b861f909d0e3683ec91ea1c[17][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia73bc9712b861f909d0e3683ec91ea1c[17] + 1 :
                                             Ia73bc9712b861f909d0e3683ec91ea1c[17] ;
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[17]  <=  Ia73bc9712b861f909d0e3683ec91ea1c[17][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[18]        <=  Ia73bc9712b861f909d0e3683ec91ea1c[18][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia73bc9712b861f909d0e3683ec91ea1c[18] + 1 :
                                             Ia73bc9712b861f909d0e3683ec91ea1c[18] ;
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[18]  <=  Ia73bc9712b861f909d0e3683ec91ea1c[18][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[19]        <=  Ia73bc9712b861f909d0e3683ec91ea1c[19][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia73bc9712b861f909d0e3683ec91ea1c[19] + 1 :
                                             Ia73bc9712b861f909d0e3683ec91ea1c[19] ;
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[19]  <=  Ia73bc9712b861f909d0e3683ec91ea1c[19][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[20]        <=  Ia73bc9712b861f909d0e3683ec91ea1c[20][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia73bc9712b861f909d0e3683ec91ea1c[20] + 1 :
                                             Ia73bc9712b861f909d0e3683ec91ea1c[20] ;
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[20]  <=  Ia73bc9712b861f909d0e3683ec91ea1c[20][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[21]        <=  Ia73bc9712b861f909d0e3683ec91ea1c[21][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia73bc9712b861f909d0e3683ec91ea1c[21] + 1 :
                                             Ia73bc9712b861f909d0e3683ec91ea1c[21] ;
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[21]  <=  Ia73bc9712b861f909d0e3683ec91ea1c[21][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic8a3b3e2aacd0eb24cbc429e9bb734ee[22]        <=  Ia73bc9712b861f909d0e3683ec91ea1c[22][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia73bc9712b861f909d0e3683ec91ea1c[22] + 1 :
                                             Ia73bc9712b861f909d0e3683ec91ea1c[22] ;
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[22]  <=  Ia73bc9712b861f909d0e3683ec91ea1c[22][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6ff6fafd1a3364131b269724ad273ba5[0]        <=  I97d2ee9c3120e78ebcda2f0dbb888b49[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I97d2ee9c3120e78ebcda2f0dbb888b49[0] + 1 :
                                             I97d2ee9c3120e78ebcda2f0dbb888b49[0] ;
            I5b7caaeb34c43e66e8d095a859e708fe[0]  <=  I97d2ee9c3120e78ebcda2f0dbb888b49[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6ff6fafd1a3364131b269724ad273ba5[1]        <=  I97d2ee9c3120e78ebcda2f0dbb888b49[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I97d2ee9c3120e78ebcda2f0dbb888b49[1] + 1 :
                                             I97d2ee9c3120e78ebcda2f0dbb888b49[1] ;
            I5b7caaeb34c43e66e8d095a859e708fe[1]  <=  I97d2ee9c3120e78ebcda2f0dbb888b49[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6ff6fafd1a3364131b269724ad273ba5[2]        <=  I97d2ee9c3120e78ebcda2f0dbb888b49[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I97d2ee9c3120e78ebcda2f0dbb888b49[2] + 1 :
                                             I97d2ee9c3120e78ebcda2f0dbb888b49[2] ;
            I5b7caaeb34c43e66e8d095a859e708fe[2]  <=  I97d2ee9c3120e78ebcda2f0dbb888b49[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6ff6fafd1a3364131b269724ad273ba5[3]        <=  I97d2ee9c3120e78ebcda2f0dbb888b49[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I97d2ee9c3120e78ebcda2f0dbb888b49[3] + 1 :
                                             I97d2ee9c3120e78ebcda2f0dbb888b49[3] ;
            I5b7caaeb34c43e66e8d095a859e708fe[3]  <=  I97d2ee9c3120e78ebcda2f0dbb888b49[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6ff6fafd1a3364131b269724ad273ba5[4]        <=  I97d2ee9c3120e78ebcda2f0dbb888b49[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I97d2ee9c3120e78ebcda2f0dbb888b49[4] + 1 :
                                             I97d2ee9c3120e78ebcda2f0dbb888b49[4] ;
            I5b7caaeb34c43e66e8d095a859e708fe[4]  <=  I97d2ee9c3120e78ebcda2f0dbb888b49[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6ff6fafd1a3364131b269724ad273ba5[5]        <=  I97d2ee9c3120e78ebcda2f0dbb888b49[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I97d2ee9c3120e78ebcda2f0dbb888b49[5] + 1 :
                                             I97d2ee9c3120e78ebcda2f0dbb888b49[5] ;
            I5b7caaeb34c43e66e8d095a859e708fe[5]  <=  I97d2ee9c3120e78ebcda2f0dbb888b49[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6ff6fafd1a3364131b269724ad273ba5[6]        <=  I97d2ee9c3120e78ebcda2f0dbb888b49[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I97d2ee9c3120e78ebcda2f0dbb888b49[6] + 1 :
                                             I97d2ee9c3120e78ebcda2f0dbb888b49[6] ;
            I5b7caaeb34c43e66e8d095a859e708fe[6]  <=  I97d2ee9c3120e78ebcda2f0dbb888b49[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6ff6fafd1a3364131b269724ad273ba5[7]        <=  I97d2ee9c3120e78ebcda2f0dbb888b49[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I97d2ee9c3120e78ebcda2f0dbb888b49[7] + 1 :
                                             I97d2ee9c3120e78ebcda2f0dbb888b49[7] ;
            I5b7caaeb34c43e66e8d095a859e708fe[7]  <=  I97d2ee9c3120e78ebcda2f0dbb888b49[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6ff6fafd1a3364131b269724ad273ba5[8]        <=  I97d2ee9c3120e78ebcda2f0dbb888b49[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I97d2ee9c3120e78ebcda2f0dbb888b49[8] + 1 :
                                             I97d2ee9c3120e78ebcda2f0dbb888b49[8] ;
            I5b7caaeb34c43e66e8d095a859e708fe[8]  <=  I97d2ee9c3120e78ebcda2f0dbb888b49[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6ff6fafd1a3364131b269724ad273ba5[9]        <=  I97d2ee9c3120e78ebcda2f0dbb888b49[9][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I97d2ee9c3120e78ebcda2f0dbb888b49[9] + 1 :
                                             I97d2ee9c3120e78ebcda2f0dbb888b49[9] ;
            I5b7caaeb34c43e66e8d095a859e708fe[9]  <=  I97d2ee9c3120e78ebcda2f0dbb888b49[9][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6ff6fafd1a3364131b269724ad273ba5[10]        <=  I97d2ee9c3120e78ebcda2f0dbb888b49[10][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I97d2ee9c3120e78ebcda2f0dbb888b49[10] + 1 :
                                             I97d2ee9c3120e78ebcda2f0dbb888b49[10] ;
            I5b7caaeb34c43e66e8d095a859e708fe[10]  <=  I97d2ee9c3120e78ebcda2f0dbb888b49[10][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6ff6fafd1a3364131b269724ad273ba5[11]        <=  I97d2ee9c3120e78ebcda2f0dbb888b49[11][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I97d2ee9c3120e78ebcda2f0dbb888b49[11] + 1 :
                                             I97d2ee9c3120e78ebcda2f0dbb888b49[11] ;
            I5b7caaeb34c43e66e8d095a859e708fe[11]  <=  I97d2ee9c3120e78ebcda2f0dbb888b49[11][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6ff6fafd1a3364131b269724ad273ba5[12]        <=  I97d2ee9c3120e78ebcda2f0dbb888b49[12][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I97d2ee9c3120e78ebcda2f0dbb888b49[12] + 1 :
                                             I97d2ee9c3120e78ebcda2f0dbb888b49[12] ;
            I5b7caaeb34c43e66e8d095a859e708fe[12]  <=  I97d2ee9c3120e78ebcda2f0dbb888b49[12][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6ff6fafd1a3364131b269724ad273ba5[13]        <=  I97d2ee9c3120e78ebcda2f0dbb888b49[13][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I97d2ee9c3120e78ebcda2f0dbb888b49[13] + 1 :
                                             I97d2ee9c3120e78ebcda2f0dbb888b49[13] ;
            I5b7caaeb34c43e66e8d095a859e708fe[13]  <=  I97d2ee9c3120e78ebcda2f0dbb888b49[13][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6ff6fafd1a3364131b269724ad273ba5[14]        <=  I97d2ee9c3120e78ebcda2f0dbb888b49[14][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I97d2ee9c3120e78ebcda2f0dbb888b49[14] + 1 :
                                             I97d2ee9c3120e78ebcda2f0dbb888b49[14] ;
            I5b7caaeb34c43e66e8d095a859e708fe[14]  <=  I97d2ee9c3120e78ebcda2f0dbb888b49[14][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6ff6fafd1a3364131b269724ad273ba5[15]        <=  I97d2ee9c3120e78ebcda2f0dbb888b49[15][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I97d2ee9c3120e78ebcda2f0dbb888b49[15] + 1 :
                                             I97d2ee9c3120e78ebcda2f0dbb888b49[15] ;
            I5b7caaeb34c43e66e8d095a859e708fe[15]  <=  I97d2ee9c3120e78ebcda2f0dbb888b49[15][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6ff6fafd1a3364131b269724ad273ba5[16]        <=  I97d2ee9c3120e78ebcda2f0dbb888b49[16][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I97d2ee9c3120e78ebcda2f0dbb888b49[16] + 1 :
                                             I97d2ee9c3120e78ebcda2f0dbb888b49[16] ;
            I5b7caaeb34c43e66e8d095a859e708fe[16]  <=  I97d2ee9c3120e78ebcda2f0dbb888b49[16][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6ff6fafd1a3364131b269724ad273ba5[17]        <=  I97d2ee9c3120e78ebcda2f0dbb888b49[17][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I97d2ee9c3120e78ebcda2f0dbb888b49[17] + 1 :
                                             I97d2ee9c3120e78ebcda2f0dbb888b49[17] ;
            I5b7caaeb34c43e66e8d095a859e708fe[17]  <=  I97d2ee9c3120e78ebcda2f0dbb888b49[17][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6ff6fafd1a3364131b269724ad273ba5[18]        <=  I97d2ee9c3120e78ebcda2f0dbb888b49[18][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I97d2ee9c3120e78ebcda2f0dbb888b49[18] + 1 :
                                             I97d2ee9c3120e78ebcda2f0dbb888b49[18] ;
            I5b7caaeb34c43e66e8d095a859e708fe[18]  <=  I97d2ee9c3120e78ebcda2f0dbb888b49[18][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6ff6fafd1a3364131b269724ad273ba5[19]        <=  I97d2ee9c3120e78ebcda2f0dbb888b49[19][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I97d2ee9c3120e78ebcda2f0dbb888b49[19] + 1 :
                                             I97d2ee9c3120e78ebcda2f0dbb888b49[19] ;
            I5b7caaeb34c43e66e8d095a859e708fe[19]  <=  I97d2ee9c3120e78ebcda2f0dbb888b49[19][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6ff6fafd1a3364131b269724ad273ba5[20]        <=  I97d2ee9c3120e78ebcda2f0dbb888b49[20][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I97d2ee9c3120e78ebcda2f0dbb888b49[20] + 1 :
                                             I97d2ee9c3120e78ebcda2f0dbb888b49[20] ;
            I5b7caaeb34c43e66e8d095a859e708fe[20]  <=  I97d2ee9c3120e78ebcda2f0dbb888b49[20][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6ff6fafd1a3364131b269724ad273ba5[21]        <=  I97d2ee9c3120e78ebcda2f0dbb888b49[21][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I97d2ee9c3120e78ebcda2f0dbb888b49[21] + 1 :
                                             I97d2ee9c3120e78ebcda2f0dbb888b49[21] ;
            I5b7caaeb34c43e66e8d095a859e708fe[21]  <=  I97d2ee9c3120e78ebcda2f0dbb888b49[21][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6ff6fafd1a3364131b269724ad273ba5[22]        <=  I97d2ee9c3120e78ebcda2f0dbb888b49[22][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I97d2ee9c3120e78ebcda2f0dbb888b49[22] + 1 :
                                             I97d2ee9c3120e78ebcda2f0dbb888b49[22] ;
            I5b7caaeb34c43e66e8d095a859e708fe[22]  <=  I97d2ee9c3120e78ebcda2f0dbb888b49[22][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I154fcd3171f1231e825ee603d53ecfe8[0]        <=  I07b2a00225c337eed1e5a350f3361240[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I07b2a00225c337eed1e5a350f3361240[0] + 1 :
                                             I07b2a00225c337eed1e5a350f3361240[0] ;
            Ib0bf69cc797f330fb2546eb46d2d6f76[0]  <=  I07b2a00225c337eed1e5a350f3361240[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I154fcd3171f1231e825ee603d53ecfe8[1]        <=  I07b2a00225c337eed1e5a350f3361240[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I07b2a00225c337eed1e5a350f3361240[1] + 1 :
                                             I07b2a00225c337eed1e5a350f3361240[1] ;
            Ib0bf69cc797f330fb2546eb46d2d6f76[1]  <=  I07b2a00225c337eed1e5a350f3361240[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I154fcd3171f1231e825ee603d53ecfe8[2]        <=  I07b2a00225c337eed1e5a350f3361240[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I07b2a00225c337eed1e5a350f3361240[2] + 1 :
                                             I07b2a00225c337eed1e5a350f3361240[2] ;
            Ib0bf69cc797f330fb2546eb46d2d6f76[2]  <=  I07b2a00225c337eed1e5a350f3361240[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I154fcd3171f1231e825ee603d53ecfe8[3]        <=  I07b2a00225c337eed1e5a350f3361240[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I07b2a00225c337eed1e5a350f3361240[3] + 1 :
                                             I07b2a00225c337eed1e5a350f3361240[3] ;
            Ib0bf69cc797f330fb2546eb46d2d6f76[3]  <=  I07b2a00225c337eed1e5a350f3361240[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I154fcd3171f1231e825ee603d53ecfe8[4]        <=  I07b2a00225c337eed1e5a350f3361240[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I07b2a00225c337eed1e5a350f3361240[4] + 1 :
                                             I07b2a00225c337eed1e5a350f3361240[4] ;
            Ib0bf69cc797f330fb2546eb46d2d6f76[4]  <=  I07b2a00225c337eed1e5a350f3361240[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I154fcd3171f1231e825ee603d53ecfe8[5]        <=  I07b2a00225c337eed1e5a350f3361240[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I07b2a00225c337eed1e5a350f3361240[5] + 1 :
                                             I07b2a00225c337eed1e5a350f3361240[5] ;
            Ib0bf69cc797f330fb2546eb46d2d6f76[5]  <=  I07b2a00225c337eed1e5a350f3361240[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I154fcd3171f1231e825ee603d53ecfe8[6]        <=  I07b2a00225c337eed1e5a350f3361240[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I07b2a00225c337eed1e5a350f3361240[6] + 1 :
                                             I07b2a00225c337eed1e5a350f3361240[6] ;
            Ib0bf69cc797f330fb2546eb46d2d6f76[6]  <=  I07b2a00225c337eed1e5a350f3361240[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I154fcd3171f1231e825ee603d53ecfe8[7]        <=  I07b2a00225c337eed1e5a350f3361240[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I07b2a00225c337eed1e5a350f3361240[7] + 1 :
                                             I07b2a00225c337eed1e5a350f3361240[7] ;
            Ib0bf69cc797f330fb2546eb46d2d6f76[7]  <=  I07b2a00225c337eed1e5a350f3361240[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I154fcd3171f1231e825ee603d53ecfe8[8]        <=  I07b2a00225c337eed1e5a350f3361240[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I07b2a00225c337eed1e5a350f3361240[8] + 1 :
                                             I07b2a00225c337eed1e5a350f3361240[8] ;
            Ib0bf69cc797f330fb2546eb46d2d6f76[8]  <=  I07b2a00225c337eed1e5a350f3361240[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I154fcd3171f1231e825ee603d53ecfe8[9]        <=  I07b2a00225c337eed1e5a350f3361240[9][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I07b2a00225c337eed1e5a350f3361240[9] + 1 :
                                             I07b2a00225c337eed1e5a350f3361240[9] ;
            Ib0bf69cc797f330fb2546eb46d2d6f76[9]  <=  I07b2a00225c337eed1e5a350f3361240[9][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I489e70342dbba4a551097e3064dc9835[0]        <=  I64c650bb94f04521a5a33efa937d9cfc[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I64c650bb94f04521a5a33efa937d9cfc[0] + 1 :
                                             I64c650bb94f04521a5a33efa937d9cfc[0] ;
            Iec7404bc79c58d4d2538fcdf659e9134[0]  <=  I64c650bb94f04521a5a33efa937d9cfc[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I489e70342dbba4a551097e3064dc9835[1]        <=  I64c650bb94f04521a5a33efa937d9cfc[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I64c650bb94f04521a5a33efa937d9cfc[1] + 1 :
                                             I64c650bb94f04521a5a33efa937d9cfc[1] ;
            Iec7404bc79c58d4d2538fcdf659e9134[1]  <=  I64c650bb94f04521a5a33efa937d9cfc[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I489e70342dbba4a551097e3064dc9835[2]        <=  I64c650bb94f04521a5a33efa937d9cfc[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I64c650bb94f04521a5a33efa937d9cfc[2] + 1 :
                                             I64c650bb94f04521a5a33efa937d9cfc[2] ;
            Iec7404bc79c58d4d2538fcdf659e9134[2]  <=  I64c650bb94f04521a5a33efa937d9cfc[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I489e70342dbba4a551097e3064dc9835[3]        <=  I64c650bb94f04521a5a33efa937d9cfc[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I64c650bb94f04521a5a33efa937d9cfc[3] + 1 :
                                             I64c650bb94f04521a5a33efa937d9cfc[3] ;
            Iec7404bc79c58d4d2538fcdf659e9134[3]  <=  I64c650bb94f04521a5a33efa937d9cfc[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I489e70342dbba4a551097e3064dc9835[4]        <=  I64c650bb94f04521a5a33efa937d9cfc[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I64c650bb94f04521a5a33efa937d9cfc[4] + 1 :
                                             I64c650bb94f04521a5a33efa937d9cfc[4] ;
            Iec7404bc79c58d4d2538fcdf659e9134[4]  <=  I64c650bb94f04521a5a33efa937d9cfc[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I489e70342dbba4a551097e3064dc9835[5]        <=  I64c650bb94f04521a5a33efa937d9cfc[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I64c650bb94f04521a5a33efa937d9cfc[5] + 1 :
                                             I64c650bb94f04521a5a33efa937d9cfc[5] ;
            Iec7404bc79c58d4d2538fcdf659e9134[5]  <=  I64c650bb94f04521a5a33efa937d9cfc[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I489e70342dbba4a551097e3064dc9835[6]        <=  I64c650bb94f04521a5a33efa937d9cfc[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I64c650bb94f04521a5a33efa937d9cfc[6] + 1 :
                                             I64c650bb94f04521a5a33efa937d9cfc[6] ;
            Iec7404bc79c58d4d2538fcdf659e9134[6]  <=  I64c650bb94f04521a5a33efa937d9cfc[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I489e70342dbba4a551097e3064dc9835[7]        <=  I64c650bb94f04521a5a33efa937d9cfc[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I64c650bb94f04521a5a33efa937d9cfc[7] + 1 :
                                             I64c650bb94f04521a5a33efa937d9cfc[7] ;
            Iec7404bc79c58d4d2538fcdf659e9134[7]  <=  I64c650bb94f04521a5a33efa937d9cfc[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I489e70342dbba4a551097e3064dc9835[8]        <=  I64c650bb94f04521a5a33efa937d9cfc[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I64c650bb94f04521a5a33efa937d9cfc[8] + 1 :
                                             I64c650bb94f04521a5a33efa937d9cfc[8] ;
            Iec7404bc79c58d4d2538fcdf659e9134[8]  <=  I64c650bb94f04521a5a33efa937d9cfc[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I489e70342dbba4a551097e3064dc9835[9]        <=  I64c650bb94f04521a5a33efa937d9cfc[9][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I64c650bb94f04521a5a33efa937d9cfc[9] + 1 :
                                             I64c650bb94f04521a5a33efa937d9cfc[9] ;
            Iec7404bc79c58d4d2538fcdf659e9134[9]  <=  I64c650bb94f04521a5a33efa937d9cfc[9][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0b0a1f577a212bd9024c8b9a44c92e00[0]        <=  I34152d4ef2dadfcc943a004e81d175f1[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I34152d4ef2dadfcc943a004e81d175f1[0] + 1 :
                                             I34152d4ef2dadfcc943a004e81d175f1[0] ;
            Ie1cd04c7668d3f450c387a6c1ad778c7[0]  <=  I34152d4ef2dadfcc943a004e81d175f1[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0b0a1f577a212bd9024c8b9a44c92e00[1]        <=  I34152d4ef2dadfcc943a004e81d175f1[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I34152d4ef2dadfcc943a004e81d175f1[1] + 1 :
                                             I34152d4ef2dadfcc943a004e81d175f1[1] ;
            Ie1cd04c7668d3f450c387a6c1ad778c7[1]  <=  I34152d4ef2dadfcc943a004e81d175f1[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0b0a1f577a212bd9024c8b9a44c92e00[2]        <=  I34152d4ef2dadfcc943a004e81d175f1[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I34152d4ef2dadfcc943a004e81d175f1[2] + 1 :
                                             I34152d4ef2dadfcc943a004e81d175f1[2] ;
            Ie1cd04c7668d3f450c387a6c1ad778c7[2]  <=  I34152d4ef2dadfcc943a004e81d175f1[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0b0a1f577a212bd9024c8b9a44c92e00[3]        <=  I34152d4ef2dadfcc943a004e81d175f1[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I34152d4ef2dadfcc943a004e81d175f1[3] + 1 :
                                             I34152d4ef2dadfcc943a004e81d175f1[3] ;
            Ie1cd04c7668d3f450c387a6c1ad778c7[3]  <=  I34152d4ef2dadfcc943a004e81d175f1[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0b0a1f577a212bd9024c8b9a44c92e00[4]        <=  I34152d4ef2dadfcc943a004e81d175f1[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I34152d4ef2dadfcc943a004e81d175f1[4] + 1 :
                                             I34152d4ef2dadfcc943a004e81d175f1[4] ;
            Ie1cd04c7668d3f450c387a6c1ad778c7[4]  <=  I34152d4ef2dadfcc943a004e81d175f1[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0b0a1f577a212bd9024c8b9a44c92e00[5]        <=  I34152d4ef2dadfcc943a004e81d175f1[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I34152d4ef2dadfcc943a004e81d175f1[5] + 1 :
                                             I34152d4ef2dadfcc943a004e81d175f1[5] ;
            Ie1cd04c7668d3f450c387a6c1ad778c7[5]  <=  I34152d4ef2dadfcc943a004e81d175f1[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0b0a1f577a212bd9024c8b9a44c92e00[6]        <=  I34152d4ef2dadfcc943a004e81d175f1[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I34152d4ef2dadfcc943a004e81d175f1[6] + 1 :
                                             I34152d4ef2dadfcc943a004e81d175f1[6] ;
            Ie1cd04c7668d3f450c387a6c1ad778c7[6]  <=  I34152d4ef2dadfcc943a004e81d175f1[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0b0a1f577a212bd9024c8b9a44c92e00[7]        <=  I34152d4ef2dadfcc943a004e81d175f1[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I34152d4ef2dadfcc943a004e81d175f1[7] + 1 :
                                             I34152d4ef2dadfcc943a004e81d175f1[7] ;
            Ie1cd04c7668d3f450c387a6c1ad778c7[7]  <=  I34152d4ef2dadfcc943a004e81d175f1[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0b0a1f577a212bd9024c8b9a44c92e00[8]        <=  I34152d4ef2dadfcc943a004e81d175f1[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I34152d4ef2dadfcc943a004e81d175f1[8] + 1 :
                                             I34152d4ef2dadfcc943a004e81d175f1[8] ;
            Ie1cd04c7668d3f450c387a6c1ad778c7[8]  <=  I34152d4ef2dadfcc943a004e81d175f1[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0b0a1f577a212bd9024c8b9a44c92e00[9]        <=  I34152d4ef2dadfcc943a004e81d175f1[9][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I34152d4ef2dadfcc943a004e81d175f1[9] + 1 :
                                             I34152d4ef2dadfcc943a004e81d175f1[9] ;
            Ie1cd04c7668d3f450c387a6c1ad778c7[9]  <=  I34152d4ef2dadfcc943a004e81d175f1[9][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I40d311bab75b73e3788c50115a205270[0]        <=  I745f84653760acc2d83607dcbe1eec73[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I745f84653760acc2d83607dcbe1eec73[0] + 1 :
                                             I745f84653760acc2d83607dcbe1eec73[0] ;
            If511a6ea6aa5cda5353658d8e192791f[0]  <=  I745f84653760acc2d83607dcbe1eec73[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I40d311bab75b73e3788c50115a205270[1]        <=  I745f84653760acc2d83607dcbe1eec73[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I745f84653760acc2d83607dcbe1eec73[1] + 1 :
                                             I745f84653760acc2d83607dcbe1eec73[1] ;
            If511a6ea6aa5cda5353658d8e192791f[1]  <=  I745f84653760acc2d83607dcbe1eec73[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I40d311bab75b73e3788c50115a205270[2]        <=  I745f84653760acc2d83607dcbe1eec73[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I745f84653760acc2d83607dcbe1eec73[2] + 1 :
                                             I745f84653760acc2d83607dcbe1eec73[2] ;
            If511a6ea6aa5cda5353658d8e192791f[2]  <=  I745f84653760acc2d83607dcbe1eec73[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I40d311bab75b73e3788c50115a205270[3]        <=  I745f84653760acc2d83607dcbe1eec73[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I745f84653760acc2d83607dcbe1eec73[3] + 1 :
                                             I745f84653760acc2d83607dcbe1eec73[3] ;
            If511a6ea6aa5cda5353658d8e192791f[3]  <=  I745f84653760acc2d83607dcbe1eec73[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I40d311bab75b73e3788c50115a205270[4]        <=  I745f84653760acc2d83607dcbe1eec73[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I745f84653760acc2d83607dcbe1eec73[4] + 1 :
                                             I745f84653760acc2d83607dcbe1eec73[4] ;
            If511a6ea6aa5cda5353658d8e192791f[4]  <=  I745f84653760acc2d83607dcbe1eec73[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I40d311bab75b73e3788c50115a205270[5]        <=  I745f84653760acc2d83607dcbe1eec73[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I745f84653760acc2d83607dcbe1eec73[5] + 1 :
                                             I745f84653760acc2d83607dcbe1eec73[5] ;
            If511a6ea6aa5cda5353658d8e192791f[5]  <=  I745f84653760acc2d83607dcbe1eec73[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I40d311bab75b73e3788c50115a205270[6]        <=  I745f84653760acc2d83607dcbe1eec73[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I745f84653760acc2d83607dcbe1eec73[6] + 1 :
                                             I745f84653760acc2d83607dcbe1eec73[6] ;
            If511a6ea6aa5cda5353658d8e192791f[6]  <=  I745f84653760acc2d83607dcbe1eec73[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I40d311bab75b73e3788c50115a205270[7]        <=  I745f84653760acc2d83607dcbe1eec73[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I745f84653760acc2d83607dcbe1eec73[7] + 1 :
                                             I745f84653760acc2d83607dcbe1eec73[7] ;
            If511a6ea6aa5cda5353658d8e192791f[7]  <=  I745f84653760acc2d83607dcbe1eec73[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I40d311bab75b73e3788c50115a205270[8]        <=  I745f84653760acc2d83607dcbe1eec73[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I745f84653760acc2d83607dcbe1eec73[8] + 1 :
                                             I745f84653760acc2d83607dcbe1eec73[8] ;
            If511a6ea6aa5cda5353658d8e192791f[8]  <=  I745f84653760acc2d83607dcbe1eec73[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I40d311bab75b73e3788c50115a205270[9]        <=  I745f84653760acc2d83607dcbe1eec73[9][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I745f84653760acc2d83607dcbe1eec73[9] + 1 :
                                             I745f84653760acc2d83607dcbe1eec73[9] ;
            If511a6ea6aa5cda5353658d8e192791f[9]  <=  I745f84653760acc2d83607dcbe1eec73[9][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5fa015a360308bffc46921d119b60c1b[0]        <=  I9efcf5ce8571b24b590d2d4c8161d49d[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I9efcf5ce8571b24b590d2d4c8161d49d[0] + 1 :
                                             I9efcf5ce8571b24b590d2d4c8161d49d[0] ;
            Id88b9265ff08e0730e6a41abe1f80a32[0]  <=  I9efcf5ce8571b24b590d2d4c8161d49d[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5fa015a360308bffc46921d119b60c1b[1]        <=  I9efcf5ce8571b24b590d2d4c8161d49d[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I9efcf5ce8571b24b590d2d4c8161d49d[1] + 1 :
                                             I9efcf5ce8571b24b590d2d4c8161d49d[1] ;
            Id88b9265ff08e0730e6a41abe1f80a32[1]  <=  I9efcf5ce8571b24b590d2d4c8161d49d[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5fa015a360308bffc46921d119b60c1b[2]        <=  I9efcf5ce8571b24b590d2d4c8161d49d[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I9efcf5ce8571b24b590d2d4c8161d49d[2] + 1 :
                                             I9efcf5ce8571b24b590d2d4c8161d49d[2] ;
            Id88b9265ff08e0730e6a41abe1f80a32[2]  <=  I9efcf5ce8571b24b590d2d4c8161d49d[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5fa015a360308bffc46921d119b60c1b[3]        <=  I9efcf5ce8571b24b590d2d4c8161d49d[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I9efcf5ce8571b24b590d2d4c8161d49d[3] + 1 :
                                             I9efcf5ce8571b24b590d2d4c8161d49d[3] ;
            Id88b9265ff08e0730e6a41abe1f80a32[3]  <=  I9efcf5ce8571b24b590d2d4c8161d49d[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5fa015a360308bffc46921d119b60c1b[4]        <=  I9efcf5ce8571b24b590d2d4c8161d49d[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I9efcf5ce8571b24b590d2d4c8161d49d[4] + 1 :
                                             I9efcf5ce8571b24b590d2d4c8161d49d[4] ;
            Id88b9265ff08e0730e6a41abe1f80a32[4]  <=  I9efcf5ce8571b24b590d2d4c8161d49d[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9e42bc767599ce3cc4e2d886e5ef2e62[0]        <=  I60a6ef79e3a8244ad32b9833a6ec196b[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I60a6ef79e3a8244ad32b9833a6ec196b[0] + 1 :
                                             I60a6ef79e3a8244ad32b9833a6ec196b[0] ;
            I6330943c9295298c53e889d47c7904d9[0]  <=  I60a6ef79e3a8244ad32b9833a6ec196b[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9e42bc767599ce3cc4e2d886e5ef2e62[1]        <=  I60a6ef79e3a8244ad32b9833a6ec196b[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I60a6ef79e3a8244ad32b9833a6ec196b[1] + 1 :
                                             I60a6ef79e3a8244ad32b9833a6ec196b[1] ;
            I6330943c9295298c53e889d47c7904d9[1]  <=  I60a6ef79e3a8244ad32b9833a6ec196b[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9e42bc767599ce3cc4e2d886e5ef2e62[2]        <=  I60a6ef79e3a8244ad32b9833a6ec196b[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I60a6ef79e3a8244ad32b9833a6ec196b[2] + 1 :
                                             I60a6ef79e3a8244ad32b9833a6ec196b[2] ;
            I6330943c9295298c53e889d47c7904d9[2]  <=  I60a6ef79e3a8244ad32b9833a6ec196b[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9e42bc767599ce3cc4e2d886e5ef2e62[3]        <=  I60a6ef79e3a8244ad32b9833a6ec196b[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I60a6ef79e3a8244ad32b9833a6ec196b[3] + 1 :
                                             I60a6ef79e3a8244ad32b9833a6ec196b[3] ;
            I6330943c9295298c53e889d47c7904d9[3]  <=  I60a6ef79e3a8244ad32b9833a6ec196b[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9e42bc767599ce3cc4e2d886e5ef2e62[4]        <=  I60a6ef79e3a8244ad32b9833a6ec196b[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I60a6ef79e3a8244ad32b9833a6ec196b[4] + 1 :
                                             I60a6ef79e3a8244ad32b9833a6ec196b[4] ;
            I6330943c9295298c53e889d47c7904d9[4]  <=  I60a6ef79e3a8244ad32b9833a6ec196b[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iea43b150eabf3c7781275821eee3e0c1[0]        <=  I849584bb1c2436f764968afcbb14a61b[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I849584bb1c2436f764968afcbb14a61b[0] + 1 :
                                             I849584bb1c2436f764968afcbb14a61b[0] ;
            I5686b595177e07dd5bf231a35ee41659[0]  <=  I849584bb1c2436f764968afcbb14a61b[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iea43b150eabf3c7781275821eee3e0c1[1]        <=  I849584bb1c2436f764968afcbb14a61b[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I849584bb1c2436f764968afcbb14a61b[1] + 1 :
                                             I849584bb1c2436f764968afcbb14a61b[1] ;
            I5686b595177e07dd5bf231a35ee41659[1]  <=  I849584bb1c2436f764968afcbb14a61b[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iea43b150eabf3c7781275821eee3e0c1[2]        <=  I849584bb1c2436f764968afcbb14a61b[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I849584bb1c2436f764968afcbb14a61b[2] + 1 :
                                             I849584bb1c2436f764968afcbb14a61b[2] ;
            I5686b595177e07dd5bf231a35ee41659[2]  <=  I849584bb1c2436f764968afcbb14a61b[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iea43b150eabf3c7781275821eee3e0c1[3]        <=  I849584bb1c2436f764968afcbb14a61b[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I849584bb1c2436f764968afcbb14a61b[3] + 1 :
                                             I849584bb1c2436f764968afcbb14a61b[3] ;
            I5686b595177e07dd5bf231a35ee41659[3]  <=  I849584bb1c2436f764968afcbb14a61b[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iea43b150eabf3c7781275821eee3e0c1[4]        <=  I849584bb1c2436f764968afcbb14a61b[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I849584bb1c2436f764968afcbb14a61b[4] + 1 :
                                             I849584bb1c2436f764968afcbb14a61b[4] ;
            I5686b595177e07dd5bf231a35ee41659[4]  <=  I849584bb1c2436f764968afcbb14a61b[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8012eea3d53fa4e000eb28b121e02ada[0]        <=  I3ed70f2b460f9278ddeebaf6919b77e8[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I3ed70f2b460f9278ddeebaf6919b77e8[0] + 1 :
                                             I3ed70f2b460f9278ddeebaf6919b77e8[0] ;
            I9c0b88a0be66d62f8ab061aeaee7e60f[0]  <=  I3ed70f2b460f9278ddeebaf6919b77e8[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8012eea3d53fa4e000eb28b121e02ada[1]        <=  I3ed70f2b460f9278ddeebaf6919b77e8[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I3ed70f2b460f9278ddeebaf6919b77e8[1] + 1 :
                                             I3ed70f2b460f9278ddeebaf6919b77e8[1] ;
            I9c0b88a0be66d62f8ab061aeaee7e60f[1]  <=  I3ed70f2b460f9278ddeebaf6919b77e8[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8012eea3d53fa4e000eb28b121e02ada[2]        <=  I3ed70f2b460f9278ddeebaf6919b77e8[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I3ed70f2b460f9278ddeebaf6919b77e8[2] + 1 :
                                             I3ed70f2b460f9278ddeebaf6919b77e8[2] ;
            I9c0b88a0be66d62f8ab061aeaee7e60f[2]  <=  I3ed70f2b460f9278ddeebaf6919b77e8[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8012eea3d53fa4e000eb28b121e02ada[3]        <=  I3ed70f2b460f9278ddeebaf6919b77e8[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I3ed70f2b460f9278ddeebaf6919b77e8[3] + 1 :
                                             I3ed70f2b460f9278ddeebaf6919b77e8[3] ;
            I9c0b88a0be66d62f8ab061aeaee7e60f[3]  <=  I3ed70f2b460f9278ddeebaf6919b77e8[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8012eea3d53fa4e000eb28b121e02ada[4]        <=  I3ed70f2b460f9278ddeebaf6919b77e8[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I3ed70f2b460f9278ddeebaf6919b77e8[4] + 1 :
                                             I3ed70f2b460f9278ddeebaf6919b77e8[4] ;
            I9c0b88a0be66d62f8ab061aeaee7e60f[4]  <=  I3ed70f2b460f9278ddeebaf6919b77e8[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I49804415d20c0c087f802b25dd609887[0]        <=  I37b4978577c93e476e4a0bc15b9008c9[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I37b4978577c93e476e4a0bc15b9008c9[0] + 1 :
                                             I37b4978577c93e476e4a0bc15b9008c9[0] ;
            I9ef21ef20099af28d9a8c794f70d45a5[0]  <=  I37b4978577c93e476e4a0bc15b9008c9[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I49804415d20c0c087f802b25dd609887[1]        <=  I37b4978577c93e476e4a0bc15b9008c9[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I37b4978577c93e476e4a0bc15b9008c9[1] + 1 :
                                             I37b4978577c93e476e4a0bc15b9008c9[1] ;
            I9ef21ef20099af28d9a8c794f70d45a5[1]  <=  I37b4978577c93e476e4a0bc15b9008c9[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I49804415d20c0c087f802b25dd609887[2]        <=  I37b4978577c93e476e4a0bc15b9008c9[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I37b4978577c93e476e4a0bc15b9008c9[2] + 1 :
                                             I37b4978577c93e476e4a0bc15b9008c9[2] ;
            I9ef21ef20099af28d9a8c794f70d45a5[2]  <=  I37b4978577c93e476e4a0bc15b9008c9[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I49804415d20c0c087f802b25dd609887[3]        <=  I37b4978577c93e476e4a0bc15b9008c9[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I37b4978577c93e476e4a0bc15b9008c9[3] + 1 :
                                             I37b4978577c93e476e4a0bc15b9008c9[3] ;
            I9ef21ef20099af28d9a8c794f70d45a5[3]  <=  I37b4978577c93e476e4a0bc15b9008c9[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I49804415d20c0c087f802b25dd609887[4]        <=  I37b4978577c93e476e4a0bc15b9008c9[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I37b4978577c93e476e4a0bc15b9008c9[4] + 1 :
                                             I37b4978577c93e476e4a0bc15b9008c9[4] ;
            I9ef21ef20099af28d9a8c794f70d45a5[4]  <=  I37b4978577c93e476e4a0bc15b9008c9[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id270f05bf5c3fc0bb211d1665d149044[0]        <=  Ieeaf46eef680115f0d2d108b84b5d3da[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ieeaf46eef680115f0d2d108b84b5d3da[0] + 1 :
                                             Ieeaf46eef680115f0d2d108b84b5d3da[0] ;
            Ic2941d16ae6a5cbce70e8546a18ca4ff[0]  <=  Ieeaf46eef680115f0d2d108b84b5d3da[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id270f05bf5c3fc0bb211d1665d149044[1]        <=  Ieeaf46eef680115f0d2d108b84b5d3da[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ieeaf46eef680115f0d2d108b84b5d3da[1] + 1 :
                                             Ieeaf46eef680115f0d2d108b84b5d3da[1] ;
            Ic2941d16ae6a5cbce70e8546a18ca4ff[1]  <=  Ieeaf46eef680115f0d2d108b84b5d3da[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id270f05bf5c3fc0bb211d1665d149044[2]        <=  Ieeaf46eef680115f0d2d108b84b5d3da[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ieeaf46eef680115f0d2d108b84b5d3da[2] + 1 :
                                             Ieeaf46eef680115f0d2d108b84b5d3da[2] ;
            Ic2941d16ae6a5cbce70e8546a18ca4ff[2]  <=  Ieeaf46eef680115f0d2d108b84b5d3da[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id270f05bf5c3fc0bb211d1665d149044[3]        <=  Ieeaf46eef680115f0d2d108b84b5d3da[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ieeaf46eef680115f0d2d108b84b5d3da[3] + 1 :
                                             Ieeaf46eef680115f0d2d108b84b5d3da[3] ;
            Ic2941d16ae6a5cbce70e8546a18ca4ff[3]  <=  Ieeaf46eef680115f0d2d108b84b5d3da[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id270f05bf5c3fc0bb211d1665d149044[4]        <=  Ieeaf46eef680115f0d2d108b84b5d3da[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ieeaf46eef680115f0d2d108b84b5d3da[4] + 1 :
                                             Ieeaf46eef680115f0d2d108b84b5d3da[4] ;
            Ic2941d16ae6a5cbce70e8546a18ca4ff[4]  <=  Ieeaf46eef680115f0d2d108b84b5d3da[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If091fe044c792be711325c103b84cf1d[0]        <=  I8b4ff33c17efa28c7eff64664384cffe[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8b4ff33c17efa28c7eff64664384cffe[0] + 1 :
                                             I8b4ff33c17efa28c7eff64664384cffe[0] ;
            I8e29ebe9ee25ea8ef3e52ff56fc29157[0]  <=  I8b4ff33c17efa28c7eff64664384cffe[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If091fe044c792be711325c103b84cf1d[1]        <=  I8b4ff33c17efa28c7eff64664384cffe[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8b4ff33c17efa28c7eff64664384cffe[1] + 1 :
                                             I8b4ff33c17efa28c7eff64664384cffe[1] ;
            I8e29ebe9ee25ea8ef3e52ff56fc29157[1]  <=  I8b4ff33c17efa28c7eff64664384cffe[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If091fe044c792be711325c103b84cf1d[2]        <=  I8b4ff33c17efa28c7eff64664384cffe[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8b4ff33c17efa28c7eff64664384cffe[2] + 1 :
                                             I8b4ff33c17efa28c7eff64664384cffe[2] ;
            I8e29ebe9ee25ea8ef3e52ff56fc29157[2]  <=  I8b4ff33c17efa28c7eff64664384cffe[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If091fe044c792be711325c103b84cf1d[3]        <=  I8b4ff33c17efa28c7eff64664384cffe[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8b4ff33c17efa28c7eff64664384cffe[3] + 1 :
                                             I8b4ff33c17efa28c7eff64664384cffe[3] ;
            I8e29ebe9ee25ea8ef3e52ff56fc29157[3]  <=  I8b4ff33c17efa28c7eff64664384cffe[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If091fe044c792be711325c103b84cf1d[4]        <=  I8b4ff33c17efa28c7eff64664384cffe[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8b4ff33c17efa28c7eff64664384cffe[4] + 1 :
                                             I8b4ff33c17efa28c7eff64664384cffe[4] ;
            I8e29ebe9ee25ea8ef3e52ff56fc29157[4]  <=  I8b4ff33c17efa28c7eff64664384cffe[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1550db301291ab131a5536147fb938f6[0]        <=  Ia453e66ce9c1335efac95deebe00c249[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia453e66ce9c1335efac95deebe00c249[0] + 1 :
                                             Ia453e66ce9c1335efac95deebe00c249[0] ;
            Ic3742290179b27b9865f9d1f88d66266[0]  <=  Ia453e66ce9c1335efac95deebe00c249[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1550db301291ab131a5536147fb938f6[1]        <=  Ia453e66ce9c1335efac95deebe00c249[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia453e66ce9c1335efac95deebe00c249[1] + 1 :
                                             Ia453e66ce9c1335efac95deebe00c249[1] ;
            Ic3742290179b27b9865f9d1f88d66266[1]  <=  Ia453e66ce9c1335efac95deebe00c249[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1550db301291ab131a5536147fb938f6[2]        <=  Ia453e66ce9c1335efac95deebe00c249[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia453e66ce9c1335efac95deebe00c249[2] + 1 :
                                             Ia453e66ce9c1335efac95deebe00c249[2] ;
            Ic3742290179b27b9865f9d1f88d66266[2]  <=  Ia453e66ce9c1335efac95deebe00c249[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1550db301291ab131a5536147fb938f6[3]        <=  Ia453e66ce9c1335efac95deebe00c249[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia453e66ce9c1335efac95deebe00c249[3] + 1 :
                                             Ia453e66ce9c1335efac95deebe00c249[3] ;
            Ic3742290179b27b9865f9d1f88d66266[3]  <=  Ia453e66ce9c1335efac95deebe00c249[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1550db301291ab131a5536147fb938f6[4]        <=  Ia453e66ce9c1335efac95deebe00c249[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia453e66ce9c1335efac95deebe00c249[4] + 1 :
                                             Ia453e66ce9c1335efac95deebe00c249[4] ;
            Ic3742290179b27b9865f9d1f88d66266[4]  <=  Ia453e66ce9c1335efac95deebe00c249[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I74d1345ee56f5688f875823a5d7c1f4f[0]        <=  I9c5decf5be3d3e4222559a9c244afc6b[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I9c5decf5be3d3e4222559a9c244afc6b[0] + 1 :
                                             I9c5decf5be3d3e4222559a9c244afc6b[0] ;
            I04302edb2671c5bc0ca2673cd53935e1[0]  <=  I9c5decf5be3d3e4222559a9c244afc6b[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I74d1345ee56f5688f875823a5d7c1f4f[1]        <=  I9c5decf5be3d3e4222559a9c244afc6b[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I9c5decf5be3d3e4222559a9c244afc6b[1] + 1 :
                                             I9c5decf5be3d3e4222559a9c244afc6b[1] ;
            I04302edb2671c5bc0ca2673cd53935e1[1]  <=  I9c5decf5be3d3e4222559a9c244afc6b[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I74d1345ee56f5688f875823a5d7c1f4f[2]        <=  I9c5decf5be3d3e4222559a9c244afc6b[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I9c5decf5be3d3e4222559a9c244afc6b[2] + 1 :
                                             I9c5decf5be3d3e4222559a9c244afc6b[2] ;
            I04302edb2671c5bc0ca2673cd53935e1[2]  <=  I9c5decf5be3d3e4222559a9c244afc6b[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I74d1345ee56f5688f875823a5d7c1f4f[3]        <=  I9c5decf5be3d3e4222559a9c244afc6b[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I9c5decf5be3d3e4222559a9c244afc6b[3] + 1 :
                                             I9c5decf5be3d3e4222559a9c244afc6b[3] ;
            I04302edb2671c5bc0ca2673cd53935e1[3]  <=  I9c5decf5be3d3e4222559a9c244afc6b[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I74d1345ee56f5688f875823a5d7c1f4f[4]        <=  I9c5decf5be3d3e4222559a9c244afc6b[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I9c5decf5be3d3e4222559a9c244afc6b[4] + 1 :
                                             I9c5decf5be3d3e4222559a9c244afc6b[4] ;
            I04302edb2671c5bc0ca2673cd53935e1[4]  <=  I9c5decf5be3d3e4222559a9c244afc6b[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I74d1345ee56f5688f875823a5d7c1f4f[5]        <=  I9c5decf5be3d3e4222559a9c244afc6b[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I9c5decf5be3d3e4222559a9c244afc6b[5] + 1 :
                                             I9c5decf5be3d3e4222559a9c244afc6b[5] ;
            I04302edb2671c5bc0ca2673cd53935e1[5]  <=  I9c5decf5be3d3e4222559a9c244afc6b[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I74d1345ee56f5688f875823a5d7c1f4f[6]        <=  I9c5decf5be3d3e4222559a9c244afc6b[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I9c5decf5be3d3e4222559a9c244afc6b[6] + 1 :
                                             I9c5decf5be3d3e4222559a9c244afc6b[6] ;
            I04302edb2671c5bc0ca2673cd53935e1[6]  <=  I9c5decf5be3d3e4222559a9c244afc6b[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I74d1345ee56f5688f875823a5d7c1f4f[7]        <=  I9c5decf5be3d3e4222559a9c244afc6b[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I9c5decf5be3d3e4222559a9c244afc6b[7] + 1 :
                                             I9c5decf5be3d3e4222559a9c244afc6b[7] ;
            I04302edb2671c5bc0ca2673cd53935e1[7]  <=  I9c5decf5be3d3e4222559a9c244afc6b[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I74d1345ee56f5688f875823a5d7c1f4f[8]        <=  I9c5decf5be3d3e4222559a9c244afc6b[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I9c5decf5be3d3e4222559a9c244afc6b[8] + 1 :
                                             I9c5decf5be3d3e4222559a9c244afc6b[8] ;
            I04302edb2671c5bc0ca2673cd53935e1[8]  <=  I9c5decf5be3d3e4222559a9c244afc6b[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I74d1345ee56f5688f875823a5d7c1f4f[9]        <=  I9c5decf5be3d3e4222559a9c244afc6b[9][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I9c5decf5be3d3e4222559a9c244afc6b[9] + 1 :
                                             I9c5decf5be3d3e4222559a9c244afc6b[9] ;
            I04302edb2671c5bc0ca2673cd53935e1[9]  <=  I9c5decf5be3d3e4222559a9c244afc6b[9][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I74d1345ee56f5688f875823a5d7c1f4f[10]        <=  I9c5decf5be3d3e4222559a9c244afc6b[10][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I9c5decf5be3d3e4222559a9c244afc6b[10] + 1 :
                                             I9c5decf5be3d3e4222559a9c244afc6b[10] ;
            I04302edb2671c5bc0ca2673cd53935e1[10]  <=  I9c5decf5be3d3e4222559a9c244afc6b[10][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I74d1345ee56f5688f875823a5d7c1f4f[11]        <=  I9c5decf5be3d3e4222559a9c244afc6b[11][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I9c5decf5be3d3e4222559a9c244afc6b[11] + 1 :
                                             I9c5decf5be3d3e4222559a9c244afc6b[11] ;
            I04302edb2671c5bc0ca2673cd53935e1[11]  <=  I9c5decf5be3d3e4222559a9c244afc6b[11][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I74d1345ee56f5688f875823a5d7c1f4f[12]        <=  I9c5decf5be3d3e4222559a9c244afc6b[12][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I9c5decf5be3d3e4222559a9c244afc6b[12] + 1 :
                                             I9c5decf5be3d3e4222559a9c244afc6b[12] ;
            I04302edb2671c5bc0ca2673cd53935e1[12]  <=  I9c5decf5be3d3e4222559a9c244afc6b[12][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I74d1345ee56f5688f875823a5d7c1f4f[13]        <=  I9c5decf5be3d3e4222559a9c244afc6b[13][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I9c5decf5be3d3e4222559a9c244afc6b[13] + 1 :
                                             I9c5decf5be3d3e4222559a9c244afc6b[13] ;
            I04302edb2671c5bc0ca2673cd53935e1[13]  <=  I9c5decf5be3d3e4222559a9c244afc6b[13][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I187371a49a27a988920854b2bb61bea5[0]        <=  I56c4270727a90e00c295c578183a4dce[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I56c4270727a90e00c295c578183a4dce[0] + 1 :
                                             I56c4270727a90e00c295c578183a4dce[0] ;
            I480a0f6d6c3eb936de10a72749f6cd3f[0]  <=  I56c4270727a90e00c295c578183a4dce[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I187371a49a27a988920854b2bb61bea5[1]        <=  I56c4270727a90e00c295c578183a4dce[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I56c4270727a90e00c295c578183a4dce[1] + 1 :
                                             I56c4270727a90e00c295c578183a4dce[1] ;
            I480a0f6d6c3eb936de10a72749f6cd3f[1]  <=  I56c4270727a90e00c295c578183a4dce[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I187371a49a27a988920854b2bb61bea5[2]        <=  I56c4270727a90e00c295c578183a4dce[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I56c4270727a90e00c295c578183a4dce[2] + 1 :
                                             I56c4270727a90e00c295c578183a4dce[2] ;
            I480a0f6d6c3eb936de10a72749f6cd3f[2]  <=  I56c4270727a90e00c295c578183a4dce[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I187371a49a27a988920854b2bb61bea5[3]        <=  I56c4270727a90e00c295c578183a4dce[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I56c4270727a90e00c295c578183a4dce[3] + 1 :
                                             I56c4270727a90e00c295c578183a4dce[3] ;
            I480a0f6d6c3eb936de10a72749f6cd3f[3]  <=  I56c4270727a90e00c295c578183a4dce[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I187371a49a27a988920854b2bb61bea5[4]        <=  I56c4270727a90e00c295c578183a4dce[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I56c4270727a90e00c295c578183a4dce[4] + 1 :
                                             I56c4270727a90e00c295c578183a4dce[4] ;
            I480a0f6d6c3eb936de10a72749f6cd3f[4]  <=  I56c4270727a90e00c295c578183a4dce[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I187371a49a27a988920854b2bb61bea5[5]        <=  I56c4270727a90e00c295c578183a4dce[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I56c4270727a90e00c295c578183a4dce[5] + 1 :
                                             I56c4270727a90e00c295c578183a4dce[5] ;
            I480a0f6d6c3eb936de10a72749f6cd3f[5]  <=  I56c4270727a90e00c295c578183a4dce[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I187371a49a27a988920854b2bb61bea5[6]        <=  I56c4270727a90e00c295c578183a4dce[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I56c4270727a90e00c295c578183a4dce[6] + 1 :
                                             I56c4270727a90e00c295c578183a4dce[6] ;
            I480a0f6d6c3eb936de10a72749f6cd3f[6]  <=  I56c4270727a90e00c295c578183a4dce[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I187371a49a27a988920854b2bb61bea5[7]        <=  I56c4270727a90e00c295c578183a4dce[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I56c4270727a90e00c295c578183a4dce[7] + 1 :
                                             I56c4270727a90e00c295c578183a4dce[7] ;
            I480a0f6d6c3eb936de10a72749f6cd3f[7]  <=  I56c4270727a90e00c295c578183a4dce[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I187371a49a27a988920854b2bb61bea5[8]        <=  I56c4270727a90e00c295c578183a4dce[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I56c4270727a90e00c295c578183a4dce[8] + 1 :
                                             I56c4270727a90e00c295c578183a4dce[8] ;
            I480a0f6d6c3eb936de10a72749f6cd3f[8]  <=  I56c4270727a90e00c295c578183a4dce[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I187371a49a27a988920854b2bb61bea5[9]        <=  I56c4270727a90e00c295c578183a4dce[9][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I56c4270727a90e00c295c578183a4dce[9] + 1 :
                                             I56c4270727a90e00c295c578183a4dce[9] ;
            I480a0f6d6c3eb936de10a72749f6cd3f[9]  <=  I56c4270727a90e00c295c578183a4dce[9][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I187371a49a27a988920854b2bb61bea5[10]        <=  I56c4270727a90e00c295c578183a4dce[10][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I56c4270727a90e00c295c578183a4dce[10] + 1 :
                                             I56c4270727a90e00c295c578183a4dce[10] ;
            I480a0f6d6c3eb936de10a72749f6cd3f[10]  <=  I56c4270727a90e00c295c578183a4dce[10][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I187371a49a27a988920854b2bb61bea5[11]        <=  I56c4270727a90e00c295c578183a4dce[11][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I56c4270727a90e00c295c578183a4dce[11] + 1 :
                                             I56c4270727a90e00c295c578183a4dce[11] ;
            I480a0f6d6c3eb936de10a72749f6cd3f[11]  <=  I56c4270727a90e00c295c578183a4dce[11][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I187371a49a27a988920854b2bb61bea5[12]        <=  I56c4270727a90e00c295c578183a4dce[12][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I56c4270727a90e00c295c578183a4dce[12] + 1 :
                                             I56c4270727a90e00c295c578183a4dce[12] ;
            I480a0f6d6c3eb936de10a72749f6cd3f[12]  <=  I56c4270727a90e00c295c578183a4dce[12][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I187371a49a27a988920854b2bb61bea5[13]        <=  I56c4270727a90e00c295c578183a4dce[13][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I56c4270727a90e00c295c578183a4dce[13] + 1 :
                                             I56c4270727a90e00c295c578183a4dce[13] ;
            I480a0f6d6c3eb936de10a72749f6cd3f[13]  <=  I56c4270727a90e00c295c578183a4dce[13][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I48c4c6e7414394e3aeff9d17ec25d020[0]        <=  Ib3e1c6976da60eb724a8d00f19368423[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib3e1c6976da60eb724a8d00f19368423[0] + 1 :
                                             Ib3e1c6976da60eb724a8d00f19368423[0] ;
            I50976b0051e84b6a42fc1dbabd7d20ae[0]  <=  Ib3e1c6976da60eb724a8d00f19368423[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I48c4c6e7414394e3aeff9d17ec25d020[1]        <=  Ib3e1c6976da60eb724a8d00f19368423[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib3e1c6976da60eb724a8d00f19368423[1] + 1 :
                                             Ib3e1c6976da60eb724a8d00f19368423[1] ;
            I50976b0051e84b6a42fc1dbabd7d20ae[1]  <=  Ib3e1c6976da60eb724a8d00f19368423[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I48c4c6e7414394e3aeff9d17ec25d020[2]        <=  Ib3e1c6976da60eb724a8d00f19368423[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib3e1c6976da60eb724a8d00f19368423[2] + 1 :
                                             Ib3e1c6976da60eb724a8d00f19368423[2] ;
            I50976b0051e84b6a42fc1dbabd7d20ae[2]  <=  Ib3e1c6976da60eb724a8d00f19368423[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I48c4c6e7414394e3aeff9d17ec25d020[3]        <=  Ib3e1c6976da60eb724a8d00f19368423[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib3e1c6976da60eb724a8d00f19368423[3] + 1 :
                                             Ib3e1c6976da60eb724a8d00f19368423[3] ;
            I50976b0051e84b6a42fc1dbabd7d20ae[3]  <=  Ib3e1c6976da60eb724a8d00f19368423[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I48c4c6e7414394e3aeff9d17ec25d020[4]        <=  Ib3e1c6976da60eb724a8d00f19368423[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib3e1c6976da60eb724a8d00f19368423[4] + 1 :
                                             Ib3e1c6976da60eb724a8d00f19368423[4] ;
            I50976b0051e84b6a42fc1dbabd7d20ae[4]  <=  Ib3e1c6976da60eb724a8d00f19368423[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I48c4c6e7414394e3aeff9d17ec25d020[5]        <=  Ib3e1c6976da60eb724a8d00f19368423[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib3e1c6976da60eb724a8d00f19368423[5] + 1 :
                                             Ib3e1c6976da60eb724a8d00f19368423[5] ;
            I50976b0051e84b6a42fc1dbabd7d20ae[5]  <=  Ib3e1c6976da60eb724a8d00f19368423[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I48c4c6e7414394e3aeff9d17ec25d020[6]        <=  Ib3e1c6976da60eb724a8d00f19368423[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib3e1c6976da60eb724a8d00f19368423[6] + 1 :
                                             Ib3e1c6976da60eb724a8d00f19368423[6] ;
            I50976b0051e84b6a42fc1dbabd7d20ae[6]  <=  Ib3e1c6976da60eb724a8d00f19368423[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I48c4c6e7414394e3aeff9d17ec25d020[7]        <=  Ib3e1c6976da60eb724a8d00f19368423[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib3e1c6976da60eb724a8d00f19368423[7] + 1 :
                                             Ib3e1c6976da60eb724a8d00f19368423[7] ;
            I50976b0051e84b6a42fc1dbabd7d20ae[7]  <=  Ib3e1c6976da60eb724a8d00f19368423[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I48c4c6e7414394e3aeff9d17ec25d020[8]        <=  Ib3e1c6976da60eb724a8d00f19368423[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib3e1c6976da60eb724a8d00f19368423[8] + 1 :
                                             Ib3e1c6976da60eb724a8d00f19368423[8] ;
            I50976b0051e84b6a42fc1dbabd7d20ae[8]  <=  Ib3e1c6976da60eb724a8d00f19368423[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I48c4c6e7414394e3aeff9d17ec25d020[9]        <=  Ib3e1c6976da60eb724a8d00f19368423[9][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib3e1c6976da60eb724a8d00f19368423[9] + 1 :
                                             Ib3e1c6976da60eb724a8d00f19368423[9] ;
            I50976b0051e84b6a42fc1dbabd7d20ae[9]  <=  Ib3e1c6976da60eb724a8d00f19368423[9][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I48c4c6e7414394e3aeff9d17ec25d020[10]        <=  Ib3e1c6976da60eb724a8d00f19368423[10][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib3e1c6976da60eb724a8d00f19368423[10] + 1 :
                                             Ib3e1c6976da60eb724a8d00f19368423[10] ;
            I50976b0051e84b6a42fc1dbabd7d20ae[10]  <=  Ib3e1c6976da60eb724a8d00f19368423[10][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I48c4c6e7414394e3aeff9d17ec25d020[11]        <=  Ib3e1c6976da60eb724a8d00f19368423[11][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib3e1c6976da60eb724a8d00f19368423[11] + 1 :
                                             Ib3e1c6976da60eb724a8d00f19368423[11] ;
            I50976b0051e84b6a42fc1dbabd7d20ae[11]  <=  Ib3e1c6976da60eb724a8d00f19368423[11][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I48c4c6e7414394e3aeff9d17ec25d020[12]        <=  Ib3e1c6976da60eb724a8d00f19368423[12][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib3e1c6976da60eb724a8d00f19368423[12] + 1 :
                                             Ib3e1c6976da60eb724a8d00f19368423[12] ;
            I50976b0051e84b6a42fc1dbabd7d20ae[12]  <=  Ib3e1c6976da60eb724a8d00f19368423[12][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I48c4c6e7414394e3aeff9d17ec25d020[13]        <=  Ib3e1c6976da60eb724a8d00f19368423[13][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib3e1c6976da60eb724a8d00f19368423[13] + 1 :
                                             Ib3e1c6976da60eb724a8d00f19368423[13] ;
            I50976b0051e84b6a42fc1dbabd7d20ae[13]  <=  Ib3e1c6976da60eb724a8d00f19368423[13][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3cba0f4c2ca8c7c200df8e1071ab429d[0]        <=  Ib53ea6bc0e3ac45d5a8eecd5dce775d8[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib53ea6bc0e3ac45d5a8eecd5dce775d8[0] + 1 :
                                             Ib53ea6bc0e3ac45d5a8eecd5dce775d8[0] ;
            I82e0e091fba6f79cef97eacac4b43ecb[0]  <=  Ib53ea6bc0e3ac45d5a8eecd5dce775d8[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3cba0f4c2ca8c7c200df8e1071ab429d[1]        <=  Ib53ea6bc0e3ac45d5a8eecd5dce775d8[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib53ea6bc0e3ac45d5a8eecd5dce775d8[1] + 1 :
                                             Ib53ea6bc0e3ac45d5a8eecd5dce775d8[1] ;
            I82e0e091fba6f79cef97eacac4b43ecb[1]  <=  Ib53ea6bc0e3ac45d5a8eecd5dce775d8[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3cba0f4c2ca8c7c200df8e1071ab429d[2]        <=  Ib53ea6bc0e3ac45d5a8eecd5dce775d8[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib53ea6bc0e3ac45d5a8eecd5dce775d8[2] + 1 :
                                             Ib53ea6bc0e3ac45d5a8eecd5dce775d8[2] ;
            I82e0e091fba6f79cef97eacac4b43ecb[2]  <=  Ib53ea6bc0e3ac45d5a8eecd5dce775d8[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3cba0f4c2ca8c7c200df8e1071ab429d[3]        <=  Ib53ea6bc0e3ac45d5a8eecd5dce775d8[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib53ea6bc0e3ac45d5a8eecd5dce775d8[3] + 1 :
                                             Ib53ea6bc0e3ac45d5a8eecd5dce775d8[3] ;
            I82e0e091fba6f79cef97eacac4b43ecb[3]  <=  Ib53ea6bc0e3ac45d5a8eecd5dce775d8[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3cba0f4c2ca8c7c200df8e1071ab429d[4]        <=  Ib53ea6bc0e3ac45d5a8eecd5dce775d8[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib53ea6bc0e3ac45d5a8eecd5dce775d8[4] + 1 :
                                             Ib53ea6bc0e3ac45d5a8eecd5dce775d8[4] ;
            I82e0e091fba6f79cef97eacac4b43ecb[4]  <=  Ib53ea6bc0e3ac45d5a8eecd5dce775d8[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3cba0f4c2ca8c7c200df8e1071ab429d[5]        <=  Ib53ea6bc0e3ac45d5a8eecd5dce775d8[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib53ea6bc0e3ac45d5a8eecd5dce775d8[5] + 1 :
                                             Ib53ea6bc0e3ac45d5a8eecd5dce775d8[5] ;
            I82e0e091fba6f79cef97eacac4b43ecb[5]  <=  Ib53ea6bc0e3ac45d5a8eecd5dce775d8[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3cba0f4c2ca8c7c200df8e1071ab429d[6]        <=  Ib53ea6bc0e3ac45d5a8eecd5dce775d8[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib53ea6bc0e3ac45d5a8eecd5dce775d8[6] + 1 :
                                             Ib53ea6bc0e3ac45d5a8eecd5dce775d8[6] ;
            I82e0e091fba6f79cef97eacac4b43ecb[6]  <=  Ib53ea6bc0e3ac45d5a8eecd5dce775d8[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3cba0f4c2ca8c7c200df8e1071ab429d[7]        <=  Ib53ea6bc0e3ac45d5a8eecd5dce775d8[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib53ea6bc0e3ac45d5a8eecd5dce775d8[7] + 1 :
                                             Ib53ea6bc0e3ac45d5a8eecd5dce775d8[7] ;
            I82e0e091fba6f79cef97eacac4b43ecb[7]  <=  Ib53ea6bc0e3ac45d5a8eecd5dce775d8[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3cba0f4c2ca8c7c200df8e1071ab429d[8]        <=  Ib53ea6bc0e3ac45d5a8eecd5dce775d8[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib53ea6bc0e3ac45d5a8eecd5dce775d8[8] + 1 :
                                             Ib53ea6bc0e3ac45d5a8eecd5dce775d8[8] ;
            I82e0e091fba6f79cef97eacac4b43ecb[8]  <=  Ib53ea6bc0e3ac45d5a8eecd5dce775d8[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3cba0f4c2ca8c7c200df8e1071ab429d[9]        <=  Ib53ea6bc0e3ac45d5a8eecd5dce775d8[9][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib53ea6bc0e3ac45d5a8eecd5dce775d8[9] + 1 :
                                             Ib53ea6bc0e3ac45d5a8eecd5dce775d8[9] ;
            I82e0e091fba6f79cef97eacac4b43ecb[9]  <=  Ib53ea6bc0e3ac45d5a8eecd5dce775d8[9][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3cba0f4c2ca8c7c200df8e1071ab429d[10]        <=  Ib53ea6bc0e3ac45d5a8eecd5dce775d8[10][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib53ea6bc0e3ac45d5a8eecd5dce775d8[10] + 1 :
                                             Ib53ea6bc0e3ac45d5a8eecd5dce775d8[10] ;
            I82e0e091fba6f79cef97eacac4b43ecb[10]  <=  Ib53ea6bc0e3ac45d5a8eecd5dce775d8[10][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3cba0f4c2ca8c7c200df8e1071ab429d[11]        <=  Ib53ea6bc0e3ac45d5a8eecd5dce775d8[11][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib53ea6bc0e3ac45d5a8eecd5dce775d8[11] + 1 :
                                             Ib53ea6bc0e3ac45d5a8eecd5dce775d8[11] ;
            I82e0e091fba6f79cef97eacac4b43ecb[11]  <=  Ib53ea6bc0e3ac45d5a8eecd5dce775d8[11][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3cba0f4c2ca8c7c200df8e1071ab429d[12]        <=  Ib53ea6bc0e3ac45d5a8eecd5dce775d8[12][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib53ea6bc0e3ac45d5a8eecd5dce775d8[12] + 1 :
                                             Ib53ea6bc0e3ac45d5a8eecd5dce775d8[12] ;
            I82e0e091fba6f79cef97eacac4b43ecb[12]  <=  Ib53ea6bc0e3ac45d5a8eecd5dce775d8[12][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3cba0f4c2ca8c7c200df8e1071ab429d[13]        <=  Ib53ea6bc0e3ac45d5a8eecd5dce775d8[13][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib53ea6bc0e3ac45d5a8eecd5dce775d8[13] + 1 :
                                             Ib53ea6bc0e3ac45d5a8eecd5dce775d8[13] ;
            I82e0e091fba6f79cef97eacac4b43ecb[13]  <=  Ib53ea6bc0e3ac45d5a8eecd5dce775d8[13][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I35688678e1a83ec39d737d9cdfd44ba3[0]        <=  I922408509703b8175883356d89806972[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I922408509703b8175883356d89806972[0] + 1 :
                                             I922408509703b8175883356d89806972[0] ;
            I3d50cfeaa4b69c09bb648b8873a6bc24[0]  <=  I922408509703b8175883356d89806972[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I35688678e1a83ec39d737d9cdfd44ba3[1]        <=  I922408509703b8175883356d89806972[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I922408509703b8175883356d89806972[1] + 1 :
                                             I922408509703b8175883356d89806972[1] ;
            I3d50cfeaa4b69c09bb648b8873a6bc24[1]  <=  I922408509703b8175883356d89806972[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I35688678e1a83ec39d737d9cdfd44ba3[2]        <=  I922408509703b8175883356d89806972[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I922408509703b8175883356d89806972[2] + 1 :
                                             I922408509703b8175883356d89806972[2] ;
            I3d50cfeaa4b69c09bb648b8873a6bc24[2]  <=  I922408509703b8175883356d89806972[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I35688678e1a83ec39d737d9cdfd44ba3[3]        <=  I922408509703b8175883356d89806972[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I922408509703b8175883356d89806972[3] + 1 :
                                             I922408509703b8175883356d89806972[3] ;
            I3d50cfeaa4b69c09bb648b8873a6bc24[3]  <=  I922408509703b8175883356d89806972[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I35688678e1a83ec39d737d9cdfd44ba3[4]        <=  I922408509703b8175883356d89806972[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I922408509703b8175883356d89806972[4] + 1 :
                                             I922408509703b8175883356d89806972[4] ;
            I3d50cfeaa4b69c09bb648b8873a6bc24[4]  <=  I922408509703b8175883356d89806972[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I35688678e1a83ec39d737d9cdfd44ba3[5]        <=  I922408509703b8175883356d89806972[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I922408509703b8175883356d89806972[5] + 1 :
                                             I922408509703b8175883356d89806972[5] ;
            I3d50cfeaa4b69c09bb648b8873a6bc24[5]  <=  I922408509703b8175883356d89806972[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I35688678e1a83ec39d737d9cdfd44ba3[6]        <=  I922408509703b8175883356d89806972[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I922408509703b8175883356d89806972[6] + 1 :
                                             I922408509703b8175883356d89806972[6] ;
            I3d50cfeaa4b69c09bb648b8873a6bc24[6]  <=  I922408509703b8175883356d89806972[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I94b86d31e8226723950096e91855b6d3[0]        <=  I6cabc68155bc4aef952a07f101ea2802[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I6cabc68155bc4aef952a07f101ea2802[0] + 1 :
                                             I6cabc68155bc4aef952a07f101ea2802[0] ;
            I33a6ffad80ddf99a4d316a049078244d[0]  <=  I6cabc68155bc4aef952a07f101ea2802[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I94b86d31e8226723950096e91855b6d3[1]        <=  I6cabc68155bc4aef952a07f101ea2802[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I6cabc68155bc4aef952a07f101ea2802[1] + 1 :
                                             I6cabc68155bc4aef952a07f101ea2802[1] ;
            I33a6ffad80ddf99a4d316a049078244d[1]  <=  I6cabc68155bc4aef952a07f101ea2802[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I94b86d31e8226723950096e91855b6d3[2]        <=  I6cabc68155bc4aef952a07f101ea2802[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I6cabc68155bc4aef952a07f101ea2802[2] + 1 :
                                             I6cabc68155bc4aef952a07f101ea2802[2] ;
            I33a6ffad80ddf99a4d316a049078244d[2]  <=  I6cabc68155bc4aef952a07f101ea2802[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I94b86d31e8226723950096e91855b6d3[3]        <=  I6cabc68155bc4aef952a07f101ea2802[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I6cabc68155bc4aef952a07f101ea2802[3] + 1 :
                                             I6cabc68155bc4aef952a07f101ea2802[3] ;
            I33a6ffad80ddf99a4d316a049078244d[3]  <=  I6cabc68155bc4aef952a07f101ea2802[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I94b86d31e8226723950096e91855b6d3[4]        <=  I6cabc68155bc4aef952a07f101ea2802[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I6cabc68155bc4aef952a07f101ea2802[4] + 1 :
                                             I6cabc68155bc4aef952a07f101ea2802[4] ;
            I33a6ffad80ddf99a4d316a049078244d[4]  <=  I6cabc68155bc4aef952a07f101ea2802[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I94b86d31e8226723950096e91855b6d3[5]        <=  I6cabc68155bc4aef952a07f101ea2802[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I6cabc68155bc4aef952a07f101ea2802[5] + 1 :
                                             I6cabc68155bc4aef952a07f101ea2802[5] ;
            I33a6ffad80ddf99a4d316a049078244d[5]  <=  I6cabc68155bc4aef952a07f101ea2802[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I94b86d31e8226723950096e91855b6d3[6]        <=  I6cabc68155bc4aef952a07f101ea2802[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I6cabc68155bc4aef952a07f101ea2802[6] + 1 :
                                             I6cabc68155bc4aef952a07f101ea2802[6] ;
            I33a6ffad80ddf99a4d316a049078244d[6]  <=  I6cabc68155bc4aef952a07f101ea2802[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0ea7c4721ee0c13ad15a9b0fa7b15ad3[0]        <=  Ia894c8a3585def468e93aa51039d405c[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia894c8a3585def468e93aa51039d405c[0] + 1 :
                                             Ia894c8a3585def468e93aa51039d405c[0] ;
            I980165c1147ac5ff86619c841c6031dc[0]  <=  Ia894c8a3585def468e93aa51039d405c[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0ea7c4721ee0c13ad15a9b0fa7b15ad3[1]        <=  Ia894c8a3585def468e93aa51039d405c[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia894c8a3585def468e93aa51039d405c[1] + 1 :
                                             Ia894c8a3585def468e93aa51039d405c[1] ;
            I980165c1147ac5ff86619c841c6031dc[1]  <=  Ia894c8a3585def468e93aa51039d405c[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0ea7c4721ee0c13ad15a9b0fa7b15ad3[2]        <=  Ia894c8a3585def468e93aa51039d405c[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia894c8a3585def468e93aa51039d405c[2] + 1 :
                                             Ia894c8a3585def468e93aa51039d405c[2] ;
            I980165c1147ac5ff86619c841c6031dc[2]  <=  Ia894c8a3585def468e93aa51039d405c[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0ea7c4721ee0c13ad15a9b0fa7b15ad3[3]        <=  Ia894c8a3585def468e93aa51039d405c[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia894c8a3585def468e93aa51039d405c[3] + 1 :
                                             Ia894c8a3585def468e93aa51039d405c[3] ;
            I980165c1147ac5ff86619c841c6031dc[3]  <=  Ia894c8a3585def468e93aa51039d405c[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0ea7c4721ee0c13ad15a9b0fa7b15ad3[4]        <=  Ia894c8a3585def468e93aa51039d405c[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia894c8a3585def468e93aa51039d405c[4] + 1 :
                                             Ia894c8a3585def468e93aa51039d405c[4] ;
            I980165c1147ac5ff86619c841c6031dc[4]  <=  Ia894c8a3585def468e93aa51039d405c[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0ea7c4721ee0c13ad15a9b0fa7b15ad3[5]        <=  Ia894c8a3585def468e93aa51039d405c[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia894c8a3585def468e93aa51039d405c[5] + 1 :
                                             Ia894c8a3585def468e93aa51039d405c[5] ;
            I980165c1147ac5ff86619c841c6031dc[5]  <=  Ia894c8a3585def468e93aa51039d405c[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0ea7c4721ee0c13ad15a9b0fa7b15ad3[6]        <=  Ia894c8a3585def468e93aa51039d405c[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia894c8a3585def468e93aa51039d405c[6] + 1 :
                                             Ia894c8a3585def468e93aa51039d405c[6] ;
            I980165c1147ac5ff86619c841c6031dc[6]  <=  Ia894c8a3585def468e93aa51039d405c[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I29dd5fb1c2673cd4daa9cafaf24d8e7c[0]        <=  Iaf1c895fc85487f017d3c084e125551c[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Iaf1c895fc85487f017d3c084e125551c[0] + 1 :
                                             Iaf1c895fc85487f017d3c084e125551c[0] ;
            I19df055705f322292a3601fa63f0e5f9[0]  <=  Iaf1c895fc85487f017d3c084e125551c[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I29dd5fb1c2673cd4daa9cafaf24d8e7c[1]        <=  Iaf1c895fc85487f017d3c084e125551c[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Iaf1c895fc85487f017d3c084e125551c[1] + 1 :
                                             Iaf1c895fc85487f017d3c084e125551c[1] ;
            I19df055705f322292a3601fa63f0e5f9[1]  <=  Iaf1c895fc85487f017d3c084e125551c[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I29dd5fb1c2673cd4daa9cafaf24d8e7c[2]        <=  Iaf1c895fc85487f017d3c084e125551c[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Iaf1c895fc85487f017d3c084e125551c[2] + 1 :
                                             Iaf1c895fc85487f017d3c084e125551c[2] ;
            I19df055705f322292a3601fa63f0e5f9[2]  <=  Iaf1c895fc85487f017d3c084e125551c[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I29dd5fb1c2673cd4daa9cafaf24d8e7c[3]        <=  Iaf1c895fc85487f017d3c084e125551c[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Iaf1c895fc85487f017d3c084e125551c[3] + 1 :
                                             Iaf1c895fc85487f017d3c084e125551c[3] ;
            I19df055705f322292a3601fa63f0e5f9[3]  <=  Iaf1c895fc85487f017d3c084e125551c[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I29dd5fb1c2673cd4daa9cafaf24d8e7c[4]        <=  Iaf1c895fc85487f017d3c084e125551c[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Iaf1c895fc85487f017d3c084e125551c[4] + 1 :
                                             Iaf1c895fc85487f017d3c084e125551c[4] ;
            I19df055705f322292a3601fa63f0e5f9[4]  <=  Iaf1c895fc85487f017d3c084e125551c[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I29dd5fb1c2673cd4daa9cafaf24d8e7c[5]        <=  Iaf1c895fc85487f017d3c084e125551c[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Iaf1c895fc85487f017d3c084e125551c[5] + 1 :
                                             Iaf1c895fc85487f017d3c084e125551c[5] ;
            I19df055705f322292a3601fa63f0e5f9[5]  <=  Iaf1c895fc85487f017d3c084e125551c[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I29dd5fb1c2673cd4daa9cafaf24d8e7c[6]        <=  Iaf1c895fc85487f017d3c084e125551c[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Iaf1c895fc85487f017d3c084e125551c[6] + 1 :
                                             Iaf1c895fc85487f017d3c084e125551c[6] ;
            I19df055705f322292a3601fa63f0e5f9[6]  <=  Iaf1c895fc85487f017d3c084e125551c[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iead4c81d836e3befae55049797c30d6b[0]        <=  I63d67a9bf5a46800216b38df1eb185eb[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I63d67a9bf5a46800216b38df1eb185eb[0] + 1 :
                                             I63d67a9bf5a46800216b38df1eb185eb[0] ;
            I0e0b15868b02ca52b260f17f150d237e[0]  <=  I63d67a9bf5a46800216b38df1eb185eb[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iead4c81d836e3befae55049797c30d6b[1]        <=  I63d67a9bf5a46800216b38df1eb185eb[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I63d67a9bf5a46800216b38df1eb185eb[1] + 1 :
                                             I63d67a9bf5a46800216b38df1eb185eb[1] ;
            I0e0b15868b02ca52b260f17f150d237e[1]  <=  I63d67a9bf5a46800216b38df1eb185eb[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iead4c81d836e3befae55049797c30d6b[2]        <=  I63d67a9bf5a46800216b38df1eb185eb[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I63d67a9bf5a46800216b38df1eb185eb[2] + 1 :
                                             I63d67a9bf5a46800216b38df1eb185eb[2] ;
            I0e0b15868b02ca52b260f17f150d237e[2]  <=  I63d67a9bf5a46800216b38df1eb185eb[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iead4c81d836e3befae55049797c30d6b[3]        <=  I63d67a9bf5a46800216b38df1eb185eb[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I63d67a9bf5a46800216b38df1eb185eb[3] + 1 :
                                             I63d67a9bf5a46800216b38df1eb185eb[3] ;
            I0e0b15868b02ca52b260f17f150d237e[3]  <=  I63d67a9bf5a46800216b38df1eb185eb[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iead4c81d836e3befae55049797c30d6b[4]        <=  I63d67a9bf5a46800216b38df1eb185eb[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I63d67a9bf5a46800216b38df1eb185eb[4] + 1 :
                                             I63d67a9bf5a46800216b38df1eb185eb[4] ;
            I0e0b15868b02ca52b260f17f150d237e[4]  <=  I63d67a9bf5a46800216b38df1eb185eb[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iead4c81d836e3befae55049797c30d6b[5]        <=  I63d67a9bf5a46800216b38df1eb185eb[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I63d67a9bf5a46800216b38df1eb185eb[5] + 1 :
                                             I63d67a9bf5a46800216b38df1eb185eb[5] ;
            I0e0b15868b02ca52b260f17f150d237e[5]  <=  I63d67a9bf5a46800216b38df1eb185eb[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iead4c81d836e3befae55049797c30d6b[6]        <=  I63d67a9bf5a46800216b38df1eb185eb[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I63d67a9bf5a46800216b38df1eb185eb[6] + 1 :
                                             I63d67a9bf5a46800216b38df1eb185eb[6] ;
            I0e0b15868b02ca52b260f17f150d237e[6]  <=  I63d67a9bf5a46800216b38df1eb185eb[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iead4c81d836e3befae55049797c30d6b[7]        <=  I63d67a9bf5a46800216b38df1eb185eb[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I63d67a9bf5a46800216b38df1eb185eb[7] + 1 :
                                             I63d67a9bf5a46800216b38df1eb185eb[7] ;
            I0e0b15868b02ca52b260f17f150d237e[7]  <=  I63d67a9bf5a46800216b38df1eb185eb[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iead4c81d836e3befae55049797c30d6b[8]        <=  I63d67a9bf5a46800216b38df1eb185eb[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I63d67a9bf5a46800216b38df1eb185eb[8] + 1 :
                                             I63d67a9bf5a46800216b38df1eb185eb[8] ;
            I0e0b15868b02ca52b260f17f150d237e[8]  <=  I63d67a9bf5a46800216b38df1eb185eb[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iead4c81d836e3befae55049797c30d6b[9]        <=  I63d67a9bf5a46800216b38df1eb185eb[9][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I63d67a9bf5a46800216b38df1eb185eb[9] + 1 :
                                             I63d67a9bf5a46800216b38df1eb185eb[9] ;
            I0e0b15868b02ca52b260f17f150d237e[9]  <=  I63d67a9bf5a46800216b38df1eb185eb[9][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iead4c81d836e3befae55049797c30d6b[10]        <=  I63d67a9bf5a46800216b38df1eb185eb[10][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I63d67a9bf5a46800216b38df1eb185eb[10] + 1 :
                                             I63d67a9bf5a46800216b38df1eb185eb[10] ;
            I0e0b15868b02ca52b260f17f150d237e[10]  <=  I63d67a9bf5a46800216b38df1eb185eb[10][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iead4c81d836e3befae55049797c30d6b[11]        <=  I63d67a9bf5a46800216b38df1eb185eb[11][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I63d67a9bf5a46800216b38df1eb185eb[11] + 1 :
                                             I63d67a9bf5a46800216b38df1eb185eb[11] ;
            I0e0b15868b02ca52b260f17f150d237e[11]  <=  I63d67a9bf5a46800216b38df1eb185eb[11][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iead4c81d836e3befae55049797c30d6b[12]        <=  I63d67a9bf5a46800216b38df1eb185eb[12][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I63d67a9bf5a46800216b38df1eb185eb[12] + 1 :
                                             I63d67a9bf5a46800216b38df1eb185eb[12] ;
            I0e0b15868b02ca52b260f17f150d237e[12]  <=  I63d67a9bf5a46800216b38df1eb185eb[12][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I23e22f44791c167acaba27c91ef3b497[0]        <=  Ic087eef7b3d2a51f34f317a6b9e49144[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic087eef7b3d2a51f34f317a6b9e49144[0] + 1 :
                                             Ic087eef7b3d2a51f34f317a6b9e49144[0] ;
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[0]  <=  Ic087eef7b3d2a51f34f317a6b9e49144[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I23e22f44791c167acaba27c91ef3b497[1]        <=  Ic087eef7b3d2a51f34f317a6b9e49144[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic087eef7b3d2a51f34f317a6b9e49144[1] + 1 :
                                             Ic087eef7b3d2a51f34f317a6b9e49144[1] ;
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[1]  <=  Ic087eef7b3d2a51f34f317a6b9e49144[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I23e22f44791c167acaba27c91ef3b497[2]        <=  Ic087eef7b3d2a51f34f317a6b9e49144[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic087eef7b3d2a51f34f317a6b9e49144[2] + 1 :
                                             Ic087eef7b3d2a51f34f317a6b9e49144[2] ;
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[2]  <=  Ic087eef7b3d2a51f34f317a6b9e49144[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I23e22f44791c167acaba27c91ef3b497[3]        <=  Ic087eef7b3d2a51f34f317a6b9e49144[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic087eef7b3d2a51f34f317a6b9e49144[3] + 1 :
                                             Ic087eef7b3d2a51f34f317a6b9e49144[3] ;
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[3]  <=  Ic087eef7b3d2a51f34f317a6b9e49144[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I23e22f44791c167acaba27c91ef3b497[4]        <=  Ic087eef7b3d2a51f34f317a6b9e49144[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic087eef7b3d2a51f34f317a6b9e49144[4] + 1 :
                                             Ic087eef7b3d2a51f34f317a6b9e49144[4] ;
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[4]  <=  Ic087eef7b3d2a51f34f317a6b9e49144[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I23e22f44791c167acaba27c91ef3b497[5]        <=  Ic087eef7b3d2a51f34f317a6b9e49144[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic087eef7b3d2a51f34f317a6b9e49144[5] + 1 :
                                             Ic087eef7b3d2a51f34f317a6b9e49144[5] ;
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[5]  <=  Ic087eef7b3d2a51f34f317a6b9e49144[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I23e22f44791c167acaba27c91ef3b497[6]        <=  Ic087eef7b3d2a51f34f317a6b9e49144[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic087eef7b3d2a51f34f317a6b9e49144[6] + 1 :
                                             Ic087eef7b3d2a51f34f317a6b9e49144[6] ;
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[6]  <=  Ic087eef7b3d2a51f34f317a6b9e49144[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I23e22f44791c167acaba27c91ef3b497[7]        <=  Ic087eef7b3d2a51f34f317a6b9e49144[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic087eef7b3d2a51f34f317a6b9e49144[7] + 1 :
                                             Ic087eef7b3d2a51f34f317a6b9e49144[7] ;
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[7]  <=  Ic087eef7b3d2a51f34f317a6b9e49144[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I23e22f44791c167acaba27c91ef3b497[8]        <=  Ic087eef7b3d2a51f34f317a6b9e49144[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic087eef7b3d2a51f34f317a6b9e49144[8] + 1 :
                                             Ic087eef7b3d2a51f34f317a6b9e49144[8] ;
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[8]  <=  Ic087eef7b3d2a51f34f317a6b9e49144[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I23e22f44791c167acaba27c91ef3b497[9]        <=  Ic087eef7b3d2a51f34f317a6b9e49144[9][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic087eef7b3d2a51f34f317a6b9e49144[9] + 1 :
                                             Ic087eef7b3d2a51f34f317a6b9e49144[9] ;
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[9]  <=  Ic087eef7b3d2a51f34f317a6b9e49144[9][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I23e22f44791c167acaba27c91ef3b497[10]        <=  Ic087eef7b3d2a51f34f317a6b9e49144[10][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic087eef7b3d2a51f34f317a6b9e49144[10] + 1 :
                                             Ic087eef7b3d2a51f34f317a6b9e49144[10] ;
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[10]  <=  Ic087eef7b3d2a51f34f317a6b9e49144[10][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I23e22f44791c167acaba27c91ef3b497[11]        <=  Ic087eef7b3d2a51f34f317a6b9e49144[11][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic087eef7b3d2a51f34f317a6b9e49144[11] + 1 :
                                             Ic087eef7b3d2a51f34f317a6b9e49144[11] ;
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[11]  <=  Ic087eef7b3d2a51f34f317a6b9e49144[11][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I23e22f44791c167acaba27c91ef3b497[12]        <=  Ic087eef7b3d2a51f34f317a6b9e49144[12][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic087eef7b3d2a51f34f317a6b9e49144[12] + 1 :
                                             Ic087eef7b3d2a51f34f317a6b9e49144[12] ;
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[12]  <=  Ic087eef7b3d2a51f34f317a6b9e49144[12][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic91f087829e0b9e0c964229a2dc567bc[0]        <=  I6d360540762be9eab571c0bfe0500f67[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I6d360540762be9eab571c0bfe0500f67[0] + 1 :
                                             I6d360540762be9eab571c0bfe0500f67[0] ;
            I8e591d83170c8ba46d31c61935311b22[0]  <=  I6d360540762be9eab571c0bfe0500f67[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic91f087829e0b9e0c964229a2dc567bc[1]        <=  I6d360540762be9eab571c0bfe0500f67[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I6d360540762be9eab571c0bfe0500f67[1] + 1 :
                                             I6d360540762be9eab571c0bfe0500f67[1] ;
            I8e591d83170c8ba46d31c61935311b22[1]  <=  I6d360540762be9eab571c0bfe0500f67[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic91f087829e0b9e0c964229a2dc567bc[2]        <=  I6d360540762be9eab571c0bfe0500f67[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I6d360540762be9eab571c0bfe0500f67[2] + 1 :
                                             I6d360540762be9eab571c0bfe0500f67[2] ;
            I8e591d83170c8ba46d31c61935311b22[2]  <=  I6d360540762be9eab571c0bfe0500f67[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic91f087829e0b9e0c964229a2dc567bc[3]        <=  I6d360540762be9eab571c0bfe0500f67[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I6d360540762be9eab571c0bfe0500f67[3] + 1 :
                                             I6d360540762be9eab571c0bfe0500f67[3] ;
            I8e591d83170c8ba46d31c61935311b22[3]  <=  I6d360540762be9eab571c0bfe0500f67[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic91f087829e0b9e0c964229a2dc567bc[4]        <=  I6d360540762be9eab571c0bfe0500f67[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I6d360540762be9eab571c0bfe0500f67[4] + 1 :
                                             I6d360540762be9eab571c0bfe0500f67[4] ;
            I8e591d83170c8ba46d31c61935311b22[4]  <=  I6d360540762be9eab571c0bfe0500f67[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic91f087829e0b9e0c964229a2dc567bc[5]        <=  I6d360540762be9eab571c0bfe0500f67[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I6d360540762be9eab571c0bfe0500f67[5] + 1 :
                                             I6d360540762be9eab571c0bfe0500f67[5] ;
            I8e591d83170c8ba46d31c61935311b22[5]  <=  I6d360540762be9eab571c0bfe0500f67[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic91f087829e0b9e0c964229a2dc567bc[6]        <=  I6d360540762be9eab571c0bfe0500f67[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I6d360540762be9eab571c0bfe0500f67[6] + 1 :
                                             I6d360540762be9eab571c0bfe0500f67[6] ;
            I8e591d83170c8ba46d31c61935311b22[6]  <=  I6d360540762be9eab571c0bfe0500f67[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic91f087829e0b9e0c964229a2dc567bc[7]        <=  I6d360540762be9eab571c0bfe0500f67[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I6d360540762be9eab571c0bfe0500f67[7] + 1 :
                                             I6d360540762be9eab571c0bfe0500f67[7] ;
            I8e591d83170c8ba46d31c61935311b22[7]  <=  I6d360540762be9eab571c0bfe0500f67[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic91f087829e0b9e0c964229a2dc567bc[8]        <=  I6d360540762be9eab571c0bfe0500f67[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I6d360540762be9eab571c0bfe0500f67[8] + 1 :
                                             I6d360540762be9eab571c0bfe0500f67[8] ;
            I8e591d83170c8ba46d31c61935311b22[8]  <=  I6d360540762be9eab571c0bfe0500f67[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic91f087829e0b9e0c964229a2dc567bc[9]        <=  I6d360540762be9eab571c0bfe0500f67[9][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I6d360540762be9eab571c0bfe0500f67[9] + 1 :
                                             I6d360540762be9eab571c0bfe0500f67[9] ;
            I8e591d83170c8ba46d31c61935311b22[9]  <=  I6d360540762be9eab571c0bfe0500f67[9][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic91f087829e0b9e0c964229a2dc567bc[10]        <=  I6d360540762be9eab571c0bfe0500f67[10][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I6d360540762be9eab571c0bfe0500f67[10] + 1 :
                                             I6d360540762be9eab571c0bfe0500f67[10] ;
            I8e591d83170c8ba46d31c61935311b22[10]  <=  I6d360540762be9eab571c0bfe0500f67[10][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic91f087829e0b9e0c964229a2dc567bc[11]        <=  I6d360540762be9eab571c0bfe0500f67[11][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I6d360540762be9eab571c0bfe0500f67[11] + 1 :
                                             I6d360540762be9eab571c0bfe0500f67[11] ;
            I8e591d83170c8ba46d31c61935311b22[11]  <=  I6d360540762be9eab571c0bfe0500f67[11][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic91f087829e0b9e0c964229a2dc567bc[12]        <=  I6d360540762be9eab571c0bfe0500f67[12][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I6d360540762be9eab571c0bfe0500f67[12] + 1 :
                                             I6d360540762be9eab571c0bfe0500f67[12] ;
            I8e591d83170c8ba46d31c61935311b22[12]  <=  I6d360540762be9eab571c0bfe0500f67[12][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0fd9bcdcf8faaaabf94649881419c66f[0]        <=  Ieb702849c7e744c5d04be8f86a00a4fa[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ieb702849c7e744c5d04be8f86a00a4fa[0] + 1 :
                                             Ieb702849c7e744c5d04be8f86a00a4fa[0] ;
            I02b62fafd371de339f299f8aefec6c43[0]  <=  Ieb702849c7e744c5d04be8f86a00a4fa[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0fd9bcdcf8faaaabf94649881419c66f[1]        <=  Ieb702849c7e744c5d04be8f86a00a4fa[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ieb702849c7e744c5d04be8f86a00a4fa[1] + 1 :
                                             Ieb702849c7e744c5d04be8f86a00a4fa[1] ;
            I02b62fafd371de339f299f8aefec6c43[1]  <=  Ieb702849c7e744c5d04be8f86a00a4fa[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0fd9bcdcf8faaaabf94649881419c66f[2]        <=  Ieb702849c7e744c5d04be8f86a00a4fa[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ieb702849c7e744c5d04be8f86a00a4fa[2] + 1 :
                                             Ieb702849c7e744c5d04be8f86a00a4fa[2] ;
            I02b62fafd371de339f299f8aefec6c43[2]  <=  Ieb702849c7e744c5d04be8f86a00a4fa[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0fd9bcdcf8faaaabf94649881419c66f[3]        <=  Ieb702849c7e744c5d04be8f86a00a4fa[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ieb702849c7e744c5d04be8f86a00a4fa[3] + 1 :
                                             Ieb702849c7e744c5d04be8f86a00a4fa[3] ;
            I02b62fafd371de339f299f8aefec6c43[3]  <=  Ieb702849c7e744c5d04be8f86a00a4fa[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0fd9bcdcf8faaaabf94649881419c66f[4]        <=  Ieb702849c7e744c5d04be8f86a00a4fa[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ieb702849c7e744c5d04be8f86a00a4fa[4] + 1 :
                                             Ieb702849c7e744c5d04be8f86a00a4fa[4] ;
            I02b62fafd371de339f299f8aefec6c43[4]  <=  Ieb702849c7e744c5d04be8f86a00a4fa[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0fd9bcdcf8faaaabf94649881419c66f[5]        <=  Ieb702849c7e744c5d04be8f86a00a4fa[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ieb702849c7e744c5d04be8f86a00a4fa[5] + 1 :
                                             Ieb702849c7e744c5d04be8f86a00a4fa[5] ;
            I02b62fafd371de339f299f8aefec6c43[5]  <=  Ieb702849c7e744c5d04be8f86a00a4fa[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0fd9bcdcf8faaaabf94649881419c66f[6]        <=  Ieb702849c7e744c5d04be8f86a00a4fa[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ieb702849c7e744c5d04be8f86a00a4fa[6] + 1 :
                                             Ieb702849c7e744c5d04be8f86a00a4fa[6] ;
            I02b62fafd371de339f299f8aefec6c43[6]  <=  Ieb702849c7e744c5d04be8f86a00a4fa[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0fd9bcdcf8faaaabf94649881419c66f[7]        <=  Ieb702849c7e744c5d04be8f86a00a4fa[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ieb702849c7e744c5d04be8f86a00a4fa[7] + 1 :
                                             Ieb702849c7e744c5d04be8f86a00a4fa[7] ;
            I02b62fafd371de339f299f8aefec6c43[7]  <=  Ieb702849c7e744c5d04be8f86a00a4fa[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0fd9bcdcf8faaaabf94649881419c66f[8]        <=  Ieb702849c7e744c5d04be8f86a00a4fa[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ieb702849c7e744c5d04be8f86a00a4fa[8] + 1 :
                                             Ieb702849c7e744c5d04be8f86a00a4fa[8] ;
            I02b62fafd371de339f299f8aefec6c43[8]  <=  Ieb702849c7e744c5d04be8f86a00a4fa[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0fd9bcdcf8faaaabf94649881419c66f[9]        <=  Ieb702849c7e744c5d04be8f86a00a4fa[9][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ieb702849c7e744c5d04be8f86a00a4fa[9] + 1 :
                                             Ieb702849c7e744c5d04be8f86a00a4fa[9] ;
            I02b62fafd371de339f299f8aefec6c43[9]  <=  Ieb702849c7e744c5d04be8f86a00a4fa[9][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0fd9bcdcf8faaaabf94649881419c66f[10]        <=  Ieb702849c7e744c5d04be8f86a00a4fa[10][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ieb702849c7e744c5d04be8f86a00a4fa[10] + 1 :
                                             Ieb702849c7e744c5d04be8f86a00a4fa[10] ;
            I02b62fafd371de339f299f8aefec6c43[10]  <=  Ieb702849c7e744c5d04be8f86a00a4fa[10][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0fd9bcdcf8faaaabf94649881419c66f[11]        <=  Ieb702849c7e744c5d04be8f86a00a4fa[11][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ieb702849c7e744c5d04be8f86a00a4fa[11] + 1 :
                                             Ieb702849c7e744c5d04be8f86a00a4fa[11] ;
            I02b62fafd371de339f299f8aefec6c43[11]  <=  Ieb702849c7e744c5d04be8f86a00a4fa[11][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0fd9bcdcf8faaaabf94649881419c66f[12]        <=  Ieb702849c7e744c5d04be8f86a00a4fa[12][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ieb702849c7e744c5d04be8f86a00a4fa[12] + 1 :
                                             Ieb702849c7e744c5d04be8f86a00a4fa[12] ;
            I02b62fafd371de339f299f8aefec6c43[12]  <=  Ieb702849c7e744c5d04be8f86a00a4fa[12][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7cbcdd5018de9ceb49554b140e5665e8[0]        <=  I8519162455bacafeb7f45c170c0b5e7e[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8519162455bacafeb7f45c170c0b5e7e[0] + 1 :
                                             I8519162455bacafeb7f45c170c0b5e7e[0] ;
            I6ebab438dc55ccf6c1600313891d9c38[0]  <=  I8519162455bacafeb7f45c170c0b5e7e[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7cbcdd5018de9ceb49554b140e5665e8[1]        <=  I8519162455bacafeb7f45c170c0b5e7e[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8519162455bacafeb7f45c170c0b5e7e[1] + 1 :
                                             I8519162455bacafeb7f45c170c0b5e7e[1] ;
            I6ebab438dc55ccf6c1600313891d9c38[1]  <=  I8519162455bacafeb7f45c170c0b5e7e[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7cbcdd5018de9ceb49554b140e5665e8[2]        <=  I8519162455bacafeb7f45c170c0b5e7e[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8519162455bacafeb7f45c170c0b5e7e[2] + 1 :
                                             I8519162455bacafeb7f45c170c0b5e7e[2] ;
            I6ebab438dc55ccf6c1600313891d9c38[2]  <=  I8519162455bacafeb7f45c170c0b5e7e[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7cbcdd5018de9ceb49554b140e5665e8[3]        <=  I8519162455bacafeb7f45c170c0b5e7e[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8519162455bacafeb7f45c170c0b5e7e[3] + 1 :
                                             I8519162455bacafeb7f45c170c0b5e7e[3] ;
            I6ebab438dc55ccf6c1600313891d9c38[3]  <=  I8519162455bacafeb7f45c170c0b5e7e[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7cbcdd5018de9ceb49554b140e5665e8[4]        <=  I8519162455bacafeb7f45c170c0b5e7e[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8519162455bacafeb7f45c170c0b5e7e[4] + 1 :
                                             I8519162455bacafeb7f45c170c0b5e7e[4] ;
            I6ebab438dc55ccf6c1600313891d9c38[4]  <=  I8519162455bacafeb7f45c170c0b5e7e[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7cbcdd5018de9ceb49554b140e5665e8[5]        <=  I8519162455bacafeb7f45c170c0b5e7e[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8519162455bacafeb7f45c170c0b5e7e[5] + 1 :
                                             I8519162455bacafeb7f45c170c0b5e7e[5] ;
            I6ebab438dc55ccf6c1600313891d9c38[5]  <=  I8519162455bacafeb7f45c170c0b5e7e[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5a79c19fd2093d974b574e85245b5617[0]        <=  I0d7c184fb7627c9c50a0026ac5052448[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I0d7c184fb7627c9c50a0026ac5052448[0] + 1 :
                                             I0d7c184fb7627c9c50a0026ac5052448[0] ;
            I2fbf89398a148c47810456812dbee5a6[0]  <=  I0d7c184fb7627c9c50a0026ac5052448[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5a79c19fd2093d974b574e85245b5617[1]        <=  I0d7c184fb7627c9c50a0026ac5052448[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I0d7c184fb7627c9c50a0026ac5052448[1] + 1 :
                                             I0d7c184fb7627c9c50a0026ac5052448[1] ;
            I2fbf89398a148c47810456812dbee5a6[1]  <=  I0d7c184fb7627c9c50a0026ac5052448[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5a79c19fd2093d974b574e85245b5617[2]        <=  I0d7c184fb7627c9c50a0026ac5052448[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I0d7c184fb7627c9c50a0026ac5052448[2] + 1 :
                                             I0d7c184fb7627c9c50a0026ac5052448[2] ;
            I2fbf89398a148c47810456812dbee5a6[2]  <=  I0d7c184fb7627c9c50a0026ac5052448[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5a79c19fd2093d974b574e85245b5617[3]        <=  I0d7c184fb7627c9c50a0026ac5052448[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I0d7c184fb7627c9c50a0026ac5052448[3] + 1 :
                                             I0d7c184fb7627c9c50a0026ac5052448[3] ;
            I2fbf89398a148c47810456812dbee5a6[3]  <=  I0d7c184fb7627c9c50a0026ac5052448[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5a79c19fd2093d974b574e85245b5617[4]        <=  I0d7c184fb7627c9c50a0026ac5052448[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I0d7c184fb7627c9c50a0026ac5052448[4] + 1 :
                                             I0d7c184fb7627c9c50a0026ac5052448[4] ;
            I2fbf89398a148c47810456812dbee5a6[4]  <=  I0d7c184fb7627c9c50a0026ac5052448[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5a79c19fd2093d974b574e85245b5617[5]        <=  I0d7c184fb7627c9c50a0026ac5052448[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I0d7c184fb7627c9c50a0026ac5052448[5] + 1 :
                                             I0d7c184fb7627c9c50a0026ac5052448[5] ;
            I2fbf89398a148c47810456812dbee5a6[5]  <=  I0d7c184fb7627c9c50a0026ac5052448[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ica937143b618734fa099683949153130[0]        <=  If5cd4834f1cb99b40cd4084fea388070[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~If5cd4834f1cb99b40cd4084fea388070[0] + 1 :
                                             If5cd4834f1cb99b40cd4084fea388070[0] ;
            Icac5a9001ee113e612e3457b4b49ee68[0]  <=  If5cd4834f1cb99b40cd4084fea388070[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ica937143b618734fa099683949153130[1]        <=  If5cd4834f1cb99b40cd4084fea388070[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~If5cd4834f1cb99b40cd4084fea388070[1] + 1 :
                                             If5cd4834f1cb99b40cd4084fea388070[1] ;
            Icac5a9001ee113e612e3457b4b49ee68[1]  <=  If5cd4834f1cb99b40cd4084fea388070[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ica937143b618734fa099683949153130[2]        <=  If5cd4834f1cb99b40cd4084fea388070[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~If5cd4834f1cb99b40cd4084fea388070[2] + 1 :
                                             If5cd4834f1cb99b40cd4084fea388070[2] ;
            Icac5a9001ee113e612e3457b4b49ee68[2]  <=  If5cd4834f1cb99b40cd4084fea388070[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ica937143b618734fa099683949153130[3]        <=  If5cd4834f1cb99b40cd4084fea388070[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~If5cd4834f1cb99b40cd4084fea388070[3] + 1 :
                                             If5cd4834f1cb99b40cd4084fea388070[3] ;
            Icac5a9001ee113e612e3457b4b49ee68[3]  <=  If5cd4834f1cb99b40cd4084fea388070[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ica937143b618734fa099683949153130[4]        <=  If5cd4834f1cb99b40cd4084fea388070[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~If5cd4834f1cb99b40cd4084fea388070[4] + 1 :
                                             If5cd4834f1cb99b40cd4084fea388070[4] ;
            Icac5a9001ee113e612e3457b4b49ee68[4]  <=  If5cd4834f1cb99b40cd4084fea388070[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ica937143b618734fa099683949153130[5]        <=  If5cd4834f1cb99b40cd4084fea388070[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~If5cd4834f1cb99b40cd4084fea388070[5] + 1 :
                                             If5cd4834f1cb99b40cd4084fea388070[5] ;
            Icac5a9001ee113e612e3457b4b49ee68[5]  <=  If5cd4834f1cb99b40cd4084fea388070[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2d4d5d2694718b39e80b89b422d690cc[0]        <=  Ia3aa64fb9d2eb1168da1f7e178c05c4e[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia3aa64fb9d2eb1168da1f7e178c05c4e[0] + 1 :
                                             Ia3aa64fb9d2eb1168da1f7e178c05c4e[0] ;
            I9461e92a5880cb9e04fcece2ef4674f0[0]  <=  Ia3aa64fb9d2eb1168da1f7e178c05c4e[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2d4d5d2694718b39e80b89b422d690cc[1]        <=  Ia3aa64fb9d2eb1168da1f7e178c05c4e[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia3aa64fb9d2eb1168da1f7e178c05c4e[1] + 1 :
                                             Ia3aa64fb9d2eb1168da1f7e178c05c4e[1] ;
            I9461e92a5880cb9e04fcece2ef4674f0[1]  <=  Ia3aa64fb9d2eb1168da1f7e178c05c4e[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2d4d5d2694718b39e80b89b422d690cc[2]        <=  Ia3aa64fb9d2eb1168da1f7e178c05c4e[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia3aa64fb9d2eb1168da1f7e178c05c4e[2] + 1 :
                                             Ia3aa64fb9d2eb1168da1f7e178c05c4e[2] ;
            I9461e92a5880cb9e04fcece2ef4674f0[2]  <=  Ia3aa64fb9d2eb1168da1f7e178c05c4e[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2d4d5d2694718b39e80b89b422d690cc[3]        <=  Ia3aa64fb9d2eb1168da1f7e178c05c4e[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia3aa64fb9d2eb1168da1f7e178c05c4e[3] + 1 :
                                             Ia3aa64fb9d2eb1168da1f7e178c05c4e[3] ;
            I9461e92a5880cb9e04fcece2ef4674f0[3]  <=  Ia3aa64fb9d2eb1168da1f7e178c05c4e[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2d4d5d2694718b39e80b89b422d690cc[4]        <=  Ia3aa64fb9d2eb1168da1f7e178c05c4e[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia3aa64fb9d2eb1168da1f7e178c05c4e[4] + 1 :
                                             Ia3aa64fb9d2eb1168da1f7e178c05c4e[4] ;
            I9461e92a5880cb9e04fcece2ef4674f0[4]  <=  Ia3aa64fb9d2eb1168da1f7e178c05c4e[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2d4d5d2694718b39e80b89b422d690cc[5]        <=  Ia3aa64fb9d2eb1168da1f7e178c05c4e[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia3aa64fb9d2eb1168da1f7e178c05c4e[5] + 1 :
                                             Ia3aa64fb9d2eb1168da1f7e178c05c4e[5] ;
            I9461e92a5880cb9e04fcece2ef4674f0[5]  <=  Ia3aa64fb9d2eb1168da1f7e178c05c4e[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic2faea3d4bb97dda16ecc29c27939ca6[0]        <=  I58c319fa3e05e8f7ca440775482ba8fe[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I58c319fa3e05e8f7ca440775482ba8fe[0] + 1 :
                                             I58c319fa3e05e8f7ca440775482ba8fe[0] ;
            I07930a807994815de45864af579902c4[0]  <=  I58c319fa3e05e8f7ca440775482ba8fe[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic2faea3d4bb97dda16ecc29c27939ca6[1]        <=  I58c319fa3e05e8f7ca440775482ba8fe[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I58c319fa3e05e8f7ca440775482ba8fe[1] + 1 :
                                             I58c319fa3e05e8f7ca440775482ba8fe[1] ;
            I07930a807994815de45864af579902c4[1]  <=  I58c319fa3e05e8f7ca440775482ba8fe[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic2faea3d4bb97dda16ecc29c27939ca6[2]        <=  I58c319fa3e05e8f7ca440775482ba8fe[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I58c319fa3e05e8f7ca440775482ba8fe[2] + 1 :
                                             I58c319fa3e05e8f7ca440775482ba8fe[2] ;
            I07930a807994815de45864af579902c4[2]  <=  I58c319fa3e05e8f7ca440775482ba8fe[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic2faea3d4bb97dda16ecc29c27939ca6[3]        <=  I58c319fa3e05e8f7ca440775482ba8fe[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I58c319fa3e05e8f7ca440775482ba8fe[3] + 1 :
                                             I58c319fa3e05e8f7ca440775482ba8fe[3] ;
            I07930a807994815de45864af579902c4[3]  <=  I58c319fa3e05e8f7ca440775482ba8fe[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic2faea3d4bb97dda16ecc29c27939ca6[4]        <=  I58c319fa3e05e8f7ca440775482ba8fe[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I58c319fa3e05e8f7ca440775482ba8fe[4] + 1 :
                                             I58c319fa3e05e8f7ca440775482ba8fe[4] ;
            I07930a807994815de45864af579902c4[4]  <=  I58c319fa3e05e8f7ca440775482ba8fe[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic2faea3d4bb97dda16ecc29c27939ca6[5]        <=  I58c319fa3e05e8f7ca440775482ba8fe[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I58c319fa3e05e8f7ca440775482ba8fe[5] + 1 :
                                             I58c319fa3e05e8f7ca440775482ba8fe[5] ;
            I07930a807994815de45864af579902c4[5]  <=  I58c319fa3e05e8f7ca440775482ba8fe[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic2faea3d4bb97dda16ecc29c27939ca6[6]        <=  I58c319fa3e05e8f7ca440775482ba8fe[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I58c319fa3e05e8f7ca440775482ba8fe[6] + 1 :
                                             I58c319fa3e05e8f7ca440775482ba8fe[6] ;
            I07930a807994815de45864af579902c4[6]  <=  I58c319fa3e05e8f7ca440775482ba8fe[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic2faea3d4bb97dda16ecc29c27939ca6[7]        <=  I58c319fa3e05e8f7ca440775482ba8fe[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I58c319fa3e05e8f7ca440775482ba8fe[7] + 1 :
                                             I58c319fa3e05e8f7ca440775482ba8fe[7] ;
            I07930a807994815de45864af579902c4[7]  <=  I58c319fa3e05e8f7ca440775482ba8fe[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I503e83a1146c42d5c1ef011ecb280807[0]        <=  I23f3a4487998f2384d9323f9103f7aca[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I23f3a4487998f2384d9323f9103f7aca[0] + 1 :
                                             I23f3a4487998f2384d9323f9103f7aca[0] ;
            I72a2f42b727a0503d43332c0f22d5ae3[0]  <=  I23f3a4487998f2384d9323f9103f7aca[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I503e83a1146c42d5c1ef011ecb280807[1]        <=  I23f3a4487998f2384d9323f9103f7aca[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I23f3a4487998f2384d9323f9103f7aca[1] + 1 :
                                             I23f3a4487998f2384d9323f9103f7aca[1] ;
            I72a2f42b727a0503d43332c0f22d5ae3[1]  <=  I23f3a4487998f2384d9323f9103f7aca[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I503e83a1146c42d5c1ef011ecb280807[2]        <=  I23f3a4487998f2384d9323f9103f7aca[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I23f3a4487998f2384d9323f9103f7aca[2] + 1 :
                                             I23f3a4487998f2384d9323f9103f7aca[2] ;
            I72a2f42b727a0503d43332c0f22d5ae3[2]  <=  I23f3a4487998f2384d9323f9103f7aca[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I503e83a1146c42d5c1ef011ecb280807[3]        <=  I23f3a4487998f2384d9323f9103f7aca[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I23f3a4487998f2384d9323f9103f7aca[3] + 1 :
                                             I23f3a4487998f2384d9323f9103f7aca[3] ;
            I72a2f42b727a0503d43332c0f22d5ae3[3]  <=  I23f3a4487998f2384d9323f9103f7aca[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I503e83a1146c42d5c1ef011ecb280807[4]        <=  I23f3a4487998f2384d9323f9103f7aca[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I23f3a4487998f2384d9323f9103f7aca[4] + 1 :
                                             I23f3a4487998f2384d9323f9103f7aca[4] ;
            I72a2f42b727a0503d43332c0f22d5ae3[4]  <=  I23f3a4487998f2384d9323f9103f7aca[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I503e83a1146c42d5c1ef011ecb280807[5]        <=  I23f3a4487998f2384d9323f9103f7aca[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I23f3a4487998f2384d9323f9103f7aca[5] + 1 :
                                             I23f3a4487998f2384d9323f9103f7aca[5] ;
            I72a2f42b727a0503d43332c0f22d5ae3[5]  <=  I23f3a4487998f2384d9323f9103f7aca[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I503e83a1146c42d5c1ef011ecb280807[6]        <=  I23f3a4487998f2384d9323f9103f7aca[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I23f3a4487998f2384d9323f9103f7aca[6] + 1 :
                                             I23f3a4487998f2384d9323f9103f7aca[6] ;
            I72a2f42b727a0503d43332c0f22d5ae3[6]  <=  I23f3a4487998f2384d9323f9103f7aca[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I503e83a1146c42d5c1ef011ecb280807[7]        <=  I23f3a4487998f2384d9323f9103f7aca[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I23f3a4487998f2384d9323f9103f7aca[7] + 1 :
                                             I23f3a4487998f2384d9323f9103f7aca[7] ;
            I72a2f42b727a0503d43332c0f22d5ae3[7]  <=  I23f3a4487998f2384d9323f9103f7aca[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib9886c1fcd27ceb24afb2d0d7da85c26[0]        <=  I081087845b5c62dc79fd5b9882339572[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I081087845b5c62dc79fd5b9882339572[0] + 1 :
                                             I081087845b5c62dc79fd5b9882339572[0] ;
            I8b8b9c4777e6df3eb2b9313e69ef2c8c[0]  <=  I081087845b5c62dc79fd5b9882339572[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib9886c1fcd27ceb24afb2d0d7da85c26[1]        <=  I081087845b5c62dc79fd5b9882339572[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I081087845b5c62dc79fd5b9882339572[1] + 1 :
                                             I081087845b5c62dc79fd5b9882339572[1] ;
            I8b8b9c4777e6df3eb2b9313e69ef2c8c[1]  <=  I081087845b5c62dc79fd5b9882339572[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib9886c1fcd27ceb24afb2d0d7da85c26[2]        <=  I081087845b5c62dc79fd5b9882339572[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I081087845b5c62dc79fd5b9882339572[2] + 1 :
                                             I081087845b5c62dc79fd5b9882339572[2] ;
            I8b8b9c4777e6df3eb2b9313e69ef2c8c[2]  <=  I081087845b5c62dc79fd5b9882339572[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib9886c1fcd27ceb24afb2d0d7da85c26[3]        <=  I081087845b5c62dc79fd5b9882339572[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I081087845b5c62dc79fd5b9882339572[3] + 1 :
                                             I081087845b5c62dc79fd5b9882339572[3] ;
            I8b8b9c4777e6df3eb2b9313e69ef2c8c[3]  <=  I081087845b5c62dc79fd5b9882339572[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib9886c1fcd27ceb24afb2d0d7da85c26[4]        <=  I081087845b5c62dc79fd5b9882339572[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I081087845b5c62dc79fd5b9882339572[4] + 1 :
                                             I081087845b5c62dc79fd5b9882339572[4] ;
            I8b8b9c4777e6df3eb2b9313e69ef2c8c[4]  <=  I081087845b5c62dc79fd5b9882339572[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib9886c1fcd27ceb24afb2d0d7da85c26[5]        <=  I081087845b5c62dc79fd5b9882339572[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I081087845b5c62dc79fd5b9882339572[5] + 1 :
                                             I081087845b5c62dc79fd5b9882339572[5] ;
            I8b8b9c4777e6df3eb2b9313e69ef2c8c[5]  <=  I081087845b5c62dc79fd5b9882339572[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib9886c1fcd27ceb24afb2d0d7da85c26[6]        <=  I081087845b5c62dc79fd5b9882339572[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I081087845b5c62dc79fd5b9882339572[6] + 1 :
                                             I081087845b5c62dc79fd5b9882339572[6] ;
            I8b8b9c4777e6df3eb2b9313e69ef2c8c[6]  <=  I081087845b5c62dc79fd5b9882339572[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib9886c1fcd27ceb24afb2d0d7da85c26[7]        <=  I081087845b5c62dc79fd5b9882339572[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I081087845b5c62dc79fd5b9882339572[7] + 1 :
                                             I081087845b5c62dc79fd5b9882339572[7] ;
            I8b8b9c4777e6df3eb2b9313e69ef2c8c[7]  <=  I081087845b5c62dc79fd5b9882339572[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Icd90612c09423a2817a72f750e585309[0]        <=  I8aa441e2ed6f41bca12ddbeaac9f5c3d[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8aa441e2ed6f41bca12ddbeaac9f5c3d[0] + 1 :
                                             I8aa441e2ed6f41bca12ddbeaac9f5c3d[0] ;
            I4a16e8e7946d9a8220304fc1be3fb362[0]  <=  I8aa441e2ed6f41bca12ddbeaac9f5c3d[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Icd90612c09423a2817a72f750e585309[1]        <=  I8aa441e2ed6f41bca12ddbeaac9f5c3d[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8aa441e2ed6f41bca12ddbeaac9f5c3d[1] + 1 :
                                             I8aa441e2ed6f41bca12ddbeaac9f5c3d[1] ;
            I4a16e8e7946d9a8220304fc1be3fb362[1]  <=  I8aa441e2ed6f41bca12ddbeaac9f5c3d[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Icd90612c09423a2817a72f750e585309[2]        <=  I8aa441e2ed6f41bca12ddbeaac9f5c3d[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8aa441e2ed6f41bca12ddbeaac9f5c3d[2] + 1 :
                                             I8aa441e2ed6f41bca12ddbeaac9f5c3d[2] ;
            I4a16e8e7946d9a8220304fc1be3fb362[2]  <=  I8aa441e2ed6f41bca12ddbeaac9f5c3d[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Icd90612c09423a2817a72f750e585309[3]        <=  I8aa441e2ed6f41bca12ddbeaac9f5c3d[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8aa441e2ed6f41bca12ddbeaac9f5c3d[3] + 1 :
                                             I8aa441e2ed6f41bca12ddbeaac9f5c3d[3] ;
            I4a16e8e7946d9a8220304fc1be3fb362[3]  <=  I8aa441e2ed6f41bca12ddbeaac9f5c3d[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Icd90612c09423a2817a72f750e585309[4]        <=  I8aa441e2ed6f41bca12ddbeaac9f5c3d[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8aa441e2ed6f41bca12ddbeaac9f5c3d[4] + 1 :
                                             I8aa441e2ed6f41bca12ddbeaac9f5c3d[4] ;
            I4a16e8e7946d9a8220304fc1be3fb362[4]  <=  I8aa441e2ed6f41bca12ddbeaac9f5c3d[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Icd90612c09423a2817a72f750e585309[5]        <=  I8aa441e2ed6f41bca12ddbeaac9f5c3d[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8aa441e2ed6f41bca12ddbeaac9f5c3d[5] + 1 :
                                             I8aa441e2ed6f41bca12ddbeaac9f5c3d[5] ;
            I4a16e8e7946d9a8220304fc1be3fb362[5]  <=  I8aa441e2ed6f41bca12ddbeaac9f5c3d[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Icd90612c09423a2817a72f750e585309[6]        <=  I8aa441e2ed6f41bca12ddbeaac9f5c3d[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8aa441e2ed6f41bca12ddbeaac9f5c3d[6] + 1 :
                                             I8aa441e2ed6f41bca12ddbeaac9f5c3d[6] ;
            I4a16e8e7946d9a8220304fc1be3fb362[6]  <=  I8aa441e2ed6f41bca12ddbeaac9f5c3d[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Icd90612c09423a2817a72f750e585309[7]        <=  I8aa441e2ed6f41bca12ddbeaac9f5c3d[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8aa441e2ed6f41bca12ddbeaac9f5c3d[7] + 1 :
                                             I8aa441e2ed6f41bca12ddbeaac9f5c3d[7] ;
            I4a16e8e7946d9a8220304fc1be3fb362[7]  <=  I8aa441e2ed6f41bca12ddbeaac9f5c3d[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib7b7884d2653893806af34579f7c0760[0]        <=  I4bc30140a67bbc7b19449fcf946a17aa[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I4bc30140a67bbc7b19449fcf946a17aa[0] + 1 :
                                             I4bc30140a67bbc7b19449fcf946a17aa[0] ;
            Ic2580cbeec8c11a19bd1e2ebc29d255e[0]  <=  I4bc30140a67bbc7b19449fcf946a17aa[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib7b7884d2653893806af34579f7c0760[1]        <=  I4bc30140a67bbc7b19449fcf946a17aa[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I4bc30140a67bbc7b19449fcf946a17aa[1] + 1 :
                                             I4bc30140a67bbc7b19449fcf946a17aa[1] ;
            Ic2580cbeec8c11a19bd1e2ebc29d255e[1]  <=  I4bc30140a67bbc7b19449fcf946a17aa[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib7b7884d2653893806af34579f7c0760[2]        <=  I4bc30140a67bbc7b19449fcf946a17aa[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I4bc30140a67bbc7b19449fcf946a17aa[2] + 1 :
                                             I4bc30140a67bbc7b19449fcf946a17aa[2] ;
            Ic2580cbeec8c11a19bd1e2ebc29d255e[2]  <=  I4bc30140a67bbc7b19449fcf946a17aa[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib7b7884d2653893806af34579f7c0760[3]        <=  I4bc30140a67bbc7b19449fcf946a17aa[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I4bc30140a67bbc7b19449fcf946a17aa[3] + 1 :
                                             I4bc30140a67bbc7b19449fcf946a17aa[3] ;
            Ic2580cbeec8c11a19bd1e2ebc29d255e[3]  <=  I4bc30140a67bbc7b19449fcf946a17aa[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib7b7884d2653893806af34579f7c0760[4]        <=  I4bc30140a67bbc7b19449fcf946a17aa[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I4bc30140a67bbc7b19449fcf946a17aa[4] + 1 :
                                             I4bc30140a67bbc7b19449fcf946a17aa[4] ;
            Ic2580cbeec8c11a19bd1e2ebc29d255e[4]  <=  I4bc30140a67bbc7b19449fcf946a17aa[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib7b7884d2653893806af34579f7c0760[5]        <=  I4bc30140a67bbc7b19449fcf946a17aa[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I4bc30140a67bbc7b19449fcf946a17aa[5] + 1 :
                                             I4bc30140a67bbc7b19449fcf946a17aa[5] ;
            Ic2580cbeec8c11a19bd1e2ebc29d255e[5]  <=  I4bc30140a67bbc7b19449fcf946a17aa[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib7b7884d2653893806af34579f7c0760[6]        <=  I4bc30140a67bbc7b19449fcf946a17aa[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I4bc30140a67bbc7b19449fcf946a17aa[6] + 1 :
                                             I4bc30140a67bbc7b19449fcf946a17aa[6] ;
            Ic2580cbeec8c11a19bd1e2ebc29d255e[6]  <=  I4bc30140a67bbc7b19449fcf946a17aa[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib7b7884d2653893806af34579f7c0760[7]        <=  I4bc30140a67bbc7b19449fcf946a17aa[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I4bc30140a67bbc7b19449fcf946a17aa[7] + 1 :
                                             I4bc30140a67bbc7b19449fcf946a17aa[7] ;
            Ic2580cbeec8c11a19bd1e2ebc29d255e[7]  <=  I4bc30140a67bbc7b19449fcf946a17aa[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib7b7884d2653893806af34579f7c0760[8]        <=  I4bc30140a67bbc7b19449fcf946a17aa[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I4bc30140a67bbc7b19449fcf946a17aa[8] + 1 :
                                             I4bc30140a67bbc7b19449fcf946a17aa[8] ;
            Ic2580cbeec8c11a19bd1e2ebc29d255e[8]  <=  I4bc30140a67bbc7b19449fcf946a17aa[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic3f0ad21d8a446c31afec49309a18133[0]        <=  I943f523a14e49f42d9c6ceb3ad1dd841[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I943f523a14e49f42d9c6ceb3ad1dd841[0] + 1 :
                                             I943f523a14e49f42d9c6ceb3ad1dd841[0] ;
            If79ed5ee2b8710da0608c1e245d07d55[0]  <=  I943f523a14e49f42d9c6ceb3ad1dd841[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic3f0ad21d8a446c31afec49309a18133[1]        <=  I943f523a14e49f42d9c6ceb3ad1dd841[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I943f523a14e49f42d9c6ceb3ad1dd841[1] + 1 :
                                             I943f523a14e49f42d9c6ceb3ad1dd841[1] ;
            If79ed5ee2b8710da0608c1e245d07d55[1]  <=  I943f523a14e49f42d9c6ceb3ad1dd841[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic3f0ad21d8a446c31afec49309a18133[2]        <=  I943f523a14e49f42d9c6ceb3ad1dd841[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I943f523a14e49f42d9c6ceb3ad1dd841[2] + 1 :
                                             I943f523a14e49f42d9c6ceb3ad1dd841[2] ;
            If79ed5ee2b8710da0608c1e245d07d55[2]  <=  I943f523a14e49f42d9c6ceb3ad1dd841[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic3f0ad21d8a446c31afec49309a18133[3]        <=  I943f523a14e49f42d9c6ceb3ad1dd841[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I943f523a14e49f42d9c6ceb3ad1dd841[3] + 1 :
                                             I943f523a14e49f42d9c6ceb3ad1dd841[3] ;
            If79ed5ee2b8710da0608c1e245d07d55[3]  <=  I943f523a14e49f42d9c6ceb3ad1dd841[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic3f0ad21d8a446c31afec49309a18133[4]        <=  I943f523a14e49f42d9c6ceb3ad1dd841[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I943f523a14e49f42d9c6ceb3ad1dd841[4] + 1 :
                                             I943f523a14e49f42d9c6ceb3ad1dd841[4] ;
            If79ed5ee2b8710da0608c1e245d07d55[4]  <=  I943f523a14e49f42d9c6ceb3ad1dd841[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic3f0ad21d8a446c31afec49309a18133[5]        <=  I943f523a14e49f42d9c6ceb3ad1dd841[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I943f523a14e49f42d9c6ceb3ad1dd841[5] + 1 :
                                             I943f523a14e49f42d9c6ceb3ad1dd841[5] ;
            If79ed5ee2b8710da0608c1e245d07d55[5]  <=  I943f523a14e49f42d9c6ceb3ad1dd841[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic3f0ad21d8a446c31afec49309a18133[6]        <=  I943f523a14e49f42d9c6ceb3ad1dd841[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I943f523a14e49f42d9c6ceb3ad1dd841[6] + 1 :
                                             I943f523a14e49f42d9c6ceb3ad1dd841[6] ;
            If79ed5ee2b8710da0608c1e245d07d55[6]  <=  I943f523a14e49f42d9c6ceb3ad1dd841[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic3f0ad21d8a446c31afec49309a18133[7]        <=  I943f523a14e49f42d9c6ceb3ad1dd841[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I943f523a14e49f42d9c6ceb3ad1dd841[7] + 1 :
                                             I943f523a14e49f42d9c6ceb3ad1dd841[7] ;
            If79ed5ee2b8710da0608c1e245d07d55[7]  <=  I943f523a14e49f42d9c6ceb3ad1dd841[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic3f0ad21d8a446c31afec49309a18133[8]        <=  I943f523a14e49f42d9c6ceb3ad1dd841[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I943f523a14e49f42d9c6ceb3ad1dd841[8] + 1 :
                                             I943f523a14e49f42d9c6ceb3ad1dd841[8] ;
            If79ed5ee2b8710da0608c1e245d07d55[8]  <=  I943f523a14e49f42d9c6ceb3ad1dd841[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2dd65bec7d2bc4778b7fc48a413d2ba7[0]        <=  I10ab80965b99680e93ea304f6e261094[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I10ab80965b99680e93ea304f6e261094[0] + 1 :
                                             I10ab80965b99680e93ea304f6e261094[0] ;
            I9497bbb4f746969a95cff948a3ee9ade[0]  <=  I10ab80965b99680e93ea304f6e261094[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2dd65bec7d2bc4778b7fc48a413d2ba7[1]        <=  I10ab80965b99680e93ea304f6e261094[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I10ab80965b99680e93ea304f6e261094[1] + 1 :
                                             I10ab80965b99680e93ea304f6e261094[1] ;
            I9497bbb4f746969a95cff948a3ee9ade[1]  <=  I10ab80965b99680e93ea304f6e261094[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2dd65bec7d2bc4778b7fc48a413d2ba7[2]        <=  I10ab80965b99680e93ea304f6e261094[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I10ab80965b99680e93ea304f6e261094[2] + 1 :
                                             I10ab80965b99680e93ea304f6e261094[2] ;
            I9497bbb4f746969a95cff948a3ee9ade[2]  <=  I10ab80965b99680e93ea304f6e261094[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2dd65bec7d2bc4778b7fc48a413d2ba7[3]        <=  I10ab80965b99680e93ea304f6e261094[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I10ab80965b99680e93ea304f6e261094[3] + 1 :
                                             I10ab80965b99680e93ea304f6e261094[3] ;
            I9497bbb4f746969a95cff948a3ee9ade[3]  <=  I10ab80965b99680e93ea304f6e261094[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2dd65bec7d2bc4778b7fc48a413d2ba7[4]        <=  I10ab80965b99680e93ea304f6e261094[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I10ab80965b99680e93ea304f6e261094[4] + 1 :
                                             I10ab80965b99680e93ea304f6e261094[4] ;
            I9497bbb4f746969a95cff948a3ee9ade[4]  <=  I10ab80965b99680e93ea304f6e261094[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2dd65bec7d2bc4778b7fc48a413d2ba7[5]        <=  I10ab80965b99680e93ea304f6e261094[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I10ab80965b99680e93ea304f6e261094[5] + 1 :
                                             I10ab80965b99680e93ea304f6e261094[5] ;
            I9497bbb4f746969a95cff948a3ee9ade[5]  <=  I10ab80965b99680e93ea304f6e261094[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2dd65bec7d2bc4778b7fc48a413d2ba7[6]        <=  I10ab80965b99680e93ea304f6e261094[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I10ab80965b99680e93ea304f6e261094[6] + 1 :
                                             I10ab80965b99680e93ea304f6e261094[6] ;
            I9497bbb4f746969a95cff948a3ee9ade[6]  <=  I10ab80965b99680e93ea304f6e261094[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2dd65bec7d2bc4778b7fc48a413d2ba7[7]        <=  I10ab80965b99680e93ea304f6e261094[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I10ab80965b99680e93ea304f6e261094[7] + 1 :
                                             I10ab80965b99680e93ea304f6e261094[7] ;
            I9497bbb4f746969a95cff948a3ee9ade[7]  <=  I10ab80965b99680e93ea304f6e261094[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2dd65bec7d2bc4778b7fc48a413d2ba7[8]        <=  I10ab80965b99680e93ea304f6e261094[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I10ab80965b99680e93ea304f6e261094[8] + 1 :
                                             I10ab80965b99680e93ea304f6e261094[8] ;
            I9497bbb4f746969a95cff948a3ee9ade[8]  <=  I10ab80965b99680e93ea304f6e261094[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I36b5867a3da6f2ed529e791166640d3f[0]        <=  Ibfef15cf57c5850241c05384f18da5ea[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ibfef15cf57c5850241c05384f18da5ea[0] + 1 :
                                             Ibfef15cf57c5850241c05384f18da5ea[0] ;
            I651d700a00d7004d8728bc7356f30926[0]  <=  Ibfef15cf57c5850241c05384f18da5ea[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I36b5867a3da6f2ed529e791166640d3f[1]        <=  Ibfef15cf57c5850241c05384f18da5ea[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ibfef15cf57c5850241c05384f18da5ea[1] + 1 :
                                             Ibfef15cf57c5850241c05384f18da5ea[1] ;
            I651d700a00d7004d8728bc7356f30926[1]  <=  Ibfef15cf57c5850241c05384f18da5ea[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I36b5867a3da6f2ed529e791166640d3f[2]        <=  Ibfef15cf57c5850241c05384f18da5ea[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ibfef15cf57c5850241c05384f18da5ea[2] + 1 :
                                             Ibfef15cf57c5850241c05384f18da5ea[2] ;
            I651d700a00d7004d8728bc7356f30926[2]  <=  Ibfef15cf57c5850241c05384f18da5ea[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I36b5867a3da6f2ed529e791166640d3f[3]        <=  Ibfef15cf57c5850241c05384f18da5ea[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ibfef15cf57c5850241c05384f18da5ea[3] + 1 :
                                             Ibfef15cf57c5850241c05384f18da5ea[3] ;
            I651d700a00d7004d8728bc7356f30926[3]  <=  Ibfef15cf57c5850241c05384f18da5ea[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I36b5867a3da6f2ed529e791166640d3f[4]        <=  Ibfef15cf57c5850241c05384f18da5ea[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ibfef15cf57c5850241c05384f18da5ea[4] + 1 :
                                             Ibfef15cf57c5850241c05384f18da5ea[4] ;
            I651d700a00d7004d8728bc7356f30926[4]  <=  Ibfef15cf57c5850241c05384f18da5ea[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I36b5867a3da6f2ed529e791166640d3f[5]        <=  Ibfef15cf57c5850241c05384f18da5ea[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ibfef15cf57c5850241c05384f18da5ea[5] + 1 :
                                             Ibfef15cf57c5850241c05384f18da5ea[5] ;
            I651d700a00d7004d8728bc7356f30926[5]  <=  Ibfef15cf57c5850241c05384f18da5ea[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I36b5867a3da6f2ed529e791166640d3f[6]        <=  Ibfef15cf57c5850241c05384f18da5ea[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ibfef15cf57c5850241c05384f18da5ea[6] + 1 :
                                             Ibfef15cf57c5850241c05384f18da5ea[6] ;
            I651d700a00d7004d8728bc7356f30926[6]  <=  Ibfef15cf57c5850241c05384f18da5ea[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I36b5867a3da6f2ed529e791166640d3f[7]        <=  Ibfef15cf57c5850241c05384f18da5ea[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ibfef15cf57c5850241c05384f18da5ea[7] + 1 :
                                             Ibfef15cf57c5850241c05384f18da5ea[7] ;
            I651d700a00d7004d8728bc7356f30926[7]  <=  Ibfef15cf57c5850241c05384f18da5ea[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I36b5867a3da6f2ed529e791166640d3f[8]        <=  Ibfef15cf57c5850241c05384f18da5ea[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ibfef15cf57c5850241c05384f18da5ea[8] + 1 :
                                             Ibfef15cf57c5850241c05384f18da5ea[8] ;
            I651d700a00d7004d8728bc7356f30926[8]  <=  Ibfef15cf57c5850241c05384f18da5ea[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iedc20522d3322bbe3f55e2aa611d76df[0]        <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I0aa8bcd235f4c4f32c3075d5f39bc20f[0] + 1 :
                                             I0aa8bcd235f4c4f32c3075d5f39bc20f[0] ;
            I6f5c991e5fdcf56d582c6f80eb6731df[0]  <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iedc20522d3322bbe3f55e2aa611d76df[1]        <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I0aa8bcd235f4c4f32c3075d5f39bc20f[1] + 1 :
                                             I0aa8bcd235f4c4f32c3075d5f39bc20f[1] ;
            I6f5c991e5fdcf56d582c6f80eb6731df[1]  <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iedc20522d3322bbe3f55e2aa611d76df[2]        <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I0aa8bcd235f4c4f32c3075d5f39bc20f[2] + 1 :
                                             I0aa8bcd235f4c4f32c3075d5f39bc20f[2] ;
            I6f5c991e5fdcf56d582c6f80eb6731df[2]  <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iedc20522d3322bbe3f55e2aa611d76df[3]        <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I0aa8bcd235f4c4f32c3075d5f39bc20f[3] + 1 :
                                             I0aa8bcd235f4c4f32c3075d5f39bc20f[3] ;
            I6f5c991e5fdcf56d582c6f80eb6731df[3]  <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iedc20522d3322bbe3f55e2aa611d76df[4]        <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I0aa8bcd235f4c4f32c3075d5f39bc20f[4] + 1 :
                                             I0aa8bcd235f4c4f32c3075d5f39bc20f[4] ;
            I6f5c991e5fdcf56d582c6f80eb6731df[4]  <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iedc20522d3322bbe3f55e2aa611d76df[5]        <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I0aa8bcd235f4c4f32c3075d5f39bc20f[5] + 1 :
                                             I0aa8bcd235f4c4f32c3075d5f39bc20f[5] ;
            I6f5c991e5fdcf56d582c6f80eb6731df[5]  <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iedc20522d3322bbe3f55e2aa611d76df[6]        <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I0aa8bcd235f4c4f32c3075d5f39bc20f[6] + 1 :
                                             I0aa8bcd235f4c4f32c3075d5f39bc20f[6] ;
            I6f5c991e5fdcf56d582c6f80eb6731df[6]  <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iedc20522d3322bbe3f55e2aa611d76df[7]        <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I0aa8bcd235f4c4f32c3075d5f39bc20f[7] + 1 :
                                             I0aa8bcd235f4c4f32c3075d5f39bc20f[7] ;
            I6f5c991e5fdcf56d582c6f80eb6731df[7]  <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iedc20522d3322bbe3f55e2aa611d76df[8]        <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I0aa8bcd235f4c4f32c3075d5f39bc20f[8] + 1 :
                                             I0aa8bcd235f4c4f32c3075d5f39bc20f[8] ;
            I6f5c991e5fdcf56d582c6f80eb6731df[8]  <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iedc20522d3322bbe3f55e2aa611d76df[9]        <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[9][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I0aa8bcd235f4c4f32c3075d5f39bc20f[9] + 1 :
                                             I0aa8bcd235f4c4f32c3075d5f39bc20f[9] ;
            I6f5c991e5fdcf56d582c6f80eb6731df[9]  <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[9][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iedc20522d3322bbe3f55e2aa611d76df[10]        <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[10][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I0aa8bcd235f4c4f32c3075d5f39bc20f[10] + 1 :
                                             I0aa8bcd235f4c4f32c3075d5f39bc20f[10] ;
            I6f5c991e5fdcf56d582c6f80eb6731df[10]  <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[10][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iedc20522d3322bbe3f55e2aa611d76df[11]        <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[11][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I0aa8bcd235f4c4f32c3075d5f39bc20f[11] + 1 :
                                             I0aa8bcd235f4c4f32c3075d5f39bc20f[11] ;
            I6f5c991e5fdcf56d582c6f80eb6731df[11]  <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[11][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iedc20522d3322bbe3f55e2aa611d76df[12]        <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[12][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I0aa8bcd235f4c4f32c3075d5f39bc20f[12] + 1 :
                                             I0aa8bcd235f4c4f32c3075d5f39bc20f[12] ;
            I6f5c991e5fdcf56d582c6f80eb6731df[12]  <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[12][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iedc20522d3322bbe3f55e2aa611d76df[13]        <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[13][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I0aa8bcd235f4c4f32c3075d5f39bc20f[13] + 1 :
                                             I0aa8bcd235f4c4f32c3075d5f39bc20f[13] ;
            I6f5c991e5fdcf56d582c6f80eb6731df[13]  <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[13][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iedc20522d3322bbe3f55e2aa611d76df[14]        <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[14][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I0aa8bcd235f4c4f32c3075d5f39bc20f[14] + 1 :
                                             I0aa8bcd235f4c4f32c3075d5f39bc20f[14] ;
            I6f5c991e5fdcf56d582c6f80eb6731df[14]  <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[14][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iedc20522d3322bbe3f55e2aa611d76df[15]        <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[15][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I0aa8bcd235f4c4f32c3075d5f39bc20f[15] + 1 :
                                             I0aa8bcd235f4c4f32c3075d5f39bc20f[15] ;
            I6f5c991e5fdcf56d582c6f80eb6731df[15]  <=  I0aa8bcd235f4c4f32c3075d5f39bc20f[15][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6821e897aea31f7c237ca1a553bf0cd1[0]        <=  Ic5e951c3193081b1880ccf868e740e92[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic5e951c3193081b1880ccf868e740e92[0] + 1 :
                                             Ic5e951c3193081b1880ccf868e740e92[0] ;
            Ia5cc3055ba3365e64cf59c4d4fd3f093[0]  <=  Ic5e951c3193081b1880ccf868e740e92[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6821e897aea31f7c237ca1a553bf0cd1[1]        <=  Ic5e951c3193081b1880ccf868e740e92[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic5e951c3193081b1880ccf868e740e92[1] + 1 :
                                             Ic5e951c3193081b1880ccf868e740e92[1] ;
            Ia5cc3055ba3365e64cf59c4d4fd3f093[1]  <=  Ic5e951c3193081b1880ccf868e740e92[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6821e897aea31f7c237ca1a553bf0cd1[2]        <=  Ic5e951c3193081b1880ccf868e740e92[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic5e951c3193081b1880ccf868e740e92[2] + 1 :
                                             Ic5e951c3193081b1880ccf868e740e92[2] ;
            Ia5cc3055ba3365e64cf59c4d4fd3f093[2]  <=  Ic5e951c3193081b1880ccf868e740e92[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6821e897aea31f7c237ca1a553bf0cd1[3]        <=  Ic5e951c3193081b1880ccf868e740e92[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic5e951c3193081b1880ccf868e740e92[3] + 1 :
                                             Ic5e951c3193081b1880ccf868e740e92[3] ;
            Ia5cc3055ba3365e64cf59c4d4fd3f093[3]  <=  Ic5e951c3193081b1880ccf868e740e92[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6821e897aea31f7c237ca1a553bf0cd1[4]        <=  Ic5e951c3193081b1880ccf868e740e92[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic5e951c3193081b1880ccf868e740e92[4] + 1 :
                                             Ic5e951c3193081b1880ccf868e740e92[4] ;
            Ia5cc3055ba3365e64cf59c4d4fd3f093[4]  <=  Ic5e951c3193081b1880ccf868e740e92[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6821e897aea31f7c237ca1a553bf0cd1[5]        <=  Ic5e951c3193081b1880ccf868e740e92[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic5e951c3193081b1880ccf868e740e92[5] + 1 :
                                             Ic5e951c3193081b1880ccf868e740e92[5] ;
            Ia5cc3055ba3365e64cf59c4d4fd3f093[5]  <=  Ic5e951c3193081b1880ccf868e740e92[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6821e897aea31f7c237ca1a553bf0cd1[6]        <=  Ic5e951c3193081b1880ccf868e740e92[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic5e951c3193081b1880ccf868e740e92[6] + 1 :
                                             Ic5e951c3193081b1880ccf868e740e92[6] ;
            Ia5cc3055ba3365e64cf59c4d4fd3f093[6]  <=  Ic5e951c3193081b1880ccf868e740e92[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6821e897aea31f7c237ca1a553bf0cd1[7]        <=  Ic5e951c3193081b1880ccf868e740e92[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic5e951c3193081b1880ccf868e740e92[7] + 1 :
                                             Ic5e951c3193081b1880ccf868e740e92[7] ;
            Ia5cc3055ba3365e64cf59c4d4fd3f093[7]  <=  Ic5e951c3193081b1880ccf868e740e92[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6821e897aea31f7c237ca1a553bf0cd1[8]        <=  Ic5e951c3193081b1880ccf868e740e92[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic5e951c3193081b1880ccf868e740e92[8] + 1 :
                                             Ic5e951c3193081b1880ccf868e740e92[8] ;
            Ia5cc3055ba3365e64cf59c4d4fd3f093[8]  <=  Ic5e951c3193081b1880ccf868e740e92[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6821e897aea31f7c237ca1a553bf0cd1[9]        <=  Ic5e951c3193081b1880ccf868e740e92[9][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic5e951c3193081b1880ccf868e740e92[9] + 1 :
                                             Ic5e951c3193081b1880ccf868e740e92[9] ;
            Ia5cc3055ba3365e64cf59c4d4fd3f093[9]  <=  Ic5e951c3193081b1880ccf868e740e92[9][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6821e897aea31f7c237ca1a553bf0cd1[10]        <=  Ic5e951c3193081b1880ccf868e740e92[10][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic5e951c3193081b1880ccf868e740e92[10] + 1 :
                                             Ic5e951c3193081b1880ccf868e740e92[10] ;
            Ia5cc3055ba3365e64cf59c4d4fd3f093[10]  <=  Ic5e951c3193081b1880ccf868e740e92[10][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6821e897aea31f7c237ca1a553bf0cd1[11]        <=  Ic5e951c3193081b1880ccf868e740e92[11][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic5e951c3193081b1880ccf868e740e92[11] + 1 :
                                             Ic5e951c3193081b1880ccf868e740e92[11] ;
            Ia5cc3055ba3365e64cf59c4d4fd3f093[11]  <=  Ic5e951c3193081b1880ccf868e740e92[11][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6821e897aea31f7c237ca1a553bf0cd1[12]        <=  Ic5e951c3193081b1880ccf868e740e92[12][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic5e951c3193081b1880ccf868e740e92[12] + 1 :
                                             Ic5e951c3193081b1880ccf868e740e92[12] ;
            Ia5cc3055ba3365e64cf59c4d4fd3f093[12]  <=  Ic5e951c3193081b1880ccf868e740e92[12][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6821e897aea31f7c237ca1a553bf0cd1[13]        <=  Ic5e951c3193081b1880ccf868e740e92[13][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic5e951c3193081b1880ccf868e740e92[13] + 1 :
                                             Ic5e951c3193081b1880ccf868e740e92[13] ;
            Ia5cc3055ba3365e64cf59c4d4fd3f093[13]  <=  Ic5e951c3193081b1880ccf868e740e92[13][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6821e897aea31f7c237ca1a553bf0cd1[14]        <=  Ic5e951c3193081b1880ccf868e740e92[14][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic5e951c3193081b1880ccf868e740e92[14] + 1 :
                                             Ic5e951c3193081b1880ccf868e740e92[14] ;
            Ia5cc3055ba3365e64cf59c4d4fd3f093[14]  <=  Ic5e951c3193081b1880ccf868e740e92[14][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6821e897aea31f7c237ca1a553bf0cd1[15]        <=  Ic5e951c3193081b1880ccf868e740e92[15][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic5e951c3193081b1880ccf868e740e92[15] + 1 :
                                             Ic5e951c3193081b1880ccf868e740e92[15] ;
            Ia5cc3055ba3365e64cf59c4d4fd3f093[15]  <=  Ic5e951c3193081b1880ccf868e740e92[15][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I290499340d94dd8e234f53f9962a182b[0]        <=  Ie8edae9436451bc0a4dbdbf531401682[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie8edae9436451bc0a4dbdbf531401682[0] + 1 :
                                             Ie8edae9436451bc0a4dbdbf531401682[0] ;
            Iea7da1f43ba202d753b0edb0be8b3fcf[0]  <=  Ie8edae9436451bc0a4dbdbf531401682[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I290499340d94dd8e234f53f9962a182b[1]        <=  Ie8edae9436451bc0a4dbdbf531401682[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie8edae9436451bc0a4dbdbf531401682[1] + 1 :
                                             Ie8edae9436451bc0a4dbdbf531401682[1] ;
            Iea7da1f43ba202d753b0edb0be8b3fcf[1]  <=  Ie8edae9436451bc0a4dbdbf531401682[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I290499340d94dd8e234f53f9962a182b[2]        <=  Ie8edae9436451bc0a4dbdbf531401682[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie8edae9436451bc0a4dbdbf531401682[2] + 1 :
                                             Ie8edae9436451bc0a4dbdbf531401682[2] ;
            Iea7da1f43ba202d753b0edb0be8b3fcf[2]  <=  Ie8edae9436451bc0a4dbdbf531401682[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I290499340d94dd8e234f53f9962a182b[3]        <=  Ie8edae9436451bc0a4dbdbf531401682[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie8edae9436451bc0a4dbdbf531401682[3] + 1 :
                                             Ie8edae9436451bc0a4dbdbf531401682[3] ;
            Iea7da1f43ba202d753b0edb0be8b3fcf[3]  <=  Ie8edae9436451bc0a4dbdbf531401682[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I290499340d94dd8e234f53f9962a182b[4]        <=  Ie8edae9436451bc0a4dbdbf531401682[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie8edae9436451bc0a4dbdbf531401682[4] + 1 :
                                             Ie8edae9436451bc0a4dbdbf531401682[4] ;
            Iea7da1f43ba202d753b0edb0be8b3fcf[4]  <=  Ie8edae9436451bc0a4dbdbf531401682[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I290499340d94dd8e234f53f9962a182b[5]        <=  Ie8edae9436451bc0a4dbdbf531401682[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie8edae9436451bc0a4dbdbf531401682[5] + 1 :
                                             Ie8edae9436451bc0a4dbdbf531401682[5] ;
            Iea7da1f43ba202d753b0edb0be8b3fcf[5]  <=  Ie8edae9436451bc0a4dbdbf531401682[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I290499340d94dd8e234f53f9962a182b[6]        <=  Ie8edae9436451bc0a4dbdbf531401682[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie8edae9436451bc0a4dbdbf531401682[6] + 1 :
                                             Ie8edae9436451bc0a4dbdbf531401682[6] ;
            Iea7da1f43ba202d753b0edb0be8b3fcf[6]  <=  Ie8edae9436451bc0a4dbdbf531401682[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I290499340d94dd8e234f53f9962a182b[7]        <=  Ie8edae9436451bc0a4dbdbf531401682[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie8edae9436451bc0a4dbdbf531401682[7] + 1 :
                                             Ie8edae9436451bc0a4dbdbf531401682[7] ;
            Iea7da1f43ba202d753b0edb0be8b3fcf[7]  <=  Ie8edae9436451bc0a4dbdbf531401682[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I290499340d94dd8e234f53f9962a182b[8]        <=  Ie8edae9436451bc0a4dbdbf531401682[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie8edae9436451bc0a4dbdbf531401682[8] + 1 :
                                             Ie8edae9436451bc0a4dbdbf531401682[8] ;
            Iea7da1f43ba202d753b0edb0be8b3fcf[8]  <=  Ie8edae9436451bc0a4dbdbf531401682[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I290499340d94dd8e234f53f9962a182b[9]        <=  Ie8edae9436451bc0a4dbdbf531401682[9][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie8edae9436451bc0a4dbdbf531401682[9] + 1 :
                                             Ie8edae9436451bc0a4dbdbf531401682[9] ;
            Iea7da1f43ba202d753b0edb0be8b3fcf[9]  <=  Ie8edae9436451bc0a4dbdbf531401682[9][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I290499340d94dd8e234f53f9962a182b[10]        <=  Ie8edae9436451bc0a4dbdbf531401682[10][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie8edae9436451bc0a4dbdbf531401682[10] + 1 :
                                             Ie8edae9436451bc0a4dbdbf531401682[10] ;
            Iea7da1f43ba202d753b0edb0be8b3fcf[10]  <=  Ie8edae9436451bc0a4dbdbf531401682[10][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I290499340d94dd8e234f53f9962a182b[11]        <=  Ie8edae9436451bc0a4dbdbf531401682[11][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie8edae9436451bc0a4dbdbf531401682[11] + 1 :
                                             Ie8edae9436451bc0a4dbdbf531401682[11] ;
            Iea7da1f43ba202d753b0edb0be8b3fcf[11]  <=  Ie8edae9436451bc0a4dbdbf531401682[11][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I290499340d94dd8e234f53f9962a182b[12]        <=  Ie8edae9436451bc0a4dbdbf531401682[12][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie8edae9436451bc0a4dbdbf531401682[12] + 1 :
                                             Ie8edae9436451bc0a4dbdbf531401682[12] ;
            Iea7da1f43ba202d753b0edb0be8b3fcf[12]  <=  Ie8edae9436451bc0a4dbdbf531401682[12][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I290499340d94dd8e234f53f9962a182b[13]        <=  Ie8edae9436451bc0a4dbdbf531401682[13][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie8edae9436451bc0a4dbdbf531401682[13] + 1 :
                                             Ie8edae9436451bc0a4dbdbf531401682[13] ;
            Iea7da1f43ba202d753b0edb0be8b3fcf[13]  <=  Ie8edae9436451bc0a4dbdbf531401682[13][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I290499340d94dd8e234f53f9962a182b[14]        <=  Ie8edae9436451bc0a4dbdbf531401682[14][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie8edae9436451bc0a4dbdbf531401682[14] + 1 :
                                             Ie8edae9436451bc0a4dbdbf531401682[14] ;
            Iea7da1f43ba202d753b0edb0be8b3fcf[14]  <=  Ie8edae9436451bc0a4dbdbf531401682[14][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I290499340d94dd8e234f53f9962a182b[15]        <=  Ie8edae9436451bc0a4dbdbf531401682[15][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie8edae9436451bc0a4dbdbf531401682[15] + 1 :
                                             Ie8edae9436451bc0a4dbdbf531401682[15] ;
            Iea7da1f43ba202d753b0edb0be8b3fcf[15]  <=  Ie8edae9436451bc0a4dbdbf531401682[15][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5ce387684404cf922955e4af33ed2367[0]        <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I84a56b9dce9dfafc97fbdc2ad3b2ae68[0] + 1 :
                                             I84a56b9dce9dfafc97fbdc2ad3b2ae68[0] ;
            I872f61d20baf011e867b44dc5539fc37[0]  <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5ce387684404cf922955e4af33ed2367[1]        <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I84a56b9dce9dfafc97fbdc2ad3b2ae68[1] + 1 :
                                             I84a56b9dce9dfafc97fbdc2ad3b2ae68[1] ;
            I872f61d20baf011e867b44dc5539fc37[1]  <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5ce387684404cf922955e4af33ed2367[2]        <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I84a56b9dce9dfafc97fbdc2ad3b2ae68[2] + 1 :
                                             I84a56b9dce9dfafc97fbdc2ad3b2ae68[2] ;
            I872f61d20baf011e867b44dc5539fc37[2]  <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5ce387684404cf922955e4af33ed2367[3]        <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I84a56b9dce9dfafc97fbdc2ad3b2ae68[3] + 1 :
                                             I84a56b9dce9dfafc97fbdc2ad3b2ae68[3] ;
            I872f61d20baf011e867b44dc5539fc37[3]  <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5ce387684404cf922955e4af33ed2367[4]        <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I84a56b9dce9dfafc97fbdc2ad3b2ae68[4] + 1 :
                                             I84a56b9dce9dfafc97fbdc2ad3b2ae68[4] ;
            I872f61d20baf011e867b44dc5539fc37[4]  <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5ce387684404cf922955e4af33ed2367[5]        <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I84a56b9dce9dfafc97fbdc2ad3b2ae68[5] + 1 :
                                             I84a56b9dce9dfafc97fbdc2ad3b2ae68[5] ;
            I872f61d20baf011e867b44dc5539fc37[5]  <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5ce387684404cf922955e4af33ed2367[6]        <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I84a56b9dce9dfafc97fbdc2ad3b2ae68[6] + 1 :
                                             I84a56b9dce9dfafc97fbdc2ad3b2ae68[6] ;
            I872f61d20baf011e867b44dc5539fc37[6]  <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5ce387684404cf922955e4af33ed2367[7]        <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I84a56b9dce9dfafc97fbdc2ad3b2ae68[7] + 1 :
                                             I84a56b9dce9dfafc97fbdc2ad3b2ae68[7] ;
            I872f61d20baf011e867b44dc5539fc37[7]  <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5ce387684404cf922955e4af33ed2367[8]        <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I84a56b9dce9dfafc97fbdc2ad3b2ae68[8] + 1 :
                                             I84a56b9dce9dfafc97fbdc2ad3b2ae68[8] ;
            I872f61d20baf011e867b44dc5539fc37[8]  <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5ce387684404cf922955e4af33ed2367[9]        <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[9][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I84a56b9dce9dfafc97fbdc2ad3b2ae68[9] + 1 :
                                             I84a56b9dce9dfafc97fbdc2ad3b2ae68[9] ;
            I872f61d20baf011e867b44dc5539fc37[9]  <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[9][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5ce387684404cf922955e4af33ed2367[10]        <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[10][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I84a56b9dce9dfafc97fbdc2ad3b2ae68[10] + 1 :
                                             I84a56b9dce9dfafc97fbdc2ad3b2ae68[10] ;
            I872f61d20baf011e867b44dc5539fc37[10]  <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[10][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5ce387684404cf922955e4af33ed2367[11]        <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[11][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I84a56b9dce9dfafc97fbdc2ad3b2ae68[11] + 1 :
                                             I84a56b9dce9dfafc97fbdc2ad3b2ae68[11] ;
            I872f61d20baf011e867b44dc5539fc37[11]  <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[11][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5ce387684404cf922955e4af33ed2367[12]        <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[12][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I84a56b9dce9dfafc97fbdc2ad3b2ae68[12] + 1 :
                                             I84a56b9dce9dfafc97fbdc2ad3b2ae68[12] ;
            I872f61d20baf011e867b44dc5539fc37[12]  <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[12][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5ce387684404cf922955e4af33ed2367[13]        <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[13][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I84a56b9dce9dfafc97fbdc2ad3b2ae68[13] + 1 :
                                             I84a56b9dce9dfafc97fbdc2ad3b2ae68[13] ;
            I872f61d20baf011e867b44dc5539fc37[13]  <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[13][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5ce387684404cf922955e4af33ed2367[14]        <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[14][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I84a56b9dce9dfafc97fbdc2ad3b2ae68[14] + 1 :
                                             I84a56b9dce9dfafc97fbdc2ad3b2ae68[14] ;
            I872f61d20baf011e867b44dc5539fc37[14]  <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[14][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5ce387684404cf922955e4af33ed2367[15]        <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[15][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I84a56b9dce9dfafc97fbdc2ad3b2ae68[15] + 1 :
                                             I84a56b9dce9dfafc97fbdc2ad3b2ae68[15] ;
            I872f61d20baf011e867b44dc5539fc37[15]  <=  I84a56b9dce9dfafc97fbdc2ad3b2ae68[15][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1ae87f851f8bd64e6e1428a143e82151[0]        <=  I8afac763670df6f56525d3192e04e784[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8afac763670df6f56525d3192e04e784[0] + 1 :
                                             I8afac763670df6f56525d3192e04e784[0] ;
            Ieb244944e7ee8236a207924f56fbc689[0]  <=  I8afac763670df6f56525d3192e04e784[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1ae87f851f8bd64e6e1428a143e82151[1]        <=  I8afac763670df6f56525d3192e04e784[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8afac763670df6f56525d3192e04e784[1] + 1 :
                                             I8afac763670df6f56525d3192e04e784[1] ;
            Ieb244944e7ee8236a207924f56fbc689[1]  <=  I8afac763670df6f56525d3192e04e784[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1ae87f851f8bd64e6e1428a143e82151[2]        <=  I8afac763670df6f56525d3192e04e784[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8afac763670df6f56525d3192e04e784[2] + 1 :
                                             I8afac763670df6f56525d3192e04e784[2] ;
            Ieb244944e7ee8236a207924f56fbc689[2]  <=  I8afac763670df6f56525d3192e04e784[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1ae87f851f8bd64e6e1428a143e82151[3]        <=  I8afac763670df6f56525d3192e04e784[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8afac763670df6f56525d3192e04e784[3] + 1 :
                                             I8afac763670df6f56525d3192e04e784[3] ;
            Ieb244944e7ee8236a207924f56fbc689[3]  <=  I8afac763670df6f56525d3192e04e784[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1ae87f851f8bd64e6e1428a143e82151[4]        <=  I8afac763670df6f56525d3192e04e784[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8afac763670df6f56525d3192e04e784[4] + 1 :
                                             I8afac763670df6f56525d3192e04e784[4] ;
            Ieb244944e7ee8236a207924f56fbc689[4]  <=  I8afac763670df6f56525d3192e04e784[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1ae87f851f8bd64e6e1428a143e82151[5]        <=  I8afac763670df6f56525d3192e04e784[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8afac763670df6f56525d3192e04e784[5] + 1 :
                                             I8afac763670df6f56525d3192e04e784[5] ;
            Ieb244944e7ee8236a207924f56fbc689[5]  <=  I8afac763670df6f56525d3192e04e784[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1ae87f851f8bd64e6e1428a143e82151[6]        <=  I8afac763670df6f56525d3192e04e784[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8afac763670df6f56525d3192e04e784[6] + 1 :
                                             I8afac763670df6f56525d3192e04e784[6] ;
            Ieb244944e7ee8236a207924f56fbc689[6]  <=  I8afac763670df6f56525d3192e04e784[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1ae87f851f8bd64e6e1428a143e82151[7]        <=  I8afac763670df6f56525d3192e04e784[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8afac763670df6f56525d3192e04e784[7] + 1 :
                                             I8afac763670df6f56525d3192e04e784[7] ;
            Ieb244944e7ee8236a207924f56fbc689[7]  <=  I8afac763670df6f56525d3192e04e784[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1ae87f851f8bd64e6e1428a143e82151[8]        <=  I8afac763670df6f56525d3192e04e784[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8afac763670df6f56525d3192e04e784[8] + 1 :
                                             I8afac763670df6f56525d3192e04e784[8] ;
            Ieb244944e7ee8236a207924f56fbc689[8]  <=  I8afac763670df6f56525d3192e04e784[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I646767a2d4b3029ed7acb73a15af1682[0]        <=  I8cd574c061a4f1bb0da529d2a892324b[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8cd574c061a4f1bb0da529d2a892324b[0] + 1 :
                                             I8cd574c061a4f1bb0da529d2a892324b[0] ;
            Ie9b2be4c32334220e134e041ca8dfc06[0]  <=  I8cd574c061a4f1bb0da529d2a892324b[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I646767a2d4b3029ed7acb73a15af1682[1]        <=  I8cd574c061a4f1bb0da529d2a892324b[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8cd574c061a4f1bb0da529d2a892324b[1] + 1 :
                                             I8cd574c061a4f1bb0da529d2a892324b[1] ;
            Ie9b2be4c32334220e134e041ca8dfc06[1]  <=  I8cd574c061a4f1bb0da529d2a892324b[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I646767a2d4b3029ed7acb73a15af1682[2]        <=  I8cd574c061a4f1bb0da529d2a892324b[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8cd574c061a4f1bb0da529d2a892324b[2] + 1 :
                                             I8cd574c061a4f1bb0da529d2a892324b[2] ;
            Ie9b2be4c32334220e134e041ca8dfc06[2]  <=  I8cd574c061a4f1bb0da529d2a892324b[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I646767a2d4b3029ed7acb73a15af1682[3]        <=  I8cd574c061a4f1bb0da529d2a892324b[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8cd574c061a4f1bb0da529d2a892324b[3] + 1 :
                                             I8cd574c061a4f1bb0da529d2a892324b[3] ;
            Ie9b2be4c32334220e134e041ca8dfc06[3]  <=  I8cd574c061a4f1bb0da529d2a892324b[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I646767a2d4b3029ed7acb73a15af1682[4]        <=  I8cd574c061a4f1bb0da529d2a892324b[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8cd574c061a4f1bb0da529d2a892324b[4] + 1 :
                                             I8cd574c061a4f1bb0da529d2a892324b[4] ;
            Ie9b2be4c32334220e134e041ca8dfc06[4]  <=  I8cd574c061a4f1bb0da529d2a892324b[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I646767a2d4b3029ed7acb73a15af1682[5]        <=  I8cd574c061a4f1bb0da529d2a892324b[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8cd574c061a4f1bb0da529d2a892324b[5] + 1 :
                                             I8cd574c061a4f1bb0da529d2a892324b[5] ;
            Ie9b2be4c32334220e134e041ca8dfc06[5]  <=  I8cd574c061a4f1bb0da529d2a892324b[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I646767a2d4b3029ed7acb73a15af1682[6]        <=  I8cd574c061a4f1bb0da529d2a892324b[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8cd574c061a4f1bb0da529d2a892324b[6] + 1 :
                                             I8cd574c061a4f1bb0da529d2a892324b[6] ;
            Ie9b2be4c32334220e134e041ca8dfc06[6]  <=  I8cd574c061a4f1bb0da529d2a892324b[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I646767a2d4b3029ed7acb73a15af1682[7]        <=  I8cd574c061a4f1bb0da529d2a892324b[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8cd574c061a4f1bb0da529d2a892324b[7] + 1 :
                                             I8cd574c061a4f1bb0da529d2a892324b[7] ;
            Ie9b2be4c32334220e134e041ca8dfc06[7]  <=  I8cd574c061a4f1bb0da529d2a892324b[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I646767a2d4b3029ed7acb73a15af1682[8]        <=  I8cd574c061a4f1bb0da529d2a892324b[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8cd574c061a4f1bb0da529d2a892324b[8] + 1 :
                                             I8cd574c061a4f1bb0da529d2a892324b[8] ;
            Ie9b2be4c32334220e134e041ca8dfc06[8]  <=  I8cd574c061a4f1bb0da529d2a892324b[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I48001f5c6554999a2178308ae271b70e[0]        <=  I919a7f8471a46de33447530b4f3b591d[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I919a7f8471a46de33447530b4f3b591d[0] + 1 :
                                             I919a7f8471a46de33447530b4f3b591d[0] ;
            Id6f07dee3e47f39e3b43329c26f690f7[0]  <=  I919a7f8471a46de33447530b4f3b591d[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I48001f5c6554999a2178308ae271b70e[1]        <=  I919a7f8471a46de33447530b4f3b591d[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I919a7f8471a46de33447530b4f3b591d[1] + 1 :
                                             I919a7f8471a46de33447530b4f3b591d[1] ;
            Id6f07dee3e47f39e3b43329c26f690f7[1]  <=  I919a7f8471a46de33447530b4f3b591d[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I48001f5c6554999a2178308ae271b70e[2]        <=  I919a7f8471a46de33447530b4f3b591d[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I919a7f8471a46de33447530b4f3b591d[2] + 1 :
                                             I919a7f8471a46de33447530b4f3b591d[2] ;
            Id6f07dee3e47f39e3b43329c26f690f7[2]  <=  I919a7f8471a46de33447530b4f3b591d[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I48001f5c6554999a2178308ae271b70e[3]        <=  I919a7f8471a46de33447530b4f3b591d[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I919a7f8471a46de33447530b4f3b591d[3] + 1 :
                                             I919a7f8471a46de33447530b4f3b591d[3] ;
            Id6f07dee3e47f39e3b43329c26f690f7[3]  <=  I919a7f8471a46de33447530b4f3b591d[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I48001f5c6554999a2178308ae271b70e[4]        <=  I919a7f8471a46de33447530b4f3b591d[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I919a7f8471a46de33447530b4f3b591d[4] + 1 :
                                             I919a7f8471a46de33447530b4f3b591d[4] ;
            Id6f07dee3e47f39e3b43329c26f690f7[4]  <=  I919a7f8471a46de33447530b4f3b591d[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I48001f5c6554999a2178308ae271b70e[5]        <=  I919a7f8471a46de33447530b4f3b591d[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I919a7f8471a46de33447530b4f3b591d[5] + 1 :
                                             I919a7f8471a46de33447530b4f3b591d[5] ;
            Id6f07dee3e47f39e3b43329c26f690f7[5]  <=  I919a7f8471a46de33447530b4f3b591d[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I48001f5c6554999a2178308ae271b70e[6]        <=  I919a7f8471a46de33447530b4f3b591d[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I919a7f8471a46de33447530b4f3b591d[6] + 1 :
                                             I919a7f8471a46de33447530b4f3b591d[6] ;
            Id6f07dee3e47f39e3b43329c26f690f7[6]  <=  I919a7f8471a46de33447530b4f3b591d[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I48001f5c6554999a2178308ae271b70e[7]        <=  I919a7f8471a46de33447530b4f3b591d[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I919a7f8471a46de33447530b4f3b591d[7] + 1 :
                                             I919a7f8471a46de33447530b4f3b591d[7] ;
            Id6f07dee3e47f39e3b43329c26f690f7[7]  <=  I919a7f8471a46de33447530b4f3b591d[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I48001f5c6554999a2178308ae271b70e[8]        <=  I919a7f8471a46de33447530b4f3b591d[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I919a7f8471a46de33447530b4f3b591d[8] + 1 :
                                             I919a7f8471a46de33447530b4f3b591d[8] ;
            Id6f07dee3e47f39e3b43329c26f690f7[8]  <=  I919a7f8471a46de33447530b4f3b591d[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7fe6d853fc1c11142b64ff8f40783246[0]        <=  Ib1f53b5c820345ccdba27ab5be3fa49f[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib1f53b5c820345ccdba27ab5be3fa49f[0] + 1 :
                                             Ib1f53b5c820345ccdba27ab5be3fa49f[0] ;
            Ic7f04c065f8ff82c2288f1de77d37189[0]  <=  Ib1f53b5c820345ccdba27ab5be3fa49f[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7fe6d853fc1c11142b64ff8f40783246[1]        <=  Ib1f53b5c820345ccdba27ab5be3fa49f[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib1f53b5c820345ccdba27ab5be3fa49f[1] + 1 :
                                             Ib1f53b5c820345ccdba27ab5be3fa49f[1] ;
            Ic7f04c065f8ff82c2288f1de77d37189[1]  <=  Ib1f53b5c820345ccdba27ab5be3fa49f[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7fe6d853fc1c11142b64ff8f40783246[2]        <=  Ib1f53b5c820345ccdba27ab5be3fa49f[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib1f53b5c820345ccdba27ab5be3fa49f[2] + 1 :
                                             Ib1f53b5c820345ccdba27ab5be3fa49f[2] ;
            Ic7f04c065f8ff82c2288f1de77d37189[2]  <=  Ib1f53b5c820345ccdba27ab5be3fa49f[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7fe6d853fc1c11142b64ff8f40783246[3]        <=  Ib1f53b5c820345ccdba27ab5be3fa49f[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib1f53b5c820345ccdba27ab5be3fa49f[3] + 1 :
                                             Ib1f53b5c820345ccdba27ab5be3fa49f[3] ;
            Ic7f04c065f8ff82c2288f1de77d37189[3]  <=  Ib1f53b5c820345ccdba27ab5be3fa49f[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7fe6d853fc1c11142b64ff8f40783246[4]        <=  Ib1f53b5c820345ccdba27ab5be3fa49f[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib1f53b5c820345ccdba27ab5be3fa49f[4] + 1 :
                                             Ib1f53b5c820345ccdba27ab5be3fa49f[4] ;
            Ic7f04c065f8ff82c2288f1de77d37189[4]  <=  Ib1f53b5c820345ccdba27ab5be3fa49f[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7fe6d853fc1c11142b64ff8f40783246[5]        <=  Ib1f53b5c820345ccdba27ab5be3fa49f[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib1f53b5c820345ccdba27ab5be3fa49f[5] + 1 :
                                             Ib1f53b5c820345ccdba27ab5be3fa49f[5] ;
            Ic7f04c065f8ff82c2288f1de77d37189[5]  <=  Ib1f53b5c820345ccdba27ab5be3fa49f[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7fe6d853fc1c11142b64ff8f40783246[6]        <=  Ib1f53b5c820345ccdba27ab5be3fa49f[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib1f53b5c820345ccdba27ab5be3fa49f[6] + 1 :
                                             Ib1f53b5c820345ccdba27ab5be3fa49f[6] ;
            Ic7f04c065f8ff82c2288f1de77d37189[6]  <=  Ib1f53b5c820345ccdba27ab5be3fa49f[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7fe6d853fc1c11142b64ff8f40783246[7]        <=  Ib1f53b5c820345ccdba27ab5be3fa49f[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib1f53b5c820345ccdba27ab5be3fa49f[7] + 1 :
                                             Ib1f53b5c820345ccdba27ab5be3fa49f[7] ;
            Ic7f04c065f8ff82c2288f1de77d37189[7]  <=  Ib1f53b5c820345ccdba27ab5be3fa49f[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7fe6d853fc1c11142b64ff8f40783246[8]        <=  Ib1f53b5c820345ccdba27ab5be3fa49f[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib1f53b5c820345ccdba27ab5be3fa49f[8] + 1 :
                                             Ib1f53b5c820345ccdba27ab5be3fa49f[8] ;
            Ic7f04c065f8ff82c2288f1de77d37189[8]  <=  Ib1f53b5c820345ccdba27ab5be3fa49f[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iadc98deb917f599574e99a90e3230e88[0]        <=  I384c493c3195d97eea0a9faaec860f78[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I384c493c3195d97eea0a9faaec860f78[0] + 1 :
                                             I384c493c3195d97eea0a9faaec860f78[0] ;
            I4267622319ca65909a3b40484dc74d3a[0]  <=  I384c493c3195d97eea0a9faaec860f78[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iadc98deb917f599574e99a90e3230e88[1]        <=  I384c493c3195d97eea0a9faaec860f78[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I384c493c3195d97eea0a9faaec860f78[1] + 1 :
                                             I384c493c3195d97eea0a9faaec860f78[1] ;
            I4267622319ca65909a3b40484dc74d3a[1]  <=  I384c493c3195d97eea0a9faaec860f78[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iadc98deb917f599574e99a90e3230e88[2]        <=  I384c493c3195d97eea0a9faaec860f78[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I384c493c3195d97eea0a9faaec860f78[2] + 1 :
                                             I384c493c3195d97eea0a9faaec860f78[2] ;
            I4267622319ca65909a3b40484dc74d3a[2]  <=  I384c493c3195d97eea0a9faaec860f78[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iadc98deb917f599574e99a90e3230e88[3]        <=  I384c493c3195d97eea0a9faaec860f78[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I384c493c3195d97eea0a9faaec860f78[3] + 1 :
                                             I384c493c3195d97eea0a9faaec860f78[3] ;
            I4267622319ca65909a3b40484dc74d3a[3]  <=  I384c493c3195d97eea0a9faaec860f78[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iadc98deb917f599574e99a90e3230e88[4]        <=  I384c493c3195d97eea0a9faaec860f78[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I384c493c3195d97eea0a9faaec860f78[4] + 1 :
                                             I384c493c3195d97eea0a9faaec860f78[4] ;
            I4267622319ca65909a3b40484dc74d3a[4]  <=  I384c493c3195d97eea0a9faaec860f78[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iadc98deb917f599574e99a90e3230e88[5]        <=  I384c493c3195d97eea0a9faaec860f78[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I384c493c3195d97eea0a9faaec860f78[5] + 1 :
                                             I384c493c3195d97eea0a9faaec860f78[5] ;
            I4267622319ca65909a3b40484dc74d3a[5]  <=  I384c493c3195d97eea0a9faaec860f78[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iadc98deb917f599574e99a90e3230e88[6]        <=  I384c493c3195d97eea0a9faaec860f78[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I384c493c3195d97eea0a9faaec860f78[6] + 1 :
                                             I384c493c3195d97eea0a9faaec860f78[6] ;
            I4267622319ca65909a3b40484dc74d3a[6]  <=  I384c493c3195d97eea0a9faaec860f78[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iadc98deb917f599574e99a90e3230e88[7]        <=  I384c493c3195d97eea0a9faaec860f78[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I384c493c3195d97eea0a9faaec860f78[7] + 1 :
                                             I384c493c3195d97eea0a9faaec860f78[7] ;
            I4267622319ca65909a3b40484dc74d3a[7]  <=  I384c493c3195d97eea0a9faaec860f78[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iadc98deb917f599574e99a90e3230e88[8]        <=  I384c493c3195d97eea0a9faaec860f78[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I384c493c3195d97eea0a9faaec860f78[8] + 1 :
                                             I384c493c3195d97eea0a9faaec860f78[8] ;
            I4267622319ca65909a3b40484dc74d3a[8]  <=  I384c493c3195d97eea0a9faaec860f78[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iadc98deb917f599574e99a90e3230e88[9]        <=  I384c493c3195d97eea0a9faaec860f78[9][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I384c493c3195d97eea0a9faaec860f78[9] + 1 :
                                             I384c493c3195d97eea0a9faaec860f78[9] ;
            I4267622319ca65909a3b40484dc74d3a[9]  <=  I384c493c3195d97eea0a9faaec860f78[9][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iadc98deb917f599574e99a90e3230e88[10]        <=  I384c493c3195d97eea0a9faaec860f78[10][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I384c493c3195d97eea0a9faaec860f78[10] + 1 :
                                             I384c493c3195d97eea0a9faaec860f78[10] ;
            I4267622319ca65909a3b40484dc74d3a[10]  <=  I384c493c3195d97eea0a9faaec860f78[10][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iadc98deb917f599574e99a90e3230e88[11]        <=  I384c493c3195d97eea0a9faaec860f78[11][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I384c493c3195d97eea0a9faaec860f78[11] + 1 :
                                             I384c493c3195d97eea0a9faaec860f78[11] ;
            I4267622319ca65909a3b40484dc74d3a[11]  <=  I384c493c3195d97eea0a9faaec860f78[11][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3d79461a85cd6a58bf9f96f6e0d704ac[0]        <=  Ida1ee79b7a153e40e91549c2180d8425[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ida1ee79b7a153e40e91549c2180d8425[0] + 1 :
                                             Ida1ee79b7a153e40e91549c2180d8425[0] ;
            Iedd7d4ea8d082b40244c04946dfb14a0[0]  <=  Ida1ee79b7a153e40e91549c2180d8425[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3d79461a85cd6a58bf9f96f6e0d704ac[1]        <=  Ida1ee79b7a153e40e91549c2180d8425[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ida1ee79b7a153e40e91549c2180d8425[1] + 1 :
                                             Ida1ee79b7a153e40e91549c2180d8425[1] ;
            Iedd7d4ea8d082b40244c04946dfb14a0[1]  <=  Ida1ee79b7a153e40e91549c2180d8425[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3d79461a85cd6a58bf9f96f6e0d704ac[2]        <=  Ida1ee79b7a153e40e91549c2180d8425[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ida1ee79b7a153e40e91549c2180d8425[2] + 1 :
                                             Ida1ee79b7a153e40e91549c2180d8425[2] ;
            Iedd7d4ea8d082b40244c04946dfb14a0[2]  <=  Ida1ee79b7a153e40e91549c2180d8425[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3d79461a85cd6a58bf9f96f6e0d704ac[3]        <=  Ida1ee79b7a153e40e91549c2180d8425[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ida1ee79b7a153e40e91549c2180d8425[3] + 1 :
                                             Ida1ee79b7a153e40e91549c2180d8425[3] ;
            Iedd7d4ea8d082b40244c04946dfb14a0[3]  <=  Ida1ee79b7a153e40e91549c2180d8425[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3d79461a85cd6a58bf9f96f6e0d704ac[4]        <=  Ida1ee79b7a153e40e91549c2180d8425[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ida1ee79b7a153e40e91549c2180d8425[4] + 1 :
                                             Ida1ee79b7a153e40e91549c2180d8425[4] ;
            Iedd7d4ea8d082b40244c04946dfb14a0[4]  <=  Ida1ee79b7a153e40e91549c2180d8425[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3d79461a85cd6a58bf9f96f6e0d704ac[5]        <=  Ida1ee79b7a153e40e91549c2180d8425[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ida1ee79b7a153e40e91549c2180d8425[5] + 1 :
                                             Ida1ee79b7a153e40e91549c2180d8425[5] ;
            Iedd7d4ea8d082b40244c04946dfb14a0[5]  <=  Ida1ee79b7a153e40e91549c2180d8425[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3d79461a85cd6a58bf9f96f6e0d704ac[6]        <=  Ida1ee79b7a153e40e91549c2180d8425[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ida1ee79b7a153e40e91549c2180d8425[6] + 1 :
                                             Ida1ee79b7a153e40e91549c2180d8425[6] ;
            Iedd7d4ea8d082b40244c04946dfb14a0[6]  <=  Ida1ee79b7a153e40e91549c2180d8425[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3d79461a85cd6a58bf9f96f6e0d704ac[7]        <=  Ida1ee79b7a153e40e91549c2180d8425[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ida1ee79b7a153e40e91549c2180d8425[7] + 1 :
                                             Ida1ee79b7a153e40e91549c2180d8425[7] ;
            Iedd7d4ea8d082b40244c04946dfb14a0[7]  <=  Ida1ee79b7a153e40e91549c2180d8425[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3d79461a85cd6a58bf9f96f6e0d704ac[8]        <=  Ida1ee79b7a153e40e91549c2180d8425[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ida1ee79b7a153e40e91549c2180d8425[8] + 1 :
                                             Ida1ee79b7a153e40e91549c2180d8425[8] ;
            Iedd7d4ea8d082b40244c04946dfb14a0[8]  <=  Ida1ee79b7a153e40e91549c2180d8425[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3d79461a85cd6a58bf9f96f6e0d704ac[9]        <=  Ida1ee79b7a153e40e91549c2180d8425[9][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ida1ee79b7a153e40e91549c2180d8425[9] + 1 :
                                             Ida1ee79b7a153e40e91549c2180d8425[9] ;
            Iedd7d4ea8d082b40244c04946dfb14a0[9]  <=  Ida1ee79b7a153e40e91549c2180d8425[9][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3d79461a85cd6a58bf9f96f6e0d704ac[10]        <=  Ida1ee79b7a153e40e91549c2180d8425[10][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ida1ee79b7a153e40e91549c2180d8425[10] + 1 :
                                             Ida1ee79b7a153e40e91549c2180d8425[10] ;
            Iedd7d4ea8d082b40244c04946dfb14a0[10]  <=  Ida1ee79b7a153e40e91549c2180d8425[10][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3d79461a85cd6a58bf9f96f6e0d704ac[11]        <=  Ida1ee79b7a153e40e91549c2180d8425[11][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ida1ee79b7a153e40e91549c2180d8425[11] + 1 :
                                             Ida1ee79b7a153e40e91549c2180d8425[11] ;
            Iedd7d4ea8d082b40244c04946dfb14a0[11]  <=  Ida1ee79b7a153e40e91549c2180d8425[11][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2fcbccd884710be9c6a34f78d2ae6a18[0]        <=  Ib6bfc051a54fef77204b41e38cdfc6a8[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib6bfc051a54fef77204b41e38cdfc6a8[0] + 1 :
                                             Ib6bfc051a54fef77204b41e38cdfc6a8[0] ;
            I56e1fe0c7a62589c123876f2b4e57a26[0]  <=  Ib6bfc051a54fef77204b41e38cdfc6a8[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2fcbccd884710be9c6a34f78d2ae6a18[1]        <=  Ib6bfc051a54fef77204b41e38cdfc6a8[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib6bfc051a54fef77204b41e38cdfc6a8[1] + 1 :
                                             Ib6bfc051a54fef77204b41e38cdfc6a8[1] ;
            I56e1fe0c7a62589c123876f2b4e57a26[1]  <=  Ib6bfc051a54fef77204b41e38cdfc6a8[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2fcbccd884710be9c6a34f78d2ae6a18[2]        <=  Ib6bfc051a54fef77204b41e38cdfc6a8[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib6bfc051a54fef77204b41e38cdfc6a8[2] + 1 :
                                             Ib6bfc051a54fef77204b41e38cdfc6a8[2] ;
            I56e1fe0c7a62589c123876f2b4e57a26[2]  <=  Ib6bfc051a54fef77204b41e38cdfc6a8[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2fcbccd884710be9c6a34f78d2ae6a18[3]        <=  Ib6bfc051a54fef77204b41e38cdfc6a8[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib6bfc051a54fef77204b41e38cdfc6a8[3] + 1 :
                                             Ib6bfc051a54fef77204b41e38cdfc6a8[3] ;
            I56e1fe0c7a62589c123876f2b4e57a26[3]  <=  Ib6bfc051a54fef77204b41e38cdfc6a8[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2fcbccd884710be9c6a34f78d2ae6a18[4]        <=  Ib6bfc051a54fef77204b41e38cdfc6a8[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib6bfc051a54fef77204b41e38cdfc6a8[4] + 1 :
                                             Ib6bfc051a54fef77204b41e38cdfc6a8[4] ;
            I56e1fe0c7a62589c123876f2b4e57a26[4]  <=  Ib6bfc051a54fef77204b41e38cdfc6a8[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2fcbccd884710be9c6a34f78d2ae6a18[5]        <=  Ib6bfc051a54fef77204b41e38cdfc6a8[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib6bfc051a54fef77204b41e38cdfc6a8[5] + 1 :
                                             Ib6bfc051a54fef77204b41e38cdfc6a8[5] ;
            I56e1fe0c7a62589c123876f2b4e57a26[5]  <=  Ib6bfc051a54fef77204b41e38cdfc6a8[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2fcbccd884710be9c6a34f78d2ae6a18[6]        <=  Ib6bfc051a54fef77204b41e38cdfc6a8[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib6bfc051a54fef77204b41e38cdfc6a8[6] + 1 :
                                             Ib6bfc051a54fef77204b41e38cdfc6a8[6] ;
            I56e1fe0c7a62589c123876f2b4e57a26[6]  <=  Ib6bfc051a54fef77204b41e38cdfc6a8[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2fcbccd884710be9c6a34f78d2ae6a18[7]        <=  Ib6bfc051a54fef77204b41e38cdfc6a8[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib6bfc051a54fef77204b41e38cdfc6a8[7] + 1 :
                                             Ib6bfc051a54fef77204b41e38cdfc6a8[7] ;
            I56e1fe0c7a62589c123876f2b4e57a26[7]  <=  Ib6bfc051a54fef77204b41e38cdfc6a8[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2fcbccd884710be9c6a34f78d2ae6a18[8]        <=  Ib6bfc051a54fef77204b41e38cdfc6a8[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib6bfc051a54fef77204b41e38cdfc6a8[8] + 1 :
                                             Ib6bfc051a54fef77204b41e38cdfc6a8[8] ;
            I56e1fe0c7a62589c123876f2b4e57a26[8]  <=  Ib6bfc051a54fef77204b41e38cdfc6a8[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2fcbccd884710be9c6a34f78d2ae6a18[9]        <=  Ib6bfc051a54fef77204b41e38cdfc6a8[9][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib6bfc051a54fef77204b41e38cdfc6a8[9] + 1 :
                                             Ib6bfc051a54fef77204b41e38cdfc6a8[9] ;
            I56e1fe0c7a62589c123876f2b4e57a26[9]  <=  Ib6bfc051a54fef77204b41e38cdfc6a8[9][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2fcbccd884710be9c6a34f78d2ae6a18[10]        <=  Ib6bfc051a54fef77204b41e38cdfc6a8[10][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib6bfc051a54fef77204b41e38cdfc6a8[10] + 1 :
                                             Ib6bfc051a54fef77204b41e38cdfc6a8[10] ;
            I56e1fe0c7a62589c123876f2b4e57a26[10]  <=  Ib6bfc051a54fef77204b41e38cdfc6a8[10][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2fcbccd884710be9c6a34f78d2ae6a18[11]        <=  Ib6bfc051a54fef77204b41e38cdfc6a8[11][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib6bfc051a54fef77204b41e38cdfc6a8[11] + 1 :
                                             Ib6bfc051a54fef77204b41e38cdfc6a8[11] ;
            I56e1fe0c7a62589c123876f2b4e57a26[11]  <=  Ib6bfc051a54fef77204b41e38cdfc6a8[11][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3d3df5d4d89adf508497bac8d75ef0c6[0]        <=  Ie6d740bc0451311c5f93f4954812613d[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie6d740bc0451311c5f93f4954812613d[0] + 1 :
                                             Ie6d740bc0451311c5f93f4954812613d[0] ;
            Ia8a468877c9f96713c8141df9205f92a[0]  <=  Ie6d740bc0451311c5f93f4954812613d[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3d3df5d4d89adf508497bac8d75ef0c6[1]        <=  Ie6d740bc0451311c5f93f4954812613d[1][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie6d740bc0451311c5f93f4954812613d[1] + 1 :
                                             Ie6d740bc0451311c5f93f4954812613d[1] ;
            Ia8a468877c9f96713c8141df9205f92a[1]  <=  Ie6d740bc0451311c5f93f4954812613d[1][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3d3df5d4d89adf508497bac8d75ef0c6[2]        <=  Ie6d740bc0451311c5f93f4954812613d[2][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie6d740bc0451311c5f93f4954812613d[2] + 1 :
                                             Ie6d740bc0451311c5f93f4954812613d[2] ;
            Ia8a468877c9f96713c8141df9205f92a[2]  <=  Ie6d740bc0451311c5f93f4954812613d[2][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3d3df5d4d89adf508497bac8d75ef0c6[3]        <=  Ie6d740bc0451311c5f93f4954812613d[3][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie6d740bc0451311c5f93f4954812613d[3] + 1 :
                                             Ie6d740bc0451311c5f93f4954812613d[3] ;
            Ia8a468877c9f96713c8141df9205f92a[3]  <=  Ie6d740bc0451311c5f93f4954812613d[3][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3d3df5d4d89adf508497bac8d75ef0c6[4]        <=  Ie6d740bc0451311c5f93f4954812613d[4][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie6d740bc0451311c5f93f4954812613d[4] + 1 :
                                             Ie6d740bc0451311c5f93f4954812613d[4] ;
            Ia8a468877c9f96713c8141df9205f92a[4]  <=  Ie6d740bc0451311c5f93f4954812613d[4][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3d3df5d4d89adf508497bac8d75ef0c6[5]        <=  Ie6d740bc0451311c5f93f4954812613d[5][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie6d740bc0451311c5f93f4954812613d[5] + 1 :
                                             Ie6d740bc0451311c5f93f4954812613d[5] ;
            Ia8a468877c9f96713c8141df9205f92a[5]  <=  Ie6d740bc0451311c5f93f4954812613d[5][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3d3df5d4d89adf508497bac8d75ef0c6[6]        <=  Ie6d740bc0451311c5f93f4954812613d[6][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie6d740bc0451311c5f93f4954812613d[6] + 1 :
                                             Ie6d740bc0451311c5f93f4954812613d[6] ;
            Ia8a468877c9f96713c8141df9205f92a[6]  <=  Ie6d740bc0451311c5f93f4954812613d[6][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3d3df5d4d89adf508497bac8d75ef0c6[7]        <=  Ie6d740bc0451311c5f93f4954812613d[7][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie6d740bc0451311c5f93f4954812613d[7] + 1 :
                                             Ie6d740bc0451311c5f93f4954812613d[7] ;
            Ia8a468877c9f96713c8141df9205f92a[7]  <=  Ie6d740bc0451311c5f93f4954812613d[7][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3d3df5d4d89adf508497bac8d75ef0c6[8]        <=  Ie6d740bc0451311c5f93f4954812613d[8][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie6d740bc0451311c5f93f4954812613d[8] + 1 :
                                             Ie6d740bc0451311c5f93f4954812613d[8] ;
            Ia8a468877c9f96713c8141df9205f92a[8]  <=  Ie6d740bc0451311c5f93f4954812613d[8][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3d3df5d4d89adf508497bac8d75ef0c6[9]        <=  Ie6d740bc0451311c5f93f4954812613d[9][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie6d740bc0451311c5f93f4954812613d[9] + 1 :
                                             Ie6d740bc0451311c5f93f4954812613d[9] ;
            Ia8a468877c9f96713c8141df9205f92a[9]  <=  Ie6d740bc0451311c5f93f4954812613d[9][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3d3df5d4d89adf508497bac8d75ef0c6[10]        <=  Ie6d740bc0451311c5f93f4954812613d[10][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie6d740bc0451311c5f93f4954812613d[10] + 1 :
                                             Ie6d740bc0451311c5f93f4954812613d[10] ;
            Ia8a468877c9f96713c8141df9205f92a[10]  <=  Ie6d740bc0451311c5f93f4954812613d[10][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3d3df5d4d89adf508497bac8d75ef0c6[11]        <=  Ie6d740bc0451311c5f93f4954812613d[11][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie6d740bc0451311c5f93f4954812613d[11] + 1 :
                                             Ie6d740bc0451311c5f93f4954812613d[11] ;
            Ia8a468877c9f96713c8141df9205f92a[11]  <=  Ie6d740bc0451311c5f93f4954812613d[11][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iadecdac113e45cd08e095317d07766e5[0]        <=  Ia6ac09257dfd071a132e96619a662f57[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia6ac09257dfd071a132e96619a662f57[0] + 1 :
                                             Ia6ac09257dfd071a132e96619a662f57[0] ;
            Ida6059c6e0890f730536f97dfb83770b[0]  <=  Ia6ac09257dfd071a132e96619a662f57[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2e4a339cb29f80caa8cbd630a0372ae8[0]        <=  Id2e5704c73c707a217875dbf2743e6f3[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Id2e5704c73c707a217875dbf2743e6f3[0] + 1 :
                                             Id2e5704c73c707a217875dbf2743e6f3[0] ;
            I1993c1ed200d7cdf838d23c72a0c1c0b[0]  <=  Id2e5704c73c707a217875dbf2743e6f3[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I423e8e9a9f19cf712372622e5c80c732[0]        <=  If152a76f9c612e979151b8f51262efc1[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~If152a76f9c612e979151b8f51262efc1[0] + 1 :
                                             If152a76f9c612e979151b8f51262efc1[0] ;
            I07e04e352df9aa1988ccf05d9cb2d1d7[0]  <=  If152a76f9c612e979151b8f51262efc1[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5434db7480d96327d98156af57961745[0]        <=  Ifdb6febe29caf3ce300d9cea4954927a[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ifdb6febe29caf3ce300d9cea4954927a[0] + 1 :
                                             Ifdb6febe29caf3ce300d9cea4954927a[0] ;
            Ic4c0ebcc3711c9844a3aa3875483d2f7[0]  <=  Ifdb6febe29caf3ce300d9cea4954927a[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I20ebcbecf2c13a53be05ff26552b4e72[0]        <=  Icfb2b3a2e096f55ba29dd2f9b5761852[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Icfb2b3a2e096f55ba29dd2f9b5761852[0] + 1 :
                                             Icfb2b3a2e096f55ba29dd2f9b5761852[0] ;
            I28e344560ba76bb3b76d01d8c53693a9[0]  <=  Icfb2b3a2e096f55ba29dd2f9b5761852[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7ba72e4bac9bd64d046733ce50f43769[0]        <=  I06c6597547e69bb46e1bede7b7b7f24a[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I06c6597547e69bb46e1bede7b7b7f24a[0] + 1 :
                                             I06c6597547e69bb46e1bede7b7b7f24a[0] ;
            I0600def6e6caada88ba6dedbb0d322ac[0]  <=  I06c6597547e69bb46e1bede7b7b7f24a[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6614526a756edaabd6a25e858b472d14[0]        <=  I325f629c52919e62b3c0075481267744[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I325f629c52919e62b3c0075481267744[0] + 1 :
                                             I325f629c52919e62b3c0075481267744[0] ;
            Iddbf50612c89b5b95a5c9efb5575cae3[0]  <=  I325f629c52919e62b3c0075481267744[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I47b2e8ee0c69e5301365a25d512b1ece[0]        <=  I56dc657b33a933d2e5d3ac517a9d1fef[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I56dc657b33a933d2e5d3ac517a9d1fef[0] + 1 :
                                             I56dc657b33a933d2e5d3ac517a9d1fef[0] ;
            Iadc8f7f87b50bfff53d2d12d82489829[0]  <=  I56dc657b33a933d2e5d3ac517a9d1fef[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ibb72eb38996b41ce253875df0f620eb7[0]        <=  Ie17d5d171cb71e3748dd0b6c800263ca[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie17d5d171cb71e3748dd0b6c800263ca[0] + 1 :
                                             Ie17d5d171cb71e3748dd0b6c800263ca[0] ;
            I53a658b443200b9f11f1830547b5f42d[0]  <=  Ie17d5d171cb71e3748dd0b6c800263ca[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I66944cd8c5bc22cd92a5cfcd68cee426[0]        <=  I9cabb772f5988b877afae0c3b65f340a[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I9cabb772f5988b877afae0c3b65f340a[0] + 1 :
                                             I9cabb772f5988b877afae0c3b65f340a[0] ;
            I170f424df45651abe215ec74d649a9eb[0]  <=  I9cabb772f5988b877afae0c3b65f340a[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8f2ff78b78e43fe7f6780f19d92ff7b8[0]        <=  Ie29294b754845c1c5602dade95c9e762[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie29294b754845c1c5602dade95c9e762[0] + 1 :
                                             Ie29294b754845c1c5602dade95c9e762[0] ;
            I3c897bfed190017a876c44fd73a7ecea[0]  <=  Ie29294b754845c1c5602dade95c9e762[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ieea0e49da41cdf0d062217a6e6591728[0]        <=  Ibfc5db8e8f393324f06568278da33b4e[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ibfc5db8e8f393324f06568278da33b4e[0] + 1 :
                                             Ibfc5db8e8f393324f06568278da33b4e[0] ;
            Iaecbbae967be2c62cacf2fa7f9801899[0]  <=  Ibfc5db8e8f393324f06568278da33b4e[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I699c35d4b3c36c35ecaadb87c8b35d9a[0]        <=  I44aace203d154a4d0fc8f10f2cdc5626[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I44aace203d154a4d0fc8f10f2cdc5626[0] + 1 :
                                             I44aace203d154a4d0fc8f10f2cdc5626[0] ;
            I52f867f1009f2e8d18b50a777942bde3[0]  <=  I44aace203d154a4d0fc8f10f2cdc5626[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie6c95c6ddde379ca7437e78c42a8245e[0]        <=  I75526eea62d190615e13ac2731e07074[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I75526eea62d190615e13ac2731e07074[0] + 1 :
                                             I75526eea62d190615e13ac2731e07074[0] ;
            I56a39a0c67b1de0a3cab6c61af3eebcf[0]  <=  I75526eea62d190615e13ac2731e07074[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I85e05de515eb28d7172a95ba55da82a2[0]        <=  I67bc090d5c81788569b837217febf22d[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I67bc090d5c81788569b837217febf22d[0] + 1 :
                                             I67bc090d5c81788569b837217febf22d[0] ;
            I490a65b3f7b30540906262ec5e12717b[0]  <=  I67bc090d5c81788569b837217febf22d[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7ed14b994ecbeae0536a721e16c88489[0]        <=  I28d725840d5db12ad4940ef965775cc4[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I28d725840d5db12ad4940ef965775cc4[0] + 1 :
                                             I28d725840d5db12ad4940ef965775cc4[0] ;
            Ib3c52fef8251d95e9abc8df0aad45d4e[0]  <=  I28d725840d5db12ad4940ef965775cc4[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iad29b892bf50a3e83e4eb9b7c271292a[0]        <=  Ia9e617fb96d7ae3706736fafa5dce67c[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia9e617fb96d7ae3706736fafa5dce67c[0] + 1 :
                                             Ia9e617fb96d7ae3706736fafa5dce67c[0] ;
            If75725e534dcb00364d73a42769539fb[0]  <=  Ia9e617fb96d7ae3706736fafa5dce67c[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I35d2bc3f0efd23ded421f195b62a6a33[0]        <=  Ie033e6fdf59cdfd67ff238b68924dfb5[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie033e6fdf59cdfd67ff238b68924dfb5[0] + 1 :
                                             Ie033e6fdf59cdfd67ff238b68924dfb5[0] ;
            I9ddc427eef437ecc3ac4a2cf52aad4c3[0]  <=  Ie033e6fdf59cdfd67ff238b68924dfb5[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I4aaa94237ac5b28ce1d0db0d4e15ff81[0]        <=  I6190c7e2fd99fcb3394fc330e0b08678[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I6190c7e2fd99fcb3394fc330e0b08678[0] + 1 :
                                             I6190c7e2fd99fcb3394fc330e0b08678[0] ;
            I8999ca1f2fe9d4a30bd38fcb0daad2a4[0]  <=  I6190c7e2fd99fcb3394fc330e0b08678[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I137145b608dfe5138d4bdbea237743bd[0]        <=  I91f50b160f3a0bc73c84123d977fa4ab[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I91f50b160f3a0bc73c84123d977fa4ab[0] + 1 :
                                             I91f50b160f3a0bc73c84123d977fa4ab[0] ;
            Ie11cf6677812bb739255b053a9c9cd56[0]  <=  I91f50b160f3a0bc73c84123d977fa4ab[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I68a784efb51b172af79e3dec88d529e1[0]        <=  Ic05ea9ae53b9396b54c4484a56c7ec79[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic05ea9ae53b9396b54c4484a56c7ec79[0] + 1 :
                                             Ic05ea9ae53b9396b54c4484a56c7ec79[0] ;
            Iacc1d5a5c7811f0c9326ef80d1154fbb[0]  <=  Ic05ea9ae53b9396b54c4484a56c7ec79[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic3036adab4495c6a59055dd34a28b2e5[0]        <=  Icf4d6deb47e202e607a07639d064ca55[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Icf4d6deb47e202e607a07639d064ca55[0] + 1 :
                                             Icf4d6deb47e202e607a07639d064ca55[0] ;
            I0efdadfd49c035a49d92243391395bca[0]  <=  Icf4d6deb47e202e607a07639d064ca55[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I84a699063d2a7944f4a1b72b67ab5b4f[0]        <=  I85ee05cc8e67b77acbd3ddc7fdfd6bca[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I85ee05cc8e67b77acbd3ddc7fdfd6bca[0] + 1 :
                                             I85ee05cc8e67b77acbd3ddc7fdfd6bca[0] ;
            Ie34d59bc77e06807937fe6f6860527e9[0]  <=  I85ee05cc8e67b77acbd3ddc7fdfd6bca[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I63acf3ed504ad084a12a219790842b4a[0]        <=  I803822a38e626e789a50bade0961edab[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I803822a38e626e789a50bade0961edab[0] + 1 :
                                             I803822a38e626e789a50bade0961edab[0] ;
            I9661cb126908d8550b585e2bad383bd6[0]  <=  I803822a38e626e789a50bade0961edab[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I23a2a7fb24650eec8812d8671d92bf2b[0]        <=  If93330fbf9bc863d2837ffc2a0466e70[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~If93330fbf9bc863d2837ffc2a0466e70[0] + 1 :
                                             If93330fbf9bc863d2837ffc2a0466e70[0] ;
            Ic0b832fbcbdb57745fefcc1ac1438808[0]  <=  If93330fbf9bc863d2837ffc2a0466e70[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6f9156b7b5e13529ec0c34da34cb2b04[0]        <=  I8ac880ea1c849c493c66a82534400d8c[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8ac880ea1c849c493c66a82534400d8c[0] + 1 :
                                             I8ac880ea1c849c493c66a82534400d8c[0] ;
            I2afd96714b26f30483c3935c2a68e64f[0]  <=  I8ac880ea1c849c493c66a82534400d8c[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I09a4c92baceef72d764c6880fb62c1f7[0]        <=  I7cf96d4e28b02fd623d8c76161410eb6[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I7cf96d4e28b02fd623d8c76161410eb6[0] + 1 :
                                             I7cf96d4e28b02fd623d8c76161410eb6[0] ;
            Id6d4165b752630a1ce7ceb77fdcee477[0]  <=  I7cf96d4e28b02fd623d8c76161410eb6[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I13a44a5dfbb198be64c99845122a6e97[0]        <=  I637636f1d78f96c75bf5c3841419e9fe[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I637636f1d78f96c75bf5c3841419e9fe[0] + 1 :
                                             I637636f1d78f96c75bf5c3841419e9fe[0] ;
            I59baaf1ad22721cde9064b8aad65ac76[0]  <=  I637636f1d78f96c75bf5c3841419e9fe[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2b57472e34677b9aafb852a3e421270d[0]        <=  Icc7d8812ba512a84d2905f1182e69d0a[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Icc7d8812ba512a84d2905f1182e69d0a[0] + 1 :
                                             Icc7d8812ba512a84d2905f1182e69d0a[0] ;
            I9094f4e9c5b60add3acee212118a1dfa[0]  <=  Icc7d8812ba512a84d2905f1182e69d0a[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic96e056f2208c211122e5008d5fd8ced[0]        <=  Iba60ce25380dc39b44ba505a04453614[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Iba60ce25380dc39b44ba505a04453614[0] + 1 :
                                             Iba60ce25380dc39b44ba505a04453614[0] ;
            I13168bab2231ed22a3509142f990e408[0]  <=  Iba60ce25380dc39b44ba505a04453614[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie6b1ee6dfca427a82e4d1016585682d9[0]        <=  I9a6a2b184e5122aaa964c2bc818c255d[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I9a6a2b184e5122aaa964c2bc818c255d[0] + 1 :
                                             I9a6a2b184e5122aaa964c2bc818c255d[0] ;
            I280145f996e5e249788cacca7caf0095[0]  <=  I9a6a2b184e5122aaa964c2bc818c255d[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ieb0276790e2d912809acc7f3a409ac37[0]        <=  I4dea7825b6a0eab3aebeb7c4889cdae9[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I4dea7825b6a0eab3aebeb7c4889cdae9[0] + 1 :
                                             I4dea7825b6a0eab3aebeb7c4889cdae9[0] ;
            Ia9db6d176e9b9579a1aa5f257cd1a9f6[0]  <=  I4dea7825b6a0eab3aebeb7c4889cdae9[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9883bdcc250c2eb1f8e691d0f18b3cbc[0]        <=  I4809ebf07d855a2e48f92df77ac08b89[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I4809ebf07d855a2e48f92df77ac08b89[0] + 1 :
                                             I4809ebf07d855a2e48f92df77ac08b89[0] ;
            I0ed43cf9eec83545457c57cfb6181d3c[0]  <=  I4809ebf07d855a2e48f92df77ac08b89[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I28f58fec52ea2df3fa3d8e4a2722468b[0]        <=  Ie0a958d83a20d204b3e7a9b4235c4b19[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie0a958d83a20d204b3e7a9b4235c4b19[0] + 1 :
                                             Ie0a958d83a20d204b3e7a9b4235c4b19[0] ;
            I5b74f5fc705a0406ff2376cb8ac11db4[0]  <=  Ie0a958d83a20d204b3e7a9b4235c4b19[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ibf1bb88a30c8519cf22f684a9bc552e9[0]        <=  I8280db7b6ab8c525afd18dc79c0715fb[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8280db7b6ab8c525afd18dc79c0715fb[0] + 1 :
                                             I8280db7b6ab8c525afd18dc79c0715fb[0] ;
            I14f0d3ad4fec9ca492d6b36eb29a5dea[0]  <=  I8280db7b6ab8c525afd18dc79c0715fb[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9d2131bc965972708385d8d79c5b1687[0]        <=  Ifd4e06675d2b57e0064369490c20b8ba[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ifd4e06675d2b57e0064369490c20b8ba[0] + 1 :
                                             Ifd4e06675d2b57e0064369490c20b8ba[0] ;
            I3a25c80d9bf7655f4ce70cf29843db43[0]  <=  Ifd4e06675d2b57e0064369490c20b8ba[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I65dc268c49445ceeef922f9c273df755[0]        <=  I887915cd3be831277d41e47417ae42e7[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I887915cd3be831277d41e47417ae42e7[0] + 1 :
                                             I887915cd3be831277d41e47417ae42e7[0] ;
            I260dc9154b3a9fe38b0948e807bdb42d[0]  <=  I887915cd3be831277d41e47417ae42e7[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7c0af5fba885dca550df150029e9ee36[0]        <=  Ic3af54bfe225c905cd146c6ccd3e34e6[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic3af54bfe225c905cd146c6ccd3e34e6[0] + 1 :
                                             Ic3af54bfe225c905cd146c6ccd3e34e6[0] ;
            Ic49b2c150e2face8c362e33f2d87f9c4[0]  <=  Ic3af54bfe225c905cd146c6ccd3e34e6[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If26299fbf3d11a469aa2bc573760fed0[0]        <=  Ida4ab0033193d0b40f4ab5d8b74d7625[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ida4ab0033193d0b40f4ab5d8b74d7625[0] + 1 :
                                             Ida4ab0033193d0b40f4ab5d8b74d7625[0] ;
            I714350b3b56a3249aad06d5f59fbb291[0]  <=  Ida4ab0033193d0b40f4ab5d8b74d7625[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2ba80daf0c2b625370644ab47cef63e9[0]        <=  Ic0c2d77062c77982f91941bd99eea68a[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic0c2d77062c77982f91941bd99eea68a[0] + 1 :
                                             Ic0c2d77062c77982f91941bd99eea68a[0] ;
            Ia318eb500b8bd71048bde375c1db65a6[0]  <=  Ic0c2d77062c77982f91941bd99eea68a[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0911e01c831a9e46568122fa6dab2357[0]        <=  I783f9d09de5fce4d69c179fb398a58ae[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I783f9d09de5fce4d69c179fb398a58ae[0] + 1 :
                                             I783f9d09de5fce4d69c179fb398a58ae[0] ;
            Ia2c4192b1e4f180402550aebcf1dcd1f[0]  <=  I783f9d09de5fce4d69c179fb398a58ae[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic8f0aa27dadc689b1bfb5b284fc13562[0]        <=  I0af2bc8f858473a4b6f9467d5635f2ed[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I0af2bc8f858473a4b6f9467d5635f2ed[0] + 1 :
                                             I0af2bc8f858473a4b6f9467d5635f2ed[0] ;
            I1686a95674ecad0c4e234b8aa6e22dd9[0]  <=  I0af2bc8f858473a4b6f9467d5635f2ed[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5ad4c6aba210a8b2d343ab17b49c38a3[0]        <=  Id882b47b85085b9603449499ecfcdb49[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Id882b47b85085b9603449499ecfcdb49[0] + 1 :
                                             Id882b47b85085b9603449499ecfcdb49[0] ;
            I5ee21680396395f8338477fa2bb314ec[0]  <=  Id882b47b85085b9603449499ecfcdb49[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I34947a54412d287f3ff730332211dc5a[0]        <=  I5b2752f489336c41887046ed4673a717[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I5b2752f489336c41887046ed4673a717[0] + 1 :
                                             I5b2752f489336c41887046ed4673a717[0] ;
            I005e89f0a9a9a52aec92752813a70f81[0]  <=  I5b2752f489336c41887046ed4673a717[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ia6ac380b9be591fb53c0f36f4d417a7e[0]        <=  I75b2328b94afd38404e28c46d7358b22[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I75b2328b94afd38404e28c46d7358b22[0] + 1 :
                                             I75b2328b94afd38404e28c46d7358b22[0] ;
            I0daca3ad02a67285295cd9fc330d8027[0]  <=  I75b2328b94afd38404e28c46d7358b22[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ia5d5342af30d46f66f0e4f41e5170b87[0]        <=  I7a642ae71b9f5454a31702d6c3197c79[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I7a642ae71b9f5454a31702d6c3197c79[0] + 1 :
                                             I7a642ae71b9f5454a31702d6c3197c79[0] ;
            I0d2ddde9edfef483482e6c177a084f6e[0]  <=  I7a642ae71b9f5454a31702d6c3197c79[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ica011579f46e949eda7f8eed2e4d3ada[0]        <=  I0f8357de84a9c9e19d35ddd0715b7be4[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I0f8357de84a9c9e19d35ddd0715b7be4[0] + 1 :
                                             I0f8357de84a9c9e19d35ddd0715b7be4[0] ;
            I932ad562b582e2c9795f241c82901188[0]  <=  I0f8357de84a9c9e19d35ddd0715b7be4[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I88b214aeebaffa768ccf7c70423fb0c3[0]        <=  I76599476765ec5b54c1ed75efddc909d[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I76599476765ec5b54c1ed75efddc909d[0] + 1 :
                                             I76599476765ec5b54c1ed75efddc909d[0] ;
            Ifee4aa12e36833c935c54ef27b1917da[0]  <=  I76599476765ec5b54c1ed75efddc909d[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If46340645f788fdde3bb8f4d176aae52[0]        <=  I9e277097d3f55ad75b5b0e819d6d3651[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I9e277097d3f55ad75b5b0e819d6d3651[0] + 1 :
                                             I9e277097d3f55ad75b5b0e819d6d3651[0] ;
            I51e5b79f738795719ac21c6a88711a01[0]  <=  I9e277097d3f55ad75b5b0e819d6d3651[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib59f285283d8c3013c20aad73ed9d148[0]        <=  Ibade670ce04ec07f3b5174fcfc67fabb[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ibade670ce04ec07f3b5174fcfc67fabb[0] + 1 :
                                             Ibade670ce04ec07f3b5174fcfc67fabb[0] ;
            I4e41e628a8af629421544cb4c6f45265[0]  <=  Ibade670ce04ec07f3b5174fcfc67fabb[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3229ea9a0c348b17fcaedf6565d6d7cc[0]        <=  I19a9636de4b8153208ebef0cfbf811ea[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I19a9636de4b8153208ebef0cfbf811ea[0] + 1 :
                                             I19a9636de4b8153208ebef0cfbf811ea[0] ;
            I9b2ec7db66661f7c9d85cfb1bc41893b[0]  <=  I19a9636de4b8153208ebef0cfbf811ea[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3ba17818aa7ea9bbfcebb2a5f405fec1[0]        <=  Ieb302f84fbd92b0fa4a5747cb1764926[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ieb302f84fbd92b0fa4a5747cb1764926[0] + 1 :
                                             Ieb302f84fbd92b0fa4a5747cb1764926[0] ;
            I0a594a36728c7ac6244c504b8ea9c9af[0]  <=  Ieb302f84fbd92b0fa4a5747cb1764926[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2ad1769ceb4cf0013f7b032c6e583745[0]        <=  If88f7bba0fc9ca004e41cf047f6e6410[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~If88f7bba0fc9ca004e41cf047f6e6410[0] + 1 :
                                             If88f7bba0fc9ca004e41cf047f6e6410[0] ;
            Ibd943ebf64fe56a1818d2bb8b9f9f8bd[0]  <=  If88f7bba0fc9ca004e41cf047f6e6410[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib35d4bfa08a9364f7f6c8be7feaf15ba[0]        <=  I5989aa844d0d73de1a11b8902002efee[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I5989aa844d0d73de1a11b8902002efee[0] + 1 :
                                             I5989aa844d0d73de1a11b8902002efee[0] ;
            I8c3ba90c84f9375001e727b711dead8d[0]  <=  I5989aa844d0d73de1a11b8902002efee[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I216edc2024d31f612d05617f6696c6c5[0]        <=  Ia683e321a3334e9668b39f5fea591cd4[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ia683e321a3334e9668b39f5fea591cd4[0] + 1 :
                                             Ia683e321a3334e9668b39f5fea591cd4[0] ;
            I387ca23d0e2183522ab041ec48bffef4[0]  <=  Ia683e321a3334e9668b39f5fea591cd4[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2be51c29373fe2ddfe456265a54bcc08[0]        <=  Ic16cfcc11cd03b06afab4b96ab13a350[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic16cfcc11cd03b06afab4b96ab13a350[0] + 1 :
                                             Ic16cfcc11cd03b06afab4b96ab13a350[0] ;
            Ib933575f5224d414f87bc71fa7498534[0]  <=  Ic16cfcc11cd03b06afab4b96ab13a350[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib3561cb8090e7787ad8c324db3a5456a[0]        <=  Icb19ea7dbeb8d826bf85e1e8518e7558[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Icb19ea7dbeb8d826bf85e1e8518e7558[0] + 1 :
                                             Icb19ea7dbeb8d826bf85e1e8518e7558[0] ;
            Ibfe1bddf32fa63ea87c68de7a3af1815[0]  <=  Icb19ea7dbeb8d826bf85e1e8518e7558[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5d701e34c6fea83dccbac286a36fcbbc[0]        <=  Ie1c0888b2c811ca399501f4669dd8267[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie1c0888b2c811ca399501f4669dd8267[0] + 1 :
                                             Ie1c0888b2c811ca399501f4669dd8267[0] ;
            I719c50f9bbc66decebe794fe6ea017dd[0]  <=  Ie1c0888b2c811ca399501f4669dd8267[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie479179aee4de4208dda8af63ed9fb66[0]        <=  I65008ba6af7af0ee93fd085692ff4705[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I65008ba6af7af0ee93fd085692ff4705[0] + 1 :
                                             I65008ba6af7af0ee93fd085692ff4705[0] ;
            I833b0433a33dac70cb215bc8cc9f4863[0]  <=  I65008ba6af7af0ee93fd085692ff4705[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0acbd9a7ed1409c7958d6c630a7f96d7[0]        <=  I0818a864ca9a381fd4b8492410037437[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I0818a864ca9a381fd4b8492410037437[0] + 1 :
                                             I0818a864ca9a381fd4b8492410037437[0] ;
            I9769761eb863e3273f9253ace4c69585[0]  <=  I0818a864ca9a381fd4b8492410037437[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I390dbe9907497b62162445c90f2f27fc[0]        <=  I11e799346dda7e851c5d48f116216d5a[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I11e799346dda7e851c5d48f116216d5a[0] + 1 :
                                             I11e799346dda7e851c5d48f116216d5a[0] ;
            I1fc63f388d047207a9375842c85e87f7[0]  <=  I11e799346dda7e851c5d48f116216d5a[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I01d386885d97d770ff2ab01da72631a0[0]        <=  I1bea6ddcb374caef97e35af1eb33d878[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I1bea6ddcb374caef97e35af1eb33d878[0] + 1 :
                                             I1bea6ddcb374caef97e35af1eb33d878[0] ;
            I414c4d389ecc00197f2138eff0b6454e[0]  <=  I1bea6ddcb374caef97e35af1eb33d878[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iedbfdad739e796202d764f909e6ac6b2[0]        <=  Iae87b81938ba6be7fcfb902e35b55ff2[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Iae87b81938ba6be7fcfb902e35b55ff2[0] + 1 :
                                             Iae87b81938ba6be7fcfb902e35b55ff2[0] ;
            Ibe387e8fe6f35588e028ba29cda5b912[0]  <=  Iae87b81938ba6be7fcfb902e35b55ff2[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I41ded014d071bd714d053a8aed21cf5a[0]        <=  I2cf76e56c5212c0921ac6725ca41be3c[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I2cf76e56c5212c0921ac6725ca41be3c[0] + 1 :
                                             I2cf76e56c5212c0921ac6725ca41be3c[0] ;
            I98191a7e6c56aae1b56e3d623004ed75[0]  <=  I2cf76e56c5212c0921ac6725ca41be3c[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1f14df209c8c73fe390873ae05063afe[0]        <=  I21cf97f59f8387bdd451934e800a501d[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I21cf97f59f8387bdd451934e800a501d[0] + 1 :
                                             I21cf97f59f8387bdd451934e800a501d[0] ;
            Icd0f5c370462670cd18d30dfc0c81c02[0]  <=  I21cf97f59f8387bdd451934e800a501d[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I510a362375a9b9c75436ad01388de6db[0]        <=  I9c91a8ca3a41b5df249ad6e0cd9b6601[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I9c91a8ca3a41b5df249ad6e0cd9b6601[0] + 1 :
                                             I9c91a8ca3a41b5df249ad6e0cd9b6601[0] ;
            I15c59dc8eba10ff8eadfa6078678773b[0]  <=  I9c91a8ca3a41b5df249ad6e0cd9b6601[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic2f0b44a83961b8b49f4637ec6750f27[0]        <=  I02e4ad55fc6e12cd60370ae782bbd36b[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I02e4ad55fc6e12cd60370ae782bbd36b[0] + 1 :
                                             I02e4ad55fc6e12cd60370ae782bbd36b[0] ;
            I3870d672343c002ad9c83c816fd40567[0]  <=  I02e4ad55fc6e12cd60370ae782bbd36b[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id5cbccb1a2ccacf28b64ece8eec0099e[0]        <=  I5192b23d7d4742e17ffcf58679d96734[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I5192b23d7d4742e17ffcf58679d96734[0] + 1 :
                                             I5192b23d7d4742e17ffcf58679d96734[0] ;
            Ic341b9d947f2d3ac57aa41f408214434[0]  <=  I5192b23d7d4742e17ffcf58679d96734[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9686b2d0e5248bfb6d3ef9b7c687ed05[0]        <=  I0aaea02d5fbc4cfe6478060df6a92441[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I0aaea02d5fbc4cfe6478060df6a92441[0] + 1 :
                                             I0aaea02d5fbc4cfe6478060df6a92441[0] ;
            Ied40f6b7847158bd08cbd932254dd6ba[0]  <=  I0aaea02d5fbc4cfe6478060df6a92441[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ibe5129eb30f626925a3ab5ed5e239bb3[0]        <=  I64476c4b13b6612ab90845870c8fcec6[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I64476c4b13b6612ab90845870c8fcec6[0] + 1 :
                                             I64476c4b13b6612ab90845870c8fcec6[0] ;
            I6ab04d323306b7290cc89ed66dbd93bf[0]  <=  I64476c4b13b6612ab90845870c8fcec6[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2a656dad40cec86a53e732e78f00c269[0]        <=  I46cb13c147e8087f9f93618f946d0f75[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I46cb13c147e8087f9f93618f946d0f75[0] + 1 :
                                             I46cb13c147e8087f9f93618f946d0f75[0] ;
            Iac4a5fdede87b021e6a8150d3bf34b66[0]  <=  I46cb13c147e8087f9f93618f946d0f75[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If06132c6a0060efdbd695b31c338faf6[0]        <=  Ida1dc39acb508dea4487357625f65a62[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ida1dc39acb508dea4487357625f65a62[0] + 1 :
                                             Ida1dc39acb508dea4487357625f65a62[0] ;
            Id92b1676e19c5818fa813d06dc9a01f3[0]  <=  Ida1dc39acb508dea4487357625f65a62[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I02fd20ab9e4fa12009b63fbe41d647fb[0]        <=  Ief0a83a4d2ab6337a9a842850ed9c8d2[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ief0a83a4d2ab6337a9a842850ed9c8d2[0] + 1 :
                                             Ief0a83a4d2ab6337a9a842850ed9c8d2[0] ;
            I93da1192f27c33e21e03b9a2748774ea[0]  <=  Ief0a83a4d2ab6337a9a842850ed9c8d2[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ibb97d541a2ed2b0cbad273a09fef5594[0]        <=  Iabc0481ca8b87650597db2ab82d9526a[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Iabc0481ca8b87650597db2ab82d9526a[0] + 1 :
                                             Iabc0481ca8b87650597db2ab82d9526a[0] ;
            I69a0c79d41af6b6340430b8b337fb0ca[0]  <=  Iabc0481ca8b87650597db2ab82d9526a[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0905c7e3678f66095194058bb72d22fe[0]        <=  I273daf63e8da53e5e9b99de802715b44[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I273daf63e8da53e5e9b99de802715b44[0] + 1 :
                                             I273daf63e8da53e5e9b99de802715b44[0] ;
            Ibd47f48d306ec44d94865a0a81e4f9dc[0]  <=  I273daf63e8da53e5e9b99de802715b44[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I81433ae67b7cb4dee0b2091f3819ea88[0]        <=  I9bec797aec01899ccab507296d7f4d53[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I9bec797aec01899ccab507296d7f4d53[0] + 1 :
                                             I9bec797aec01899ccab507296d7f4d53[0] ;
            Ia5707d1275138a5145b2a42190d95183[0]  <=  I9bec797aec01899ccab507296d7f4d53[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ia6249382442d1dd3062acc63f891465b[0]        <=  Id769ce05d2596a106b4e750d272b6d86[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Id769ce05d2596a106b4e750d272b6d86[0] + 1 :
                                             Id769ce05d2596a106b4e750d272b6d86[0] ;
            I33bc2f42d997a2963b063326eb210d1c[0]  <=  Id769ce05d2596a106b4e750d272b6d86[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie4bd4c14051455f00efdb023c3b58173[0]        <=  Ifcd0ef96ba3a7a7ef8ab4f64c5671f80[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ifcd0ef96ba3a7a7ef8ab4f64c5671f80[0] + 1 :
                                             Ifcd0ef96ba3a7a7ef8ab4f64c5671f80[0] ;
            Ib22e39b701614cd9986061c32adfbc66[0]  <=  Ifcd0ef96ba3a7a7ef8ab4f64c5671f80[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie64e67a2316af18c5835c3a32ae9290f[0]        <=  I2789f24264b92b82f7e9f34a5ccaa489[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I2789f24264b92b82f7e9f34a5ccaa489[0] + 1 :
                                             I2789f24264b92b82f7e9f34a5ccaa489[0] ;
            I9b08176fde1cd08c9d7686a659213580[0]  <=  I2789f24264b92b82f7e9f34a5ccaa489[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Icaf94b3fea3e29ff77d4793b389c9d14[0]        <=  Ic9f02e5a9bad9928c784d38980f709ff[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic9f02e5a9bad9928c784d38980f709ff[0] + 1 :
                                             Ic9f02e5a9bad9928c784d38980f709ff[0] ;
            I1b4e65357a818998d08b83d21584e18c[0]  <=  Ic9f02e5a9bad9928c784d38980f709ff[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I334991f6bfe06389e35b7a580982de1f[0]        <=  I5729f3c3121489f404f8964abb3e842a[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I5729f3c3121489f404f8964abb3e842a[0] + 1 :
                                             I5729f3c3121489f404f8964abb3e842a[0] ;
            Ibb865ea5891db706b7b54e5c6fa383d0[0]  <=  I5729f3c3121489f404f8964abb3e842a[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6390495458553670944cdbf57bd6ce7b[0]        <=  If076d265cc6b8f7baf4059ea5fa7525d[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~If076d265cc6b8f7baf4059ea5fa7525d[0] + 1 :
                                             If076d265cc6b8f7baf4059ea5fa7525d[0] ;
            I32d42cfd2d516af2e68fc2db4d5dce03[0]  <=  If076d265cc6b8f7baf4059ea5fa7525d[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ibafc73f0a3486943914e197a7af4505c[0]        <=  I7acc5316ae2768ce90598a82ad196eca[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I7acc5316ae2768ce90598a82ad196eca[0] + 1 :
                                             I7acc5316ae2768ce90598a82ad196eca[0] ;
            I4d0e8d475a5d2a7da24daca60f23f3d6[0]  <=  I7acc5316ae2768ce90598a82ad196eca[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2ec83b82756dda6035ddff10dd41fed5[0]        <=  Idc81e8df0b1b36ee2885c180c992a8db[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Idc81e8df0b1b36ee2885c180c992a8db[0] + 1 :
                                             Idc81e8df0b1b36ee2885c180c992a8db[0] ;
            Ie3850345b207e59aaaa5c944dab40b90[0]  <=  Idc81e8df0b1b36ee2885c180c992a8db[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5f6abb1000e5416dd4d43fcd052321fb[0]        <=  I2f587d7d70873b05956908ded54c36f9[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I2f587d7d70873b05956908ded54c36f9[0] + 1 :
                                             I2f587d7d70873b05956908ded54c36f9[0] ;
            I4a9a1c932db30dcf04cb105a8d7384f9[0]  <=  I2f587d7d70873b05956908ded54c36f9[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Icc865d7264dd89944317be21610dcf9d[0]        <=  I7f013f76d9fcc1b14984188e7af2ec0d[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I7f013f76d9fcc1b14984188e7af2ec0d[0] + 1 :
                                             I7f013f76d9fcc1b14984188e7af2ec0d[0] ;
            I0ef689822226332f5feaf79fcf8f6674[0]  <=  I7f013f76d9fcc1b14984188e7af2ec0d[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6a301412ef9235f3a609baf10a4200dd[0]        <=  Ica4903599938b7e1996702a51a7e9ec8[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ica4903599938b7e1996702a51a7e9ec8[0] + 1 :
                                             Ica4903599938b7e1996702a51a7e9ec8[0] ;
            Ib5744c2130bb5a9d0ccdd975fdf2ff9c[0]  <=  Ica4903599938b7e1996702a51a7e9ec8[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9840f42586460341bb39256726d39ca1[0]        <=  I53484a61ff8b4273d872779c33b292d5[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I53484a61ff8b4273d872779c33b292d5[0] + 1 :
                                             I53484a61ff8b4273d872779c33b292d5[0] ;
            I039a7ddcb25972501d80c45c938cf683[0]  <=  I53484a61ff8b4273d872779c33b292d5[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0837554bfb175a9ac8a4cb17e091fa9e[0]        <=  Iae00c13f4457b91d9a252b5b2aa67780[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Iae00c13f4457b91d9a252b5b2aa67780[0] + 1 :
                                             Iae00c13f4457b91d9a252b5b2aa67780[0] ;
            Ic5f36c15ebad061dfbd5301e02ce2ffe[0]  <=  Iae00c13f4457b91d9a252b5b2aa67780[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iacd698956b9ea6f1649063ee612c7e76[0]        <=  I208b29bdae3040b547e8e40ffdc96d34[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I208b29bdae3040b547e8e40ffdc96d34[0] + 1 :
                                             I208b29bdae3040b547e8e40ffdc96d34[0] ;
            Idf0d9dac06522293f8d7e00a93b6bbb5[0]  <=  I208b29bdae3040b547e8e40ffdc96d34[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I68928b2759202e358f75b08e162e6a68[0]        <=  Ic6378ae3bd73ac1ddfb25e7d7882c671[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic6378ae3bd73ac1ddfb25e7d7882c671[0] + 1 :
                                             Ic6378ae3bd73ac1ddfb25e7d7882c671[0] ;
            Id557db735a70dbb14504bc3088e8798e[0]  <=  Ic6378ae3bd73ac1ddfb25e7d7882c671[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I609f881624ec9034823c9f54f4fb9b6d[0]        <=  I81f95de60a5dd186e51f9f4bf0b624da[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I81f95de60a5dd186e51f9f4bf0b624da[0] + 1 :
                                             I81f95de60a5dd186e51f9f4bf0b624da[0] ;
            I150d31ef31093fdfc5f145d84bb35156[0]  <=  I81f95de60a5dd186e51f9f4bf0b624da[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I075a0a1afc1463e92edb5f7658395424[0]        <=  Ic05bdf0bf00ca3ba90c6ee7728b2d49b[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic05bdf0bf00ca3ba90c6ee7728b2d49b[0] + 1 :
                                             Ic05bdf0bf00ca3ba90c6ee7728b2d49b[0] ;
            I7e40e6f9d82d9b9fc546672e8e8621bb[0]  <=  Ic05bdf0bf00ca3ba90c6ee7728b2d49b[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Idf1030f0e2aa5e2605bcea5fbe0428f8[0]        <=  Ic74ef5ce41d9db0920015b60cd80dada[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic74ef5ce41d9db0920015b60cd80dada[0] + 1 :
                                             Ic74ef5ce41d9db0920015b60cd80dada[0] ;
            I14133cbbfa6521c5b81477fa1c229cbf[0]  <=  Ic74ef5ce41d9db0920015b60cd80dada[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1b82e98260c3bdeb5183a3af470e2d4a[0]        <=  If54ee451267f16296945fca60801b6da[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~If54ee451267f16296945fca60801b6da[0] + 1 :
                                             If54ee451267f16296945fca60801b6da[0] ;
            I3728e31a7cf48639ce873d9135dc87fb[0]  <=  If54ee451267f16296945fca60801b6da[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I75338af3ebc7b7061a499e98a5be1674[0]        <=  I22af03550c9ffd5ee75db6b34f444612[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I22af03550c9ffd5ee75db6b34f444612[0] + 1 :
                                             I22af03550c9ffd5ee75db6b34f444612[0] ;
            Ic6be12e390bd3c25c66d9b9e7c0532b8[0]  <=  I22af03550c9ffd5ee75db6b34f444612[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9f863d33f3c727e13eb52e7563ef9d1e[0]        <=  I76d5529e20b89a706595f65abe004da2[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I76d5529e20b89a706595f65abe004da2[0] + 1 :
                                             I76d5529e20b89a706595f65abe004da2[0] ;
            Icc50e1923274729fe472ca578b68c0f5[0]  <=  I76d5529e20b89a706595f65abe004da2[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I56b8e0a7e6d2229baa9908843c0208ce[0]        <=  Iebca060c7873173db59d0e1a244a5f62[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Iebca060c7873173db59d0e1a244a5f62[0] + 1 :
                                             Iebca060c7873173db59d0e1a244a5f62[0] ;
            I4d98064f544a41b977ba945d2eecdf21[0]  <=  Iebca060c7873173db59d0e1a244a5f62[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3d04bcd17aa2b98b69dcd671b9666c50[0]        <=  I39ebf0c6f66596aeb1c56eaf50bc6b55[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I39ebf0c6f66596aeb1c56eaf50bc6b55[0] + 1 :
                                             I39ebf0c6f66596aeb1c56eaf50bc6b55[0] ;
            I12f2a9f1e3e715d7e684ff39dd7942f0[0]  <=  I39ebf0c6f66596aeb1c56eaf50bc6b55[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id254880ed38db79c53facbdc0c4a6d1a[0]        <=  I685db637ba885fcd9a37a9457b56c827[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I685db637ba885fcd9a37a9457b56c827[0] + 1 :
                                             I685db637ba885fcd9a37a9457b56c827[0] ;
            Iaa4e3c53a0d55e8f42f60ff40893427e[0]  <=  I685db637ba885fcd9a37a9457b56c827[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I988a7c2c284c38fcd6682236dc2d6151[0]        <=  If659617a922c1800e53f789111d7f946[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~If659617a922c1800e53f789111d7f946[0] + 1 :
                                             If659617a922c1800e53f789111d7f946[0] ;
            I26aae317b0b320df86ca4004f64aab88[0]  <=  If659617a922c1800e53f789111d7f946[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ida4c48caeba43eccdddd1748824ec551[0]        <=  I3cde77dbb4b236619f7d00d6212d8f46[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I3cde77dbb4b236619f7d00d6212d8f46[0] + 1 :
                                             I3cde77dbb4b236619f7d00d6212d8f46[0] ;
            I9344825cc2e5864f691043a1f94f86a4[0]  <=  I3cde77dbb4b236619f7d00d6212d8f46[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If9936b476bb351a9ecbb97e2088cdd6f[0]        <=  Ic1f7f01098e573cdab8482bd3f0dfe0c[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic1f7f01098e573cdab8482bd3f0dfe0c[0] + 1 :
                                             Ic1f7f01098e573cdab8482bd3f0dfe0c[0] ;
            I82988c3879c1de76fe2140c469f6a4c1[0]  <=  Ic1f7f01098e573cdab8482bd3f0dfe0c[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6cbccfdeeb675a8a99d4c394bc8e71cd[0]        <=  Ic229657d83879de9bd470c1739254faa[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ic229657d83879de9bd470c1739254faa[0] + 1 :
                                             Ic229657d83879de9bd470c1739254faa[0] ;
            I6bdd8334512c7c6a3226ebb4e928a270[0]  <=  Ic229657d83879de9bd470c1739254faa[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I79a4a9dfcecca4073c101bdd9b738c7c[0]        <=  I3e69a3b20cf7ac74e77887b37fc3a5d7[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I3e69a3b20cf7ac74e77887b37fc3a5d7[0] + 1 :
                                             I3e69a3b20cf7ac74e77887b37fc3a5d7[0] ;
            I0debec6ace7160558cce7f111dd1bea6[0]  <=  I3e69a3b20cf7ac74e77887b37fc3a5d7[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ice57a50f53d13e7eaf25af23547b5fb0[0]        <=  Ief74f9042bd0058f17af181156b58456[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ief74f9042bd0058f17af181156b58456[0] + 1 :
                                             Ief74f9042bd0058f17af181156b58456[0] ;
            I8ee02e65ce9183683f0f3168bfd755c5[0]  <=  Ief74f9042bd0058f17af181156b58456[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8ff8106a70daac7c8932e88aeb6d198b[0]        <=  Ide1209ba9c80b0f69b0f17a1320b7a33[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ide1209ba9c80b0f69b0f17a1320b7a33[0] + 1 :
                                             Ide1209ba9c80b0f69b0f17a1320b7a33[0] ;
            I80e6d2c9c5f7b6bc6bffa063c4959115[0]  <=  Ide1209ba9c80b0f69b0f17a1320b7a33[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8f9d1ec03357f7f045196050511341a2[0]        <=  Ib8c08ba5cf3c7bd8233532cc8ecb4825[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ib8c08ba5cf3c7bd8233532cc8ecb4825[0] + 1 :
                                             Ib8c08ba5cf3c7bd8233532cc8ecb4825[0] ;
            I0f21fb041239a7a8895c9506f2754595[0]  <=  Ib8c08ba5cf3c7bd8233532cc8ecb4825[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic423bfa7639075130324da59f2cca2fc[0]        <=  I812e31439ca7c94df3d6bf578b60beaf[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I812e31439ca7c94df3d6bf578b60beaf[0] + 1 :
                                             I812e31439ca7c94df3d6bf578b60beaf[0] ;
            I8ce37a8e81b54043276835c11e394df5[0]  <=  I812e31439ca7c94df3d6bf578b60beaf[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I4eed402353a7fa22fcb11f2adbf6be03[0]        <=  Ie93978ee93511b6ed29aad9aed8ee903[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie93978ee93511b6ed29aad9aed8ee903[0] + 1 :
                                             Ie93978ee93511b6ed29aad9aed8ee903[0] ;
            Idf7d1f78735ce1e9695d99a532a7726e[0]  <=  Ie93978ee93511b6ed29aad9aed8ee903[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ieb579bed6711928456b296873c5da9cd[0]        <=  If0c12a1750d279b90738aacac5b35e04[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~If0c12a1750d279b90738aacac5b35e04[0] + 1 :
                                             If0c12a1750d279b90738aacac5b35e04[0] ;
            I96a552ed2d18c0ba3fc6cb6d6b6a0f44[0]  <=  If0c12a1750d279b90738aacac5b35e04[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ifdf316d14ef99080247091609b2c2a8f[0]        <=  I0501ec6e9230839738818ae2b19a5b65[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I0501ec6e9230839738818ae2b19a5b65[0] + 1 :
                                             I0501ec6e9230839738818ae2b19a5b65[0] ;
            I3c76936e8e3467378210a13645a401d4[0]  <=  I0501ec6e9230839738818ae2b19a5b65[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2a1afeffe5592e35349bfd4384de834e[0]        <=  I9e9c3529814bb741e0e425dba9ba0abf[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I9e9c3529814bb741e0e425dba9ba0abf[0] + 1 :
                                             I9e9c3529814bb741e0e425dba9ba0abf[0] ;
            Ic9a1d599fcfd5dd51265e5d0989719b6[0]  <=  I9e9c3529814bb741e0e425dba9ba0abf[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I93f88eac6c04d26228b5d7a3b1d00a42[0]        <=  I3898f311fc81d9bbcda50e18e7f978e1[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I3898f311fc81d9bbcda50e18e7f978e1[0] + 1 :
                                             I3898f311fc81d9bbcda50e18e7f978e1[0] ;
            I60156470e631268c392040d3c5582eca[0]  <=  I3898f311fc81d9bbcda50e18e7f978e1[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8c32ed7572af2a6a41a415ff6c580f3d[0]        <=  I4bf59374718f169f17fea6adb9d9c7e1[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I4bf59374718f169f17fea6adb9d9c7e1[0] + 1 :
                                             I4bf59374718f169f17fea6adb9d9c7e1[0] ;
            I821126d1516ad7e8191a7b2a3b5e4b47[0]  <=  I4bf59374718f169f17fea6adb9d9c7e1[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9cc4cd2860ebe1e5d43eb6024ea32dcf[0]        <=  Ide127cda229e55eca7ef703c0d794e6e[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ide127cda229e55eca7ef703c0d794e6e[0] + 1 :
                                             Ide127cda229e55eca7ef703c0d794e6e[0] ;
            Ibe72e9f6d2c3cbbcf98f6b5aa6a4f93b[0]  <=  Ide127cda229e55eca7ef703c0d794e6e[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I35b73e275ce37c06d10c227595c7c3f6[0]        <=  I482955b75319360d2646b1f712acdbde[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I482955b75319360d2646b1f712acdbde[0] + 1 :
                                             I482955b75319360d2646b1f712acdbde[0] ;
            I1e8b6306d2dfde4a36ee9b9c2caf1c85[0]  <=  I482955b75319360d2646b1f712acdbde[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iac4ee00e62d47494b2bfe3aff55506ea[0]        <=  I158984c3dfe52e5107e4aa64548c1ab5[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I158984c3dfe52e5107e4aa64548c1ab5[0] + 1 :
                                             I158984c3dfe52e5107e4aa64548c1ab5[0] ;
            I48ed92480f457fc3cc2ff0dd7d177a10[0]  <=  I158984c3dfe52e5107e4aa64548c1ab5[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6023ec90efcd1ac53ea71eeee1c996e2[0]        <=  Ibdfb487053f2567b45db76d12e9eb75a[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ibdfb487053f2567b45db76d12e9eb75a[0] + 1 :
                                             Ibdfb487053f2567b45db76d12e9eb75a[0] ;
            Iaed28d88a651f0151501ec4ea6ee3346[0]  <=  Ibdfb487053f2567b45db76d12e9eb75a[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6f2b0c5e254aeb7e967f86e914876171[0]        <=  I1fc2b706279a62a29d90f261f211c3a9[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I1fc2b706279a62a29d90f261f211c3a9[0] + 1 :
                                             I1fc2b706279a62a29d90f261f211c3a9[0] ;
            I9d94d9b5414662de841443d7866e66b1[0]  <=  I1fc2b706279a62a29d90f261f211c3a9[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie9353d9dd97f3536dfa6bcc2c662bf40[0]        <=  I988227c12ad87b2ced8fd8fd89eb138d[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I988227c12ad87b2ced8fd8fd89eb138d[0] + 1 :
                                             I988227c12ad87b2ced8fd8fd89eb138d[0] ;
            I870b8a3b11be215a8704ba05568f05e2[0]  <=  I988227c12ad87b2ced8fd8fd89eb138d[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I09fd28ae4656b1282feb899a40b9b233[0]        <=  Id537c7ec3b2e195d892f7fb1a63dcf46[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Id537c7ec3b2e195d892f7fb1a63dcf46[0] + 1 :
                                             Id537c7ec3b2e195d892f7fb1a63dcf46[0] ;
            Ia8bbf21e040b326058a9acb7d198a835[0]  <=  Id537c7ec3b2e195d892f7fb1a63dcf46[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iabbb1734d7e19cd9c7329b30cb26cd3b[0]        <=  I92a93c16158990f624973e9cc487fc00[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I92a93c16158990f624973e9cc487fc00[0] + 1 :
                                             I92a93c16158990f624973e9cc487fc00[0] ;
            Ie852f207c8f537621b080ffa0a89bfdc[0]  <=  I92a93c16158990f624973e9cc487fc00[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iacc03e49c3cd6749e4c49e13c8c8593e[0]        <=  Iab0879a7d17f0fbf2c2ed147e41d3f32[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Iab0879a7d17f0fbf2c2ed147e41d3f32[0] + 1 :
                                             Iab0879a7d17f0fbf2c2ed147e41d3f32[0] ;
            If53029b05bea46d656a6ef72fb6d6642[0]  <=  Iab0879a7d17f0fbf2c2ed147e41d3f32[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7913101e04088970adf3f1e7429cd06a[0]        <=  I762ebc964e606e803121e347086668e4[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I762ebc964e606e803121e347086668e4[0] + 1 :
                                             I762ebc964e606e803121e347086668e4[0] ;
            I8e8a740d09e000444ba1f4931b5cccf4[0]  <=  I762ebc964e606e803121e347086668e4[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ibddcea3450984eb0b3cc3ca6961fa646[0]        <=  I032010a0a18eaf23274cdff5c99442bc[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I032010a0a18eaf23274cdff5c99442bc[0] + 1 :
                                             I032010a0a18eaf23274cdff5c99442bc[0] ;
            I46605d823e06af5485e50b256b5c3f22[0]  <=  I032010a0a18eaf23274cdff5c99442bc[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0a863fcba425a8683ebbb35195ea70a4[0]        <=  I24956c032de466de716b6ab57dd8a265[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I24956c032de466de716b6ab57dd8a265[0] + 1 :
                                             I24956c032de466de716b6ab57dd8a265[0] ;
            I38344d68127f5c035193bb9030ce4d4d[0]  <=  I24956c032de466de716b6ab57dd8a265[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8138f45ab1b8a10869a2a6078b6c214c[0]        <=  If816e24bfd42448c3c0fb03b6e9e9404[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~If816e24bfd42448c3c0fb03b6e9e9404[0] + 1 :
                                             If816e24bfd42448c3c0fb03b6e9e9404[0] ;
            Iba9f33c08db89a7f120cc1e3eaf05dec[0]  <=  If816e24bfd42448c3c0fb03b6e9e9404[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie4c27f8574c8bad0b923796d2544f858[0]        <=  I0903046199323180f148f13aedaa0ab3[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I0903046199323180f148f13aedaa0ab3[0] + 1 :
                                             I0903046199323180f148f13aedaa0ab3[0] ;
            Ibde51eb91b3ca50a8a0513c94bd7be15[0]  <=  I0903046199323180f148f13aedaa0ab3[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ibea29d15c71d594e4e9cbe6a58ebc550[0]        <=  I25ec8dfa866fe300e67a01944f893bf6[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I25ec8dfa866fe300e67a01944f893bf6[0] + 1 :
                                             I25ec8dfa866fe300e67a01944f893bf6[0] ;
            Ifb94196d1653a0166567e170f06ec0db[0]  <=  I25ec8dfa866fe300e67a01944f893bf6[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0b249349485591abcc09c4587efca78d[0]        <=  I77ac8c7c5ea03d948931590d57c8d649[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I77ac8c7c5ea03d948931590d57c8d649[0] + 1 :
                                             I77ac8c7c5ea03d948931590d57c8d649[0] ;
            I9cf7557e2cac4532a77fcb212712db0f[0]  <=  I77ac8c7c5ea03d948931590d57c8d649[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6bbe05bfdabac8f312c7800eca53be62[0]        <=  Ief5d16bc74276d3aec10a56fe8234b8a[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ief5d16bc74276d3aec10a56fe8234b8a[0] + 1 :
                                             Ief5d16bc74276d3aec10a56fe8234b8a[0] ;
            I3159d7faeee1a904c409bde1967d2c21[0]  <=  Ief5d16bc74276d3aec10a56fe8234b8a[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie28e38c9881297e7ffae5c3aed4dfdd3[0]        <=  I6bec62410ca887855fafaa4be4c09d72[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I6bec62410ca887855fafaa4be4c09d72[0] + 1 :
                                             I6bec62410ca887855fafaa4be4c09d72[0] ;
            I35dfb5ece5e04504d6e74739ae99c9cc[0]  <=  I6bec62410ca887855fafaa4be4c09d72[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1358b8ab0933bd596c33b622d2f9523f[0]        <=  I290223476b30aa41df98af3016119109[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I290223476b30aa41df98af3016119109[0] + 1 :
                                             I290223476b30aa41df98af3016119109[0] ;
            Iabff939ae4acf7d7b038e028c29b6166[0]  <=  I290223476b30aa41df98af3016119109[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I46ce01ea907e88cafb7d96d22b5fffd6[0]        <=  I07e3ae59ec05fa46d6ca3398a42e287c[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I07e3ae59ec05fa46d6ca3398a42e287c[0] + 1 :
                                             I07e3ae59ec05fa46d6ca3398a42e287c[0] ;
            Ia14159444578c6dc88f2d5ea0317774b[0]  <=  I07e3ae59ec05fa46d6ca3398a42e287c[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I64c0e39b2f3c34d724ecf0f511a413c9[0]        <=  I7b019b5e5991ad8497a048367d83341f[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I7b019b5e5991ad8497a048367d83341f[0] + 1 :
                                             I7b019b5e5991ad8497a048367d83341f[0] ;
            Ie2306a5c441d621388b73195027fc118[0]  <=  I7b019b5e5991ad8497a048367d83341f[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6ffbd03867a92aea248506af197c2e86[0]        <=  I80f8ed713e4b0281f94804a0b66fadcf[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I80f8ed713e4b0281f94804a0b66fadcf[0] + 1 :
                                             I80f8ed713e4b0281f94804a0b66fadcf[0] ;
            I700a0fbf81e57d4970ce07090ec4f2e2[0]  <=  I80f8ed713e4b0281f94804a0b66fadcf[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie0a0c3e63be2145dc838faf227a84044[0]        <=  I8cd2472defb068d6e3af7070c97c25ef[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I8cd2472defb068d6e3af7070c97c25ef[0] + 1 :
                                             I8cd2472defb068d6e3af7070c97c25ef[0] ;
            I6007914b3fb3011c3ab2f9a9d7794ab2[0]  <=  I8cd2472defb068d6e3af7070c97c25ef[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I58265e8a07eede7063d5a80db2412214[0]        <=  I3689f559a9636f9dd4558e99424d6c80[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I3689f559a9636f9dd4558e99424d6c80[0] + 1 :
                                             I3689f559a9636f9dd4558e99424d6c80[0] ;
            I2096f40fe62e9d6f1ff96f258ffdbe33[0]  <=  I3689f559a9636f9dd4558e99424d6c80[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6734d5f87b795f4a05510778c22b555c[0]        <=  I77c454b260ff3c291b59ac8679966ab1[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I77c454b260ff3c291b59ac8679966ab1[0] + 1 :
                                             I77c454b260ff3c291b59ac8679966ab1[0] ;
            I93d8b7a24702bacbfc528242991516a9[0]  <=  I77c454b260ff3c291b59ac8679966ab1[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I314ced88cfc50d8b2edf129a6a3bf1a6[0]        <=  Iddb9b8c346479631362bfc4aa039b746[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Iddb9b8c346479631362bfc4aa039b746[0] + 1 :
                                             Iddb9b8c346479631362bfc4aa039b746[0] ;
            If0863fae91b2ec980ebdb26cfc90ae2e[0]  <=  Iddb9b8c346479631362bfc4aa039b746[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8cc6f1dc58a26262f18f334b751385ea[0]        <=  I3db9cdf51e4437b6e979f8c1a0be96df[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I3db9cdf51e4437b6e979f8c1a0be96df[0] + 1 :
                                             I3db9cdf51e4437b6e979f8c1a0be96df[0] ;
            I9ec29a319384efd562c2337e1857cb4e[0]  <=  I3db9cdf51e4437b6e979f8c1a0be96df[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I18d34c481f17aae6b16b6d0a5aa85357[0]        <=  I2a2352cab4f2edc64f156ef7b5e5595b[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I2a2352cab4f2edc64f156ef7b5e5595b[0] + 1 :
                                             I2a2352cab4f2edc64f156ef7b5e5595b[0] ;
            Ia56ecc024eae608d7de1509d75139dc2[0]  <=  I2a2352cab4f2edc64f156ef7b5e5595b[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib54b35abe1088393d275f4f45f7ed966[0]        <=  Iee3314c9bfca7066dcbb138d5f46d1f8[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Iee3314c9bfca7066dcbb138d5f46d1f8[0] + 1 :
                                             Iee3314c9bfca7066dcbb138d5f46d1f8[0] ;
            Iebcd65ea41cd38bfe3c8577277809acd[0]  <=  Iee3314c9bfca7066dcbb138d5f46d1f8[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie339493197828e5bd69bc49ca91aeb1d[0]        <=  I4883185d078ac45e5eb2d6dbcd2c875b[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I4883185d078ac45e5eb2d6dbcd2c875b[0] + 1 :
                                             I4883185d078ac45e5eb2d6dbcd2c875b[0] ;
            I75be12b14694ebcb5aff6e5d3e576315[0]  <=  I4883185d078ac45e5eb2d6dbcd2c875b[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic5084e34e9626f2e423283a87ea0d91d[0]        <=  Ie6242ba25d061a37a41d7ca41370e919[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Ie6242ba25d061a37a41d7ca41370e919[0] + 1 :
                                             Ie6242ba25d061a37a41d7ca41370e919[0] ;
            I8e06fe414cd04103baf3882771a63e2c[0]  <=  Ie6242ba25d061a37a41d7ca41370e919[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3fee16f7ef907bcf1e2f5b2e7ec77866[0]        <=  I99d9fb1f21a8aba32da690b3bbb786df[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I99d9fb1f21a8aba32da690b3bbb786df[0] + 1 :
                                             I99d9fb1f21a8aba32da690b3bbb786df[0] ;
            I0fe8574049166c363c7cc816b1435009[0]  <=  I99d9fb1f21a8aba32da690b3bbb786df[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iee529a0d30e79cdc9b33dd3d876a0f23[0]        <=  I1328d62797b528de9c98372d828d4af0[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I1328d62797b528de9c98372d828d4af0[0] + 1 :
                                             I1328d62797b528de9c98372d828d4af0[0] ;
            Id5f435c07240d5fe4a0e48c8f25ad0b7[0]  <=  I1328d62797b528de9c98372d828d4af0[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6c7373fafcfbb14c527e38e0f4440404[0]        <=  Id71c488586e019260c79018420d61673[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~Id71c488586e019260c79018420d61673[0] + 1 :
                                             Id71c488586e019260c79018420d61673[0] ;
            I1ae21e0db88f955c4f08f6d52f58974d[0]  <=  Id71c488586e019260c79018420d61673[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ided1b79349f8806da8f5c6898cea94bc[0]        <=  I6f2d4122c89e56e6640df3cec76c3c48[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I6f2d4122c89e56e6640df3cec76c3c48[0] + 1 :
                                             I6f2d4122c89e56e6640df3cec76c3c48[0] ;
            I92efddd59e1ea92902a295c0b8385c68[0]  <=  I6f2d4122c89e56e6640df3cec76c3c48[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id77e3ee5aded95fe141c26ad08639538[0]        <=  I37d02ddb7b52ae3495a3a182a3d4708a[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I37d02ddb7b52ae3495a3a182a3d4708a[0] + 1 :
                                             I37d02ddb7b52ae3495a3a182a3d4708a[0] ;
            I56948ad2b2cc245bb1003fd71ae5f899[0]  <=  I37d02ddb7b52ae3495a3a182a3d4708a[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3c286283659a38021c27b5e5346b59b0[0]        <=  I30b006cb2cf34c967066041123ac3698[0][SIGN_MAX_SUM_WDTH_LONG] ?
                                             ~I30b006cb2cf34c967066041123ac3698[0] + 1 :
                                             I30b006cb2cf34c967066041123ac3698[0] ;
            I5fb5081b7a2da89115c0080b0967974d[0]  <=  I30b006cb2cf34c967066041123ac3698[0][SIGN_MAX_SUM_WDTH_LONG] ;
           end
       end

   end

assign I583b1bfc712ec29d08acc68c27675882[0]      = I748f85f6680918a2e992df339b4b6558 +  ~Iea07d1adf9016a29cffd61d183e268d0 +1;
assign I583b1bfc712ec29d08acc68c27675882[1]      = I748f85f6680918a2e992df339b4b6558 +  ~If92db65b39a83e1c699e4cc6d7f9e57b +1;
assign I583b1bfc712ec29d08acc68c27675882[2]      = I748f85f6680918a2e992df339b4b6558 +  ~I8f2986bc015fcc64ac5e5395ac6dd851 +1;
assign I583b1bfc712ec29d08acc68c27675882[3]      = I748f85f6680918a2e992df339b4b6558 +  ~I355725a804e0df68b4acf96ca98f2448 +1;
assign I583b1bfc712ec29d08acc68c27675882[4]      = I748f85f6680918a2e992df339b4b6558 +  ~I78212ae965ab2dcb2eed0b060d6b253f +1;
assign I583b1bfc712ec29d08acc68c27675882[5]      = I748f85f6680918a2e992df339b4b6558 +  ~I0b56aa7a1b7549c91dddd3a06ecbaacf +1;
assign I583b1bfc712ec29d08acc68c27675882[6]      = I748f85f6680918a2e992df339b4b6558 +  ~I71412803cc5229025487255aec62ec4f +1;
assign I583b1bfc712ec29d08acc68c27675882[7]      = I748f85f6680918a2e992df339b4b6558 +  ~I32fcb28a27356bc6f403528836ea4c1f +1;
assign I583b1bfc712ec29d08acc68c27675882[8]      = I748f85f6680918a2e992df339b4b6558 +  ~Iad354d876cb9fc72fc0143e6f7da9357 +1;
assign I583b1bfc712ec29d08acc68c27675882[9]      = I748f85f6680918a2e992df339b4b6558 +  ~If6e745bb85abba7282dae1f6f701225e +1;
assign I583b1bfc712ec29d08acc68c27675882[10]      = I748f85f6680918a2e992df339b4b6558 +  ~I93bb43c1b89d4c70a57bdc019d64fd22 +1;
assign I583b1bfc712ec29d08acc68c27675882[11]      = I748f85f6680918a2e992df339b4b6558 +  ~I7a2e554d07bbea291f2cfc18694fca3a +1;
assign I583b1bfc712ec29d08acc68c27675882[12]      = I748f85f6680918a2e992df339b4b6558 +  ~I3e59b2419c7dd1553b792d536208514e +1;
assign I583b1bfc712ec29d08acc68c27675882[13]      = I748f85f6680918a2e992df339b4b6558 +  ~I46894c6526983bf1ce4b503159131b41 +1;
assign I583b1bfc712ec29d08acc68c27675882[14]      = I748f85f6680918a2e992df339b4b6558 +  ~I6404d0df952b5bf8292c753e4c6f35d8 +1;
assign I583b1bfc712ec29d08acc68c27675882[15]      = I748f85f6680918a2e992df339b4b6558 +  ~I8522c402e654d007abffcb0e904af5e6 +1;
assign I583b1bfc712ec29d08acc68c27675882[16]      = I748f85f6680918a2e992df339b4b6558 +  ~I5ed85845c39337c37791f16e718069b4 +1;
assign I583b1bfc712ec29d08acc68c27675882[17]      = I748f85f6680918a2e992df339b4b6558 +  ~I89013d61c1ea8da8b1c6071cc21c316f +1;
assign I583b1bfc712ec29d08acc68c27675882[18]      = I748f85f6680918a2e992df339b4b6558 +  ~I4102100fa5f1dd299af0190862efcc42 +1;
assign I583b1bfc712ec29d08acc68c27675882[19]      = I748f85f6680918a2e992df339b4b6558 +  ~I4939f69abb1eac56d5021e06406a93b5 +1;
assign I583b1bfc712ec29d08acc68c27675882[20]      = I748f85f6680918a2e992df339b4b6558 +  ~Iadbd245bf842aebb456417579a3e6296 +1;
assign I583b1bfc712ec29d08acc68c27675882[21]      = I748f85f6680918a2e992df339b4b6558 +  ~Ifc8ece44a4e68c3117eda9e65f3084d2 +1;
assign Ifba287889bea3585954fef5efdf5bb24[0]      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~I91679dfab57a372eddc7f9b94a231edb +1;
assign Ifba287889bea3585954fef5efdf5bb24[1]      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~I2213c1a2b831f421707a261f5a58b1b1 +1;
assign Ifba287889bea3585954fef5efdf5bb24[2]      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~Ic53b875b2ddcba11406eb2ca39354757 +1;
assign Ifba287889bea3585954fef5efdf5bb24[3]      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~I634484f00590216c0f74f975c9c83400 +1;
assign Ifba287889bea3585954fef5efdf5bb24[4]      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~Ib3b1db2d8b669988c887ed780e439b26 +1;
assign Ifba287889bea3585954fef5efdf5bb24[5]      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~I735db8b0ee0ec98e4cce0030b11508da +1;
assign Ifba287889bea3585954fef5efdf5bb24[6]      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~If1607e907e626902ee26d15020a64c21 +1;
assign Ifba287889bea3585954fef5efdf5bb24[7]      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~I081b38dbb37d4c14a6a9fd3fefa13daa +1;
assign Ifba287889bea3585954fef5efdf5bb24[8]      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~Ibac5e7b6d4bf5cd6926358318f0c418f +1;
assign Ifba287889bea3585954fef5efdf5bb24[9]      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~Iadfc60386481092ae85cc148a2c40abb +1;
assign Ifba287889bea3585954fef5efdf5bb24[10]      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~Ie0ee5445c56a5f9b41640b57422206de +1;
assign Ifba287889bea3585954fef5efdf5bb24[11]      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~Ie5f8620371236cb11c9e88c16b509ee8 +1;
assign Ifba287889bea3585954fef5efdf5bb24[12]      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~I8d7c1fe2e33bbd45379b0325a3c5e989 +1;
assign Ifba287889bea3585954fef5efdf5bb24[13]      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~I4fbdc4ee57a3be42b62d9bd43078d6ef +1;
assign Ifba287889bea3585954fef5efdf5bb24[14]      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~I5510b88bfd65811b3200adf4ef975b48 +1;
assign Ifba287889bea3585954fef5efdf5bb24[15]      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~Ib57ef2f577cca54713c16717cbbd1ce9 +1;
assign Ifba287889bea3585954fef5efdf5bb24[16]      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~I15943aa74e9fbbaebdc0d54eb6a3bffa +1;
assign Ifba287889bea3585954fef5efdf5bb24[17]      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~I6ac24c46319a787daa5c545de8c6eeea +1;
assign Ifba287889bea3585954fef5efdf5bb24[18]      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~I52403a0454e5fa002e79eaab7ea497bd +1;
assign Ifba287889bea3585954fef5efdf5bb24[19]      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~I634f0ce28934600a1a31ab0d8e59b4a9 +1;
assign Ifba287889bea3585954fef5efdf5bb24[20]      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~I7103aa739616a39c03e675ea0efb0335 +1;
assign Ifba287889bea3585954fef5efdf5bb24[21]      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~I0296d01fd3f9a269a617efd4beea9b8b +1;
assign I8e5ae9e6fa38cea8e5d320fe582c0729[0]      = If75e99660e3997f53f7b903bc366f47f +  ~I065a81ba25962785215583e7ece27661 +1;
assign I8e5ae9e6fa38cea8e5d320fe582c0729[1]      = If75e99660e3997f53f7b903bc366f47f +  ~I631a3300cb6685f47da7781940ec5d27 +1;
assign I8e5ae9e6fa38cea8e5d320fe582c0729[2]      = If75e99660e3997f53f7b903bc366f47f +  ~I8bbe1a2ace8f51aa22cca5d9fc66f136 +1;
assign I8e5ae9e6fa38cea8e5d320fe582c0729[3]      = If75e99660e3997f53f7b903bc366f47f +  ~I38c3e3e136acb79c8a0ff850bcc55f16 +1;
assign I8e5ae9e6fa38cea8e5d320fe582c0729[4]      = If75e99660e3997f53f7b903bc366f47f +  ~I35b2c7e9cdc53a98913e1c16a3a47b37 +1;
assign I8e5ae9e6fa38cea8e5d320fe582c0729[5]      = If75e99660e3997f53f7b903bc366f47f +  ~Ib1a2b31d49ae476e2f1fb9acba2d5af0 +1;
assign I8e5ae9e6fa38cea8e5d320fe582c0729[6]      = If75e99660e3997f53f7b903bc366f47f +  ~Ic72f41f9bbf470aee3c9b9b8787b31c3 +1;
assign I8e5ae9e6fa38cea8e5d320fe582c0729[7]      = If75e99660e3997f53f7b903bc366f47f +  ~I3ea4c33a9419820ed54460eb64134dff +1;
assign I8e5ae9e6fa38cea8e5d320fe582c0729[8]      = If75e99660e3997f53f7b903bc366f47f +  ~Ia0d940e16c8cbd4f7544f5a5cd7d83b2 +1;
assign I8e5ae9e6fa38cea8e5d320fe582c0729[9]      = If75e99660e3997f53f7b903bc366f47f +  ~I4a8abfa0896ce414d9b98093ef84455f +1;
assign I8e5ae9e6fa38cea8e5d320fe582c0729[10]      = If75e99660e3997f53f7b903bc366f47f +  ~I680be647bf2a62e0ee9b5d379dc87b4f +1;
assign I8e5ae9e6fa38cea8e5d320fe582c0729[11]      = If75e99660e3997f53f7b903bc366f47f +  ~If4d75f83299a21802b6fbe136913489f +1;
assign I8e5ae9e6fa38cea8e5d320fe582c0729[12]      = If75e99660e3997f53f7b903bc366f47f +  ~Ibddfda6413e3dd2f483c3174ea836b6a +1;
assign I8e5ae9e6fa38cea8e5d320fe582c0729[13]      = If75e99660e3997f53f7b903bc366f47f +  ~I33bddb0adcc2af7b12a83bf843036385 +1;
assign I8e5ae9e6fa38cea8e5d320fe582c0729[14]      = If75e99660e3997f53f7b903bc366f47f +  ~I529f92b82248efe2cf64f7da0ec8283c +1;
assign I8e5ae9e6fa38cea8e5d320fe582c0729[15]      = If75e99660e3997f53f7b903bc366f47f +  ~I2f34af0036985cd94ade9cc905bec065 +1;
assign I8e5ae9e6fa38cea8e5d320fe582c0729[16]      = If75e99660e3997f53f7b903bc366f47f +  ~Ia1a0d8d7dfd6e877f15cce773f85f5b7 +1;
assign I8e5ae9e6fa38cea8e5d320fe582c0729[17]      = If75e99660e3997f53f7b903bc366f47f +  ~I5dd29fd1a73df5662d2b636e7285bad9 +1;
assign I8e5ae9e6fa38cea8e5d320fe582c0729[18]      = If75e99660e3997f53f7b903bc366f47f +  ~Ide530e6f4622c8a7b101b6dce9650e42 +1;
assign I8e5ae9e6fa38cea8e5d320fe582c0729[19]      = If75e99660e3997f53f7b903bc366f47f +  ~Ibaf00a6780325882067a79f0c4d693d2 +1;
assign I8e5ae9e6fa38cea8e5d320fe582c0729[20]      = If75e99660e3997f53f7b903bc366f47f +  ~I16e3559c63ebfed83d6698fc9a9cd93a +1;
assign I8e5ae9e6fa38cea8e5d320fe582c0729[21]      = If75e99660e3997f53f7b903bc366f47f +  ~I9747a02384abb1c2dd1f52b3a5a999cc +1;
assign I67315420a608e257df8cfb520ef9f0a1[0]      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~Iceb7a1d4c23806b8f5824016779ad129 +1;
assign I67315420a608e257df8cfb520ef9f0a1[1]      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~I40ef50004a60ae58aedc49eb5e6797c9 +1;
assign I67315420a608e257df8cfb520ef9f0a1[2]      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~I753f92da60980736440aba814a156f1e +1;
assign I67315420a608e257df8cfb520ef9f0a1[3]      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~I4ac79b67a8904b95f7912d24af420585 +1;
assign I67315420a608e257df8cfb520ef9f0a1[4]      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~Iad44c932cfa5c249c5e59f8c706173a8 +1;
assign I67315420a608e257df8cfb520ef9f0a1[5]      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~I10f14b6433498e3b9e9bf021b60115e8 +1;
assign I67315420a608e257df8cfb520ef9f0a1[6]      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~I96008f47b9f134c9c4274cfcfb28e550 +1;
assign I67315420a608e257df8cfb520ef9f0a1[7]      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~Id0344146d1a53d418add6d2b185377dd +1;
assign I67315420a608e257df8cfb520ef9f0a1[8]      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~I1eede74f12d37331b399eb7136bc621f +1;
assign I67315420a608e257df8cfb520ef9f0a1[9]      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~I3e4754acc31d99bc71525789bdee0c1a +1;
assign I67315420a608e257df8cfb520ef9f0a1[10]      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~I11c1fc94a3bd6dffa17e1571cc6ae97c +1;
assign I67315420a608e257df8cfb520ef9f0a1[11]      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~I5395ee57418c31e11cf847f0f514ec19 +1;
assign I67315420a608e257df8cfb520ef9f0a1[12]      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~Iff125392fa39afebae1637a19c4e23ec +1;
assign I67315420a608e257df8cfb520ef9f0a1[13]      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~Ia6308e16fae5428f4ab6560f5b21479a +1;
assign I67315420a608e257df8cfb520ef9f0a1[14]      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~I5ea02b5349cd4d99ccbcb6b26f0cfdd7 +1;
assign I67315420a608e257df8cfb520ef9f0a1[15]      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~I21de4f6194dec9e3c401934db92c25e7 +1;
assign I67315420a608e257df8cfb520ef9f0a1[16]      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~I57d0920119f8901bd4dea2d5f8fb5d90 +1;
assign I67315420a608e257df8cfb520ef9f0a1[17]      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~I89537301987d6da0dbe6cff3caab3ff4 +1;
assign I67315420a608e257df8cfb520ef9f0a1[18]      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~Iaf0bbbe791bb71d0f557dc71caa5fb87 +1;
assign I67315420a608e257df8cfb520ef9f0a1[19]      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~Ic7ff9cde71054c1ee9eef81eabdd7061 +1;
assign I67315420a608e257df8cfb520ef9f0a1[20]      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~I88c10c47ae424fbdcb852fbf1e94127c +1;
assign I67315420a608e257df8cfb520ef9f0a1[21]      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~Icd2e75e47cab1d539ba9ff1b6e1d7155 +1;
assign Ic80a23c7b47f2236087fd7818d8d7c7f[0]      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~I37e6bc7aff363ed0ed1f84b23c5f3e34 +1;
assign Ic80a23c7b47f2236087fd7818d8d7c7f[1]      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~I733605337bf6972630c089d32fd7f98f +1;
assign Ic80a23c7b47f2236087fd7818d8d7c7f[2]      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~Idcb1d8bbdeaed6768c2a418c3048e6ee +1;
assign Ic80a23c7b47f2236087fd7818d8d7c7f[3]      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~Ia89da2f1890524ad3519ab403dd0686c +1;
assign Ic80a23c7b47f2236087fd7818d8d7c7f[4]      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~Ie33a780b0221084898c9fc5b237b244a +1;
assign Ic80a23c7b47f2236087fd7818d8d7c7f[5]      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~Iabbd1668e0014df518ede5216232834c +1;
assign Ic80a23c7b47f2236087fd7818d8d7c7f[6]      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~Ibd89458312687610aa166a9538968851 +1;
assign Ic80a23c7b47f2236087fd7818d8d7c7f[7]      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~Icbaf92a8e9875bcb19a1d074779a9ea5 +1;
assign Ic80a23c7b47f2236087fd7818d8d7c7f[8]      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~I80f3c8559da8e97bc5397bb8b621a0bd +1;
assign Ic80a23c7b47f2236087fd7818d8d7c7f[9]      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~I7a0eada108891aba06cecab5071232c9 +1;
assign Ic80a23c7b47f2236087fd7818d8d7c7f[10]      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~Ie21a2c9b22e7bf8425fb5c0f33e5f4f7 +1;
assign Ic80a23c7b47f2236087fd7818d8d7c7f[11]      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~Iaa5b2807e5cc2403c5787eeb3d10ca6b +1;
assign Ic80a23c7b47f2236087fd7818d8d7c7f[12]      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~I6da2b3a481ee71b85f3087b36b399288 +1;
assign Ic80a23c7b47f2236087fd7818d8d7c7f[13]      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~I11094e852295755925c3c61f1df81643 +1;
assign Ic80a23c7b47f2236087fd7818d8d7c7f[14]      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~I9c633aa620cca127b0ff8cf882178e76 +1;
assign Ic80a23c7b47f2236087fd7818d8d7c7f[15]      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~I694d471fd353eb54aae08a2afa7b645a +1;
assign Ic80a23c7b47f2236087fd7818d8d7c7f[16]      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~I816704585ad393f685731104ad3ec64f +1;
assign Ic80a23c7b47f2236087fd7818d8d7c7f[17]      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~I85d95015a9ce27a18ccbf73bbbcdbd70 +1;
assign Ic80a23c7b47f2236087fd7818d8d7c7f[18]      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~I992e7c551b4aa818606c3465d33eb798 +1;
assign Ic80a23c7b47f2236087fd7818d8d7c7f[19]      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~I2ead0e9941e2280309ab53535b1e1ac1 +1;
assign Ic80a23c7b47f2236087fd7818d8d7c7f[20]      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~I56873feb8418005b5661c7382f2dbeec +1;
assign Ic80a23c7b47f2236087fd7818d8d7c7f[21]      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~Ib6ea4a822da2ea32e0abf6cf8a33d295 +1;
assign Ic80a23c7b47f2236087fd7818d8d7c7f[22]      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~Id1659ccdeaea3e59eb2d3f65a65ebd05 +1;
assign Ie53d62e3ef9caf35092d7a63be1f565f[0]      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~Ic2171967791a0329f3e39fc19d0a6bc8 +1;
assign Ie53d62e3ef9caf35092d7a63be1f565f[1]      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~I7d5041a6796c00188f74936d283defe6 +1;
assign Ie53d62e3ef9caf35092d7a63be1f565f[2]      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~Iba7608ee0a01af103e022bcaf564bf6b +1;
assign Ie53d62e3ef9caf35092d7a63be1f565f[3]      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~Iedbe9d0e48bd36064f59faea51afddb9 +1;
assign Ie53d62e3ef9caf35092d7a63be1f565f[4]      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~Ic3871325d57b310c95ca02fcaca529eb +1;
assign Ie53d62e3ef9caf35092d7a63be1f565f[5]      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~I42f9b1f8ef24ad56c10086852678b456 +1;
assign Ie53d62e3ef9caf35092d7a63be1f565f[6]      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~I3ed5d0fca86f35b3d4b4a89c6147d0cd +1;
assign Ie53d62e3ef9caf35092d7a63be1f565f[7]      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~Ib0126fb335e32793c400a97c5a4a337c +1;
assign Ie53d62e3ef9caf35092d7a63be1f565f[8]      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~I20590d8fb97ec0b2164ffe17826136a7 +1;
assign Ie53d62e3ef9caf35092d7a63be1f565f[9]      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~I3c128efc9f80c9b8334bf7b61de71b43 +1;
assign Ie53d62e3ef9caf35092d7a63be1f565f[10]      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~Ic7147944f8835e26b9838fdbdc18ca41 +1;
assign Ie53d62e3ef9caf35092d7a63be1f565f[11]      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~I698b1dbc9d8664d1c86c7a763d97b3b7 +1;
assign Ie53d62e3ef9caf35092d7a63be1f565f[12]      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~I508bbade361787127e1a2e8687ec884c +1;
assign Ie53d62e3ef9caf35092d7a63be1f565f[13]      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~I2afeb2a7b199c0c6738938f156ae4274 +1;
assign Ie53d62e3ef9caf35092d7a63be1f565f[14]      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~I86255756ddd1f88b74e070b19f8c3bfa +1;
assign Ie53d62e3ef9caf35092d7a63be1f565f[15]      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~I7d4924388dc5373ad7936dca76797473 +1;
assign Ie53d62e3ef9caf35092d7a63be1f565f[16]      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~Ie317e5ea2ca4ba2060d0f491290af96f +1;
assign Ie53d62e3ef9caf35092d7a63be1f565f[17]      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~I56ea52c50a188ec47e48740839a031c9 +1;
assign Ie53d62e3ef9caf35092d7a63be1f565f[18]      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~Id9b9a8fe43992ec0793845715dd2226c +1;
assign Ie53d62e3ef9caf35092d7a63be1f565f[19]      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~I93b69bfb228db4b569a6772179d603be +1;
assign Ie53d62e3ef9caf35092d7a63be1f565f[20]      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~I71afab29cdb962e1f1ca21b61dfb50c6 +1;
assign Ie53d62e3ef9caf35092d7a63be1f565f[21]      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~I9905e2686b350e8a6e7f790563a91294 +1;
assign Ie53d62e3ef9caf35092d7a63be1f565f[22]      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~I524e78ae6a4204e17ba4532dba047d4b +1;
assign Ia73bc9712b861f909d0e3683ec91ea1c[0]      = Id7699f8f89380c315303644fdebacb32 +  ~I71228fe4188ab1d9796081184a422094 +1;
assign Ia73bc9712b861f909d0e3683ec91ea1c[1]      = Id7699f8f89380c315303644fdebacb32 +  ~Ie19b39200436b0bfca13502ad36c21b9 +1;
assign Ia73bc9712b861f909d0e3683ec91ea1c[2]      = Id7699f8f89380c315303644fdebacb32 +  ~If6657f90c84ca5e2ba08ec705f34be03 +1;
assign Ia73bc9712b861f909d0e3683ec91ea1c[3]      = Id7699f8f89380c315303644fdebacb32 +  ~I60ec7459bbe99fce295406bee1f2af46 +1;
assign Ia73bc9712b861f909d0e3683ec91ea1c[4]      = Id7699f8f89380c315303644fdebacb32 +  ~I29ab844f80c105d247c5c15faa35863c +1;
assign Ia73bc9712b861f909d0e3683ec91ea1c[5]      = Id7699f8f89380c315303644fdebacb32 +  ~I856fa68463aa5ef1ae53442699d38b33 +1;
assign Ia73bc9712b861f909d0e3683ec91ea1c[6]      = Id7699f8f89380c315303644fdebacb32 +  ~Ic3d00a27f15f8983a120395082854d6b +1;
assign Ia73bc9712b861f909d0e3683ec91ea1c[7]      = Id7699f8f89380c315303644fdebacb32 +  ~I6b1d01c3cb8fb51e43cdb788b89816be +1;
assign Ia73bc9712b861f909d0e3683ec91ea1c[8]      = Id7699f8f89380c315303644fdebacb32 +  ~Ib74a56900c1f8b159ad381f61acee801 +1;
assign Ia73bc9712b861f909d0e3683ec91ea1c[9]      = Id7699f8f89380c315303644fdebacb32 +  ~Ia5eba52d169755c507b9e0094e467fab +1;
assign Ia73bc9712b861f909d0e3683ec91ea1c[10]      = Id7699f8f89380c315303644fdebacb32 +  ~I0899e8fec1a7209cd94757c0b2f87c9a +1;
assign Ia73bc9712b861f909d0e3683ec91ea1c[11]      = Id7699f8f89380c315303644fdebacb32 +  ~I08ece7cd684e593e02321612b7a88cee +1;
assign Ia73bc9712b861f909d0e3683ec91ea1c[12]      = Id7699f8f89380c315303644fdebacb32 +  ~I691c84d81c60a462e28e2b2bae3ea845 +1;
assign Ia73bc9712b861f909d0e3683ec91ea1c[13]      = Id7699f8f89380c315303644fdebacb32 +  ~I58dc9cce6384160c0a85c6efb3319cdb +1;
assign Ia73bc9712b861f909d0e3683ec91ea1c[14]      = Id7699f8f89380c315303644fdebacb32 +  ~I56bf74b5890ec67090f499afdc0a9c88 +1;
assign Ia73bc9712b861f909d0e3683ec91ea1c[15]      = Id7699f8f89380c315303644fdebacb32 +  ~Ibaf2f1f8bda2f6b932dc30f8369c0e1f +1;
assign Ia73bc9712b861f909d0e3683ec91ea1c[16]      = Id7699f8f89380c315303644fdebacb32 +  ~Id9364a29fd79b52d0442e18dc0227854 +1;
assign Ia73bc9712b861f909d0e3683ec91ea1c[17]      = Id7699f8f89380c315303644fdebacb32 +  ~Ica3a41ace27f7d94377981079952f4f7 +1;
assign Ia73bc9712b861f909d0e3683ec91ea1c[18]      = Id7699f8f89380c315303644fdebacb32 +  ~Ib57795a63d642a73456324bab41384b6 +1;
assign Ia73bc9712b861f909d0e3683ec91ea1c[19]      = Id7699f8f89380c315303644fdebacb32 +  ~Iabf572c97b48c6a7dcc19e56676e3a82 +1;
assign Ia73bc9712b861f909d0e3683ec91ea1c[20]      = Id7699f8f89380c315303644fdebacb32 +  ~Iefd370d0df1a93639af482f78a1e8706 +1;
assign Ia73bc9712b861f909d0e3683ec91ea1c[21]      = Id7699f8f89380c315303644fdebacb32 +  ~I995d2809ffaf0ecda6a004d01cb9c8c4 +1;
assign Ia73bc9712b861f909d0e3683ec91ea1c[22]      = Id7699f8f89380c315303644fdebacb32 +  ~I4e8ebc46bc068c3f9889d970db131112 +1;
assign I97d2ee9c3120e78ebcda2f0dbb888b49[0]      = Ibf3e1ead3776901898d4b154aeb61267 +  ~I7b561638da1b4a45ff59be81243e4471 +1;
assign I97d2ee9c3120e78ebcda2f0dbb888b49[1]      = Ibf3e1ead3776901898d4b154aeb61267 +  ~If0a3b88a66a816b25f17ced5d0e8f775 +1;
assign I97d2ee9c3120e78ebcda2f0dbb888b49[2]      = Ibf3e1ead3776901898d4b154aeb61267 +  ~I0374ada4fe50717f2158468b7ad205d4 +1;
assign I97d2ee9c3120e78ebcda2f0dbb888b49[3]      = Ibf3e1ead3776901898d4b154aeb61267 +  ~I357137b41bb91e0659b1ac6ead9b5c12 +1;
assign I97d2ee9c3120e78ebcda2f0dbb888b49[4]      = Ibf3e1ead3776901898d4b154aeb61267 +  ~I5d70bc64cf7b3d3ef4180e082e533237 +1;
assign I97d2ee9c3120e78ebcda2f0dbb888b49[5]      = Ibf3e1ead3776901898d4b154aeb61267 +  ~I7d9ad929660cd212387d893266b681da +1;
assign I97d2ee9c3120e78ebcda2f0dbb888b49[6]      = Ibf3e1ead3776901898d4b154aeb61267 +  ~I34be4b353cf75603301372840c2f91c2 +1;
assign I97d2ee9c3120e78ebcda2f0dbb888b49[7]      = Ibf3e1ead3776901898d4b154aeb61267 +  ~I14834fc8e6489775359bcecf5a37ff4d +1;
assign I97d2ee9c3120e78ebcda2f0dbb888b49[8]      = Ibf3e1ead3776901898d4b154aeb61267 +  ~I633a74e4dfa841c9fd13dbb6564c8493 +1;
assign I97d2ee9c3120e78ebcda2f0dbb888b49[9]      = Ibf3e1ead3776901898d4b154aeb61267 +  ~I157bd468200e63385583b9045758d81e +1;
assign I97d2ee9c3120e78ebcda2f0dbb888b49[10]      = Ibf3e1ead3776901898d4b154aeb61267 +  ~I918c46173eebc5b2a95e041cfd91d958 +1;
assign I97d2ee9c3120e78ebcda2f0dbb888b49[11]      = Ibf3e1ead3776901898d4b154aeb61267 +  ~I4f8792c18bd07b23e82bbc44b4ca947f +1;
assign I97d2ee9c3120e78ebcda2f0dbb888b49[12]      = Ibf3e1ead3776901898d4b154aeb61267 +  ~I8d0a1ae4c47edf1f2b99d1175aaa7197 +1;
assign I97d2ee9c3120e78ebcda2f0dbb888b49[13]      = Ibf3e1ead3776901898d4b154aeb61267 +  ~I734e601f5f9d568a44a48834559e04db +1;
assign I97d2ee9c3120e78ebcda2f0dbb888b49[14]      = Ibf3e1ead3776901898d4b154aeb61267 +  ~Ie421da1dc5aaea57c50d0c7d9c5a2717 +1;
assign I97d2ee9c3120e78ebcda2f0dbb888b49[15]      = Ibf3e1ead3776901898d4b154aeb61267 +  ~Ief5cbddfbfb98fce4812a676849b9a98 +1;
assign I97d2ee9c3120e78ebcda2f0dbb888b49[16]      = Ibf3e1ead3776901898d4b154aeb61267 +  ~Id113cab2dd1949d32e3c1c15273185c8 +1;
assign I97d2ee9c3120e78ebcda2f0dbb888b49[17]      = Ibf3e1ead3776901898d4b154aeb61267 +  ~Icfe1a689e33b2b9aa9dba692d6d610b9 +1;
assign I97d2ee9c3120e78ebcda2f0dbb888b49[18]      = Ibf3e1ead3776901898d4b154aeb61267 +  ~Ia4b671f3360f3ce55db0dc0e4d78ddbe +1;
assign I97d2ee9c3120e78ebcda2f0dbb888b49[19]      = Ibf3e1ead3776901898d4b154aeb61267 +  ~I60cbd4369e7ba9b6532f279e5c59084c +1;
assign I97d2ee9c3120e78ebcda2f0dbb888b49[20]      = Ibf3e1ead3776901898d4b154aeb61267 +  ~Ifb6c65a00d9a2c31d8b1119b949828d8 +1;
assign I97d2ee9c3120e78ebcda2f0dbb888b49[21]      = Ibf3e1ead3776901898d4b154aeb61267 +  ~I4a777f0dd62b19dd340ad31517c4e789 +1;
assign I97d2ee9c3120e78ebcda2f0dbb888b49[22]      = Ibf3e1ead3776901898d4b154aeb61267 +  ~Ib75747cb32130d44b338ed8c8af8ca11 +1;
assign I07b2a00225c337eed1e5a350f3361240[0]      = Ie486617fc1d6354c7f347692cdbd894d +  ~Ic7e35cf8d5cd230b94c40714f16e2418 +1;
assign I07b2a00225c337eed1e5a350f3361240[1]      = Ie486617fc1d6354c7f347692cdbd894d +  ~Ic51bb9184dfd103703cd0c6ad6edff4b +1;
assign I07b2a00225c337eed1e5a350f3361240[2]      = Ie486617fc1d6354c7f347692cdbd894d +  ~I103f1449c78c47396d6a54dc1c810934 +1;
assign I07b2a00225c337eed1e5a350f3361240[3]      = Ie486617fc1d6354c7f347692cdbd894d +  ~I56b3a97dc3037f0bb2eed93a9482c813 +1;
assign I07b2a00225c337eed1e5a350f3361240[4]      = Ie486617fc1d6354c7f347692cdbd894d +  ~I51e98035b35a35fdc52f5bab8f19c152 +1;
assign I07b2a00225c337eed1e5a350f3361240[5]      = Ie486617fc1d6354c7f347692cdbd894d +  ~Ia6a7f9beaceb08d81012f0e72171252f +1;
assign I07b2a00225c337eed1e5a350f3361240[6]      = Ie486617fc1d6354c7f347692cdbd894d +  ~I21b062856ced09cb9131c01b5e166f32 +1;
assign I07b2a00225c337eed1e5a350f3361240[7]      = Ie486617fc1d6354c7f347692cdbd894d +  ~I4f1221ce7880729fe584b42ef3afe6b2 +1;
assign I07b2a00225c337eed1e5a350f3361240[8]      = Ie486617fc1d6354c7f347692cdbd894d +  ~Ie7f3f1d6cee7f02ae1b17740ed54c049 +1;
assign I07b2a00225c337eed1e5a350f3361240[9]      = Ie486617fc1d6354c7f347692cdbd894d +  ~Ib196f5bcf9152703dc32c5101076600a +1;
assign I64c650bb94f04521a5a33efa937d9cfc[0]      = I7ba403c6745e7d026282ad704e065702 +  ~Ide9ef5a16d8fe32353c2c2a30e8ee3b0 +1;
assign I64c650bb94f04521a5a33efa937d9cfc[1]      = I7ba403c6745e7d026282ad704e065702 +  ~Iee6f2484a381bd42e441ff072ec582e4 +1;
assign I64c650bb94f04521a5a33efa937d9cfc[2]      = I7ba403c6745e7d026282ad704e065702 +  ~I53121a39de0bcba91a4d0438be2ae958 +1;
assign I64c650bb94f04521a5a33efa937d9cfc[3]      = I7ba403c6745e7d026282ad704e065702 +  ~Iff7950f24f0a6b0073942c37fff49d37 +1;
assign I64c650bb94f04521a5a33efa937d9cfc[4]      = I7ba403c6745e7d026282ad704e065702 +  ~Ide86f019e9573706c25bd8b4552396a8 +1;
assign I64c650bb94f04521a5a33efa937d9cfc[5]      = I7ba403c6745e7d026282ad704e065702 +  ~I2370042234b0e93bb66e44b97fca3e43 +1;
assign I64c650bb94f04521a5a33efa937d9cfc[6]      = I7ba403c6745e7d026282ad704e065702 +  ~If9efe7a1c359ec03014a52870ac13aec +1;
assign I64c650bb94f04521a5a33efa937d9cfc[7]      = I7ba403c6745e7d026282ad704e065702 +  ~I6a6eb62960b616043415406ebfc21346 +1;
assign I64c650bb94f04521a5a33efa937d9cfc[8]      = I7ba403c6745e7d026282ad704e065702 +  ~I06c7728ef64be8311f48d10d766d0c44 +1;
assign I64c650bb94f04521a5a33efa937d9cfc[9]      = I7ba403c6745e7d026282ad704e065702 +  ~I9fe11f6c8147391aa4a5afd1a4e4f731 +1;
assign I34152d4ef2dadfcc943a004e81d175f1[0]      = I93cb3974b8594665b2e7ce5593fde69b +  ~Id50edc56fce48130247fdbc42eeff9ea +1;
assign I34152d4ef2dadfcc943a004e81d175f1[1]      = I93cb3974b8594665b2e7ce5593fde69b +  ~If3e5161254eb9056914c46263b865c10 +1;
assign I34152d4ef2dadfcc943a004e81d175f1[2]      = I93cb3974b8594665b2e7ce5593fde69b +  ~I58703e8b6d04f8c69ac38f5fcfdc4efc +1;
assign I34152d4ef2dadfcc943a004e81d175f1[3]      = I93cb3974b8594665b2e7ce5593fde69b +  ~Ie1f41720e296ced1b74cb325b666d88f +1;
assign I34152d4ef2dadfcc943a004e81d175f1[4]      = I93cb3974b8594665b2e7ce5593fde69b +  ~I5d5701435c96f1078e741921b56e3c65 +1;
assign I34152d4ef2dadfcc943a004e81d175f1[5]      = I93cb3974b8594665b2e7ce5593fde69b +  ~Id96e744d9b10dcddd1ae0115ea57a76a +1;
assign I34152d4ef2dadfcc943a004e81d175f1[6]      = I93cb3974b8594665b2e7ce5593fde69b +  ~I0c0060fe260afa3cdc72f35ffb6938ff +1;
assign I34152d4ef2dadfcc943a004e81d175f1[7]      = I93cb3974b8594665b2e7ce5593fde69b +  ~Iaec1f186cb4a65da21d41e637fc628f7 +1;
assign I34152d4ef2dadfcc943a004e81d175f1[8]      = I93cb3974b8594665b2e7ce5593fde69b +  ~I9c15a6a5c0db11ede80ff6d04c9a56d8 +1;
assign I34152d4ef2dadfcc943a004e81d175f1[9]      = I93cb3974b8594665b2e7ce5593fde69b +  ~I8922487573e02d684a3d71448c3828f5 +1;
assign I745f84653760acc2d83607dcbe1eec73[0]      = Id6a9ab06d58c3a01e1fe04fcf61406fd +  ~I47f17afcd5871fc3ac378316fd3d7ae9 +1;
assign I745f84653760acc2d83607dcbe1eec73[1]      = Id6a9ab06d58c3a01e1fe04fcf61406fd +  ~Ia9642d79bb50567348083b4435c7d66d +1;
assign I745f84653760acc2d83607dcbe1eec73[2]      = Id6a9ab06d58c3a01e1fe04fcf61406fd +  ~I2b2bd845428c49346ef8e94e95b618f8 +1;
assign I745f84653760acc2d83607dcbe1eec73[3]      = Id6a9ab06d58c3a01e1fe04fcf61406fd +  ~Ib730fdb59198f23d1e590f6d6039e96a +1;
assign I745f84653760acc2d83607dcbe1eec73[4]      = Id6a9ab06d58c3a01e1fe04fcf61406fd +  ~I644e83f0a7d432fba38ffb2d99088eca +1;
assign I745f84653760acc2d83607dcbe1eec73[5]      = Id6a9ab06d58c3a01e1fe04fcf61406fd +  ~I97f2b15ce0a74e68d5a4438111adcb0a +1;
assign I745f84653760acc2d83607dcbe1eec73[6]      = Id6a9ab06d58c3a01e1fe04fcf61406fd +  ~I84c88b631bed5311cb6e99e58941149e +1;
assign I745f84653760acc2d83607dcbe1eec73[7]      = Id6a9ab06d58c3a01e1fe04fcf61406fd +  ~I45c5e6710240685bf54b73b0d7a64271 +1;
assign I745f84653760acc2d83607dcbe1eec73[8]      = Id6a9ab06d58c3a01e1fe04fcf61406fd +  ~I5827bc87b5db1801b7db16e1e61515db +1;
assign I745f84653760acc2d83607dcbe1eec73[9]      = Id6a9ab06d58c3a01e1fe04fcf61406fd +  ~I1c85c8f73ef80a6808c6aec0c8eca8ab +1;
assign I9efcf5ce8571b24b590d2d4c8161d49d[0]      = I261bd53528b82128acabd405389c8d60 +  ~Id13c99b7f7500c8195b54627efbc4232 +1;
assign I9efcf5ce8571b24b590d2d4c8161d49d[1]      = I261bd53528b82128acabd405389c8d60 +  ~I4636821315d702a677dc93113872e647 +1;
assign I9efcf5ce8571b24b590d2d4c8161d49d[2]      = I261bd53528b82128acabd405389c8d60 +  ~I9c981b0614a29386ca5e8ebc06a17f15 +1;
assign I9efcf5ce8571b24b590d2d4c8161d49d[3]      = I261bd53528b82128acabd405389c8d60 +  ~I4df3d4dac24877b14e6d361bafc1a800 +1;
assign I9efcf5ce8571b24b590d2d4c8161d49d[4]      = I261bd53528b82128acabd405389c8d60 +  ~I913d818403024510c55b65b56a38dd89 +1;
assign I60a6ef79e3a8244ad32b9833a6ec196b[0]      = If7fa833bf1b1438e7a5bc783ee745252 +  ~I57015930f5b09a6c6b030ed01dad2177 +1;
assign I60a6ef79e3a8244ad32b9833a6ec196b[1]      = If7fa833bf1b1438e7a5bc783ee745252 +  ~Ib54d55a70605119e37e9898b940ff636 +1;
assign I60a6ef79e3a8244ad32b9833a6ec196b[2]      = If7fa833bf1b1438e7a5bc783ee745252 +  ~If7e146da4f3bd255b8457fd6902005f6 +1;
assign I60a6ef79e3a8244ad32b9833a6ec196b[3]      = If7fa833bf1b1438e7a5bc783ee745252 +  ~Ied00d87af99ae55144fdde41ebfc1357 +1;
assign I60a6ef79e3a8244ad32b9833a6ec196b[4]      = If7fa833bf1b1438e7a5bc783ee745252 +  ~I7774313f1ae5a2de98855aad572b3676 +1;
assign I849584bb1c2436f764968afcbb14a61b[0]      = Ibb103853fc21f8f3d466ca16557ccd3e +  ~I679baea452c3c6d04c53baa88edd8eb3 +1;
assign I849584bb1c2436f764968afcbb14a61b[1]      = Ibb103853fc21f8f3d466ca16557ccd3e +  ~If4132b39ddb92aa02d8d0346fb0e6691 +1;
assign I849584bb1c2436f764968afcbb14a61b[2]      = Ibb103853fc21f8f3d466ca16557ccd3e +  ~Iba70e737d52e6812a67c159520e5192f +1;
assign I849584bb1c2436f764968afcbb14a61b[3]      = Ibb103853fc21f8f3d466ca16557ccd3e +  ~Ib9ceb8315f0cd848f861bab677c2c694 +1;
assign I849584bb1c2436f764968afcbb14a61b[4]      = Ibb103853fc21f8f3d466ca16557ccd3e +  ~I7846bc2cc11e08d05f7c853c4920d555 +1;
assign I3ed70f2b460f9278ddeebaf6919b77e8[0]      = I37446eb66ccfd268cb418655b8160fe1 +  ~I0865623d3350645e63fa6e6c9b78ac57 +1;
assign I3ed70f2b460f9278ddeebaf6919b77e8[1]      = I37446eb66ccfd268cb418655b8160fe1 +  ~I0262b30a4efa9f1cfb11d1c3940de9e7 +1;
assign I3ed70f2b460f9278ddeebaf6919b77e8[2]      = I37446eb66ccfd268cb418655b8160fe1 +  ~I7a2e79d42779ad235bca6ce3757cf588 +1;
assign I3ed70f2b460f9278ddeebaf6919b77e8[3]      = I37446eb66ccfd268cb418655b8160fe1 +  ~I09e9a3cd4c12d204f760758e873a177b +1;
assign I3ed70f2b460f9278ddeebaf6919b77e8[4]      = I37446eb66ccfd268cb418655b8160fe1 +  ~I30b0b1d54912c1a41a02a25ab238bb54 +1;
assign I37b4978577c93e476e4a0bc15b9008c9[0]      = Id17f6250f8c7f1d7f75fd27f92698da3 +  ~I49fb0909ddf66fc0073e6400f1a07844 +1;
assign I37b4978577c93e476e4a0bc15b9008c9[1]      = Id17f6250f8c7f1d7f75fd27f92698da3 +  ~I9938397dc94002481984f5b560fadc58 +1;
assign I37b4978577c93e476e4a0bc15b9008c9[2]      = Id17f6250f8c7f1d7f75fd27f92698da3 +  ~I4378d139db4b710e3587aa72df22b70d +1;
assign I37b4978577c93e476e4a0bc15b9008c9[3]      = Id17f6250f8c7f1d7f75fd27f92698da3 +  ~Ifa43d74fa91b7b9884969f575ef9ca8e +1;
assign I37b4978577c93e476e4a0bc15b9008c9[4]      = Id17f6250f8c7f1d7f75fd27f92698da3 +  ~I7c19a79f441ecbb73685db5a505e7479 +1;
assign Ieeaf46eef680115f0d2d108b84b5d3da[0]      = I9957b02e8d0d888e6950eb553d9084d7 +  ~If2af8106efc1f7dd02c074af68278b3d +1;
assign Ieeaf46eef680115f0d2d108b84b5d3da[1]      = I9957b02e8d0d888e6950eb553d9084d7 +  ~I89a3f8d5f760d1a650f85814cbfdc017 +1;
assign Ieeaf46eef680115f0d2d108b84b5d3da[2]      = I9957b02e8d0d888e6950eb553d9084d7 +  ~Ifae345c79662c3df3dff0fe68ad68746 +1;
assign Ieeaf46eef680115f0d2d108b84b5d3da[3]      = I9957b02e8d0d888e6950eb553d9084d7 +  ~I88a61cf72347d695489909d0819332ab +1;
assign Ieeaf46eef680115f0d2d108b84b5d3da[4]      = I9957b02e8d0d888e6950eb553d9084d7 +  ~I9aaa036a6158d11c235bdc8406d79f4c +1;
assign I8b4ff33c17efa28c7eff64664384cffe[0]      = Ic71258b745437bc8463fb4f847c55e27 +  ~Ie8df350430970b5f1229cda772440f85 +1;
assign I8b4ff33c17efa28c7eff64664384cffe[1]      = Ic71258b745437bc8463fb4f847c55e27 +  ~I7d77ac9b64b2e8cae21c6e36947e3ca2 +1;
assign I8b4ff33c17efa28c7eff64664384cffe[2]      = Ic71258b745437bc8463fb4f847c55e27 +  ~Ic1faed76fca5a9ceb7db26c2f43623d9 +1;
assign I8b4ff33c17efa28c7eff64664384cffe[3]      = Ic71258b745437bc8463fb4f847c55e27 +  ~I3ca2b9b77ed8d78a10aff42a07a53b07 +1;
assign I8b4ff33c17efa28c7eff64664384cffe[4]      = Ic71258b745437bc8463fb4f847c55e27 +  ~I1f00849ea055a7893df386aed162a7b6 +1;
assign Ia453e66ce9c1335efac95deebe00c249[0]      = I24bb5c315eacf0f4e8c86f6582389e39 +  ~Iaf8a19fde3de660c3fa925593bebbe0c +1;
assign Ia453e66ce9c1335efac95deebe00c249[1]      = I24bb5c315eacf0f4e8c86f6582389e39 +  ~Icd1da43a4d95230e79dbd35a7ae41066 +1;
assign Ia453e66ce9c1335efac95deebe00c249[2]      = I24bb5c315eacf0f4e8c86f6582389e39 +  ~Ice9079fb6e08d629f8c0c9ce332c8f11 +1;
assign Ia453e66ce9c1335efac95deebe00c249[3]      = I24bb5c315eacf0f4e8c86f6582389e39 +  ~I15fafe2baba4d2f28037023a81ce0a81 +1;
assign Ia453e66ce9c1335efac95deebe00c249[4]      = I24bb5c315eacf0f4e8c86f6582389e39 +  ~If4d5b48882e9e628cf51ad2ac2f38c22 +1;
assign I9c5decf5be3d3e4222559a9c244afc6b[0]      = I607f203694ff76930cfee4103cb73c30 +  ~Id0eef1adba01447c14a6f005782dd9a2 +1;
assign I9c5decf5be3d3e4222559a9c244afc6b[1]      = I607f203694ff76930cfee4103cb73c30 +  ~I1d1a7c5928982c278d068ebd262254da +1;
assign I9c5decf5be3d3e4222559a9c244afc6b[2]      = I607f203694ff76930cfee4103cb73c30 +  ~I6354a0e638340378124e4df7f3d145b8 +1;
assign I9c5decf5be3d3e4222559a9c244afc6b[3]      = I607f203694ff76930cfee4103cb73c30 +  ~I0236c912c6d684bf4862b725be9d5951 +1;
assign I9c5decf5be3d3e4222559a9c244afc6b[4]      = I607f203694ff76930cfee4103cb73c30 +  ~I6f3be51d69b2b64a04e55b8946d5dd56 +1;
assign I9c5decf5be3d3e4222559a9c244afc6b[5]      = I607f203694ff76930cfee4103cb73c30 +  ~Icde3e6dbcf985682041f30903ad95572 +1;
assign I9c5decf5be3d3e4222559a9c244afc6b[6]      = I607f203694ff76930cfee4103cb73c30 +  ~I46ee30b46020d91707689f3468f00e26 +1;
assign I9c5decf5be3d3e4222559a9c244afc6b[7]      = I607f203694ff76930cfee4103cb73c30 +  ~I2605f078c1a9006c93855a9a2b0cf6b9 +1;
assign I9c5decf5be3d3e4222559a9c244afc6b[8]      = I607f203694ff76930cfee4103cb73c30 +  ~I4d226dd2f0bfcdbea6a2e6a6613c1b64 +1;
assign I9c5decf5be3d3e4222559a9c244afc6b[9]      = I607f203694ff76930cfee4103cb73c30 +  ~I5c942076b173cf527e1be2ddb8560e84 +1;
assign I9c5decf5be3d3e4222559a9c244afc6b[10]      = I607f203694ff76930cfee4103cb73c30 +  ~Ic95191bccb18e26c10e56be395ca6b1a +1;
assign I9c5decf5be3d3e4222559a9c244afc6b[11]      = I607f203694ff76930cfee4103cb73c30 +  ~Ia284f974dd8a526f31eb81ed71a06e94 +1;
assign I9c5decf5be3d3e4222559a9c244afc6b[12]      = I607f203694ff76930cfee4103cb73c30 +  ~Icc93450a007cee4c0a42717ed7600528 +1;
assign I9c5decf5be3d3e4222559a9c244afc6b[13]      = I607f203694ff76930cfee4103cb73c30 +  ~I9ec9f389d0489908d497487e44c6edcd +1;
assign I56c4270727a90e00c295c578183a4dce[0]      = Ica8e4c56ebb37e189ca8e6b3daafdb80 +  ~If8a527cc7f06a9963a80a880d225d34c +1;
assign I56c4270727a90e00c295c578183a4dce[1]      = Ica8e4c56ebb37e189ca8e6b3daafdb80 +  ~I39ff4663007dbc89b403f3b08a69bb6c +1;
assign I56c4270727a90e00c295c578183a4dce[2]      = Ica8e4c56ebb37e189ca8e6b3daafdb80 +  ~I9590eb28a81c730b83b92ef7653e71a1 +1;
assign I56c4270727a90e00c295c578183a4dce[3]      = Ica8e4c56ebb37e189ca8e6b3daafdb80 +  ~I2ba1acca919bddcc22a41a28d43a4e3e +1;
assign I56c4270727a90e00c295c578183a4dce[4]      = Ica8e4c56ebb37e189ca8e6b3daafdb80 +  ~I62d8efd4227cb3dc88aa08b6585fafc8 +1;
assign I56c4270727a90e00c295c578183a4dce[5]      = Ica8e4c56ebb37e189ca8e6b3daafdb80 +  ~I749e987266a20840bb8a4b1a2a2fc5b0 +1;
assign I56c4270727a90e00c295c578183a4dce[6]      = Ica8e4c56ebb37e189ca8e6b3daafdb80 +  ~I7607af5d98e8070e3d15cee23cdf877e +1;
assign I56c4270727a90e00c295c578183a4dce[7]      = Ica8e4c56ebb37e189ca8e6b3daafdb80 +  ~I2e11a697d7f17ac30302eadb500de72d +1;
assign I56c4270727a90e00c295c578183a4dce[8]      = Ica8e4c56ebb37e189ca8e6b3daafdb80 +  ~Ia0886ce792e062e22d0c224158cdfb7d +1;
assign I56c4270727a90e00c295c578183a4dce[9]      = Ica8e4c56ebb37e189ca8e6b3daafdb80 +  ~I6b3cd79aa87235ff174c0299b855dd3d +1;
assign I56c4270727a90e00c295c578183a4dce[10]      = Ica8e4c56ebb37e189ca8e6b3daafdb80 +  ~Ie4ae993ddb776bdffec843db0def2f5c +1;
assign I56c4270727a90e00c295c578183a4dce[11]      = Ica8e4c56ebb37e189ca8e6b3daafdb80 +  ~I3ed2da9b53daac0852a06ad1acfad21b +1;
assign I56c4270727a90e00c295c578183a4dce[12]      = Ica8e4c56ebb37e189ca8e6b3daafdb80 +  ~Idefa29d4d4e2a6e9147f84893520096f +1;
assign I56c4270727a90e00c295c578183a4dce[13]      = Ica8e4c56ebb37e189ca8e6b3daafdb80 +  ~Id1fbbe0594dae272856566522633bb3d +1;
assign Ib3e1c6976da60eb724a8d00f19368423[0]      = I7089386c94261e0febf3b4f7dc1aec30 +  ~I8070a3b7d8b1a7ae90c1a2d27aed09aa +1;
assign Ib3e1c6976da60eb724a8d00f19368423[1]      = I7089386c94261e0febf3b4f7dc1aec30 +  ~Ie88285ce2b9c71de02ebd62e8f44ca72 +1;
assign Ib3e1c6976da60eb724a8d00f19368423[2]      = I7089386c94261e0febf3b4f7dc1aec30 +  ~Ica1997c6c569c1d1f45224fbaa4e6b59 +1;
assign Ib3e1c6976da60eb724a8d00f19368423[3]      = I7089386c94261e0febf3b4f7dc1aec30 +  ~Iaf08bcaaeb15bb0c971432f7f8b16d0a +1;
assign Ib3e1c6976da60eb724a8d00f19368423[4]      = I7089386c94261e0febf3b4f7dc1aec30 +  ~Idcb37cfc357cc088c775409fb9225b51 +1;
assign Ib3e1c6976da60eb724a8d00f19368423[5]      = I7089386c94261e0febf3b4f7dc1aec30 +  ~Ic419255414995e7168afb97b051fa64f +1;
assign Ib3e1c6976da60eb724a8d00f19368423[6]      = I7089386c94261e0febf3b4f7dc1aec30 +  ~Iee6da3120d73373627b25ab7c0dedd28 +1;
assign Ib3e1c6976da60eb724a8d00f19368423[7]      = I7089386c94261e0febf3b4f7dc1aec30 +  ~I56fc99a22960232b305d6e683c66fcc7 +1;
assign Ib3e1c6976da60eb724a8d00f19368423[8]      = I7089386c94261e0febf3b4f7dc1aec30 +  ~I0a9a09b0ab43d2a0f1d1d01e13f0333c +1;
assign Ib3e1c6976da60eb724a8d00f19368423[9]      = I7089386c94261e0febf3b4f7dc1aec30 +  ~Ibc73d07e0c97a6fcae791e04106cb082 +1;
assign Ib3e1c6976da60eb724a8d00f19368423[10]      = I7089386c94261e0febf3b4f7dc1aec30 +  ~I224bbdf94ac86c5c376d1db4f4d4e060 +1;
assign Ib3e1c6976da60eb724a8d00f19368423[11]      = I7089386c94261e0febf3b4f7dc1aec30 +  ~I43f2b69c6b427de3095c44d4166b77cd +1;
assign Ib3e1c6976da60eb724a8d00f19368423[12]      = I7089386c94261e0febf3b4f7dc1aec30 +  ~I1e50c90010a3df1a8ce1cff811cc7a0c +1;
assign Ib3e1c6976da60eb724a8d00f19368423[13]      = I7089386c94261e0febf3b4f7dc1aec30 +  ~Ie1817cbf3a80dae435a5571dfbd2f5ad +1;
assign Ib53ea6bc0e3ac45d5a8eecd5dce775d8[0]      = Ia1e4f20f32f7371cb0078d6e80fe8b7e +  ~I0052d562fb3182890c8828e52d437b11 +1;
assign Ib53ea6bc0e3ac45d5a8eecd5dce775d8[1]      = Ia1e4f20f32f7371cb0078d6e80fe8b7e +  ~I1eedecb1d8ff505c75be7787199afada +1;
assign Ib53ea6bc0e3ac45d5a8eecd5dce775d8[2]      = Ia1e4f20f32f7371cb0078d6e80fe8b7e +  ~I7ef544597a185b1de63b4ffc4a1d44c2 +1;
assign Ib53ea6bc0e3ac45d5a8eecd5dce775d8[3]      = Ia1e4f20f32f7371cb0078d6e80fe8b7e +  ~Iadeedf3870f0b1eae98d0f7dbbeff04a +1;
assign Ib53ea6bc0e3ac45d5a8eecd5dce775d8[4]      = Ia1e4f20f32f7371cb0078d6e80fe8b7e +  ~I70ae07db9b44d530be220f06401d3d3d +1;
assign Ib53ea6bc0e3ac45d5a8eecd5dce775d8[5]      = Ia1e4f20f32f7371cb0078d6e80fe8b7e +  ~I7992ea31927b4f0e268462a3b0f18c5d +1;
assign Ib53ea6bc0e3ac45d5a8eecd5dce775d8[6]      = Ia1e4f20f32f7371cb0078d6e80fe8b7e +  ~Iadf927d18644a232ad1f1eba7db82934 +1;
assign Ib53ea6bc0e3ac45d5a8eecd5dce775d8[7]      = Ia1e4f20f32f7371cb0078d6e80fe8b7e +  ~I2a9c673cdd7ded79e09ada38c0f47e6f +1;
assign Ib53ea6bc0e3ac45d5a8eecd5dce775d8[8]      = Ia1e4f20f32f7371cb0078d6e80fe8b7e +  ~Ia86740e870d8063f0266b68ad6d7481d +1;
assign Ib53ea6bc0e3ac45d5a8eecd5dce775d8[9]      = Ia1e4f20f32f7371cb0078d6e80fe8b7e +  ~I6627bcdbaa8afb115123777abd45435b +1;
assign Ib53ea6bc0e3ac45d5a8eecd5dce775d8[10]      = Ia1e4f20f32f7371cb0078d6e80fe8b7e +  ~I96fe3eb633eff6958ac575b997460bb9 +1;
assign Ib53ea6bc0e3ac45d5a8eecd5dce775d8[11]      = Ia1e4f20f32f7371cb0078d6e80fe8b7e +  ~Iefdcb71f2903b11f5cb0b8857f7a1727 +1;
assign Ib53ea6bc0e3ac45d5a8eecd5dce775d8[12]      = Ia1e4f20f32f7371cb0078d6e80fe8b7e +  ~I2eb90278aaa54b9c8212b3b4af7c3617 +1;
assign Ib53ea6bc0e3ac45d5a8eecd5dce775d8[13]      = Ia1e4f20f32f7371cb0078d6e80fe8b7e +  ~I43493f70f0336453d77caf7f27503daa +1;
assign I922408509703b8175883356d89806972[0]      = I790cbca796af58b1726d0a4680cc164f +  ~I26a7fe395eb583258c1ac58aaaa3234a +1;
assign I922408509703b8175883356d89806972[1]      = I790cbca796af58b1726d0a4680cc164f +  ~I21668ff77cf75570cae97f575cbcf644 +1;
assign I922408509703b8175883356d89806972[2]      = I790cbca796af58b1726d0a4680cc164f +  ~Ie48be9e6b6fd63baa104d0a6a4561a1a +1;
assign I922408509703b8175883356d89806972[3]      = I790cbca796af58b1726d0a4680cc164f +  ~I05370777439b01811fe7f750d2f724f4 +1;
assign I922408509703b8175883356d89806972[4]      = I790cbca796af58b1726d0a4680cc164f +  ~Icdcd83341f6b5c404f91ec7e97d0550c +1;
assign I922408509703b8175883356d89806972[5]      = I790cbca796af58b1726d0a4680cc164f +  ~Ibba4e82d1510ddc16eb4ef64893cec02 +1;
assign I922408509703b8175883356d89806972[6]      = I790cbca796af58b1726d0a4680cc164f +  ~Ifb00ae47340bc99669c71da34cccc59e +1;
assign I6cabc68155bc4aef952a07f101ea2802[0]      = I0a93f095f9efb1542116a295c0db9c8b +  ~I75a4cf2948bebc58e12bb039ed273ff2 +1;
assign I6cabc68155bc4aef952a07f101ea2802[1]      = I0a93f095f9efb1542116a295c0db9c8b +  ~I5a9fdec7d7ff99fe33ad6cd8afd9e059 +1;
assign I6cabc68155bc4aef952a07f101ea2802[2]      = I0a93f095f9efb1542116a295c0db9c8b +  ~I47b1695a74e4d27389b97543415dcc67 +1;
assign I6cabc68155bc4aef952a07f101ea2802[3]      = I0a93f095f9efb1542116a295c0db9c8b +  ~Ieb38fa62119a5a77c060d6634e051298 +1;
assign I6cabc68155bc4aef952a07f101ea2802[4]      = I0a93f095f9efb1542116a295c0db9c8b +  ~I3459d98131faef5a5040a03847890b55 +1;
assign I6cabc68155bc4aef952a07f101ea2802[5]      = I0a93f095f9efb1542116a295c0db9c8b +  ~Ie9b9221b2122087cd5f309570b6d31ca +1;
assign I6cabc68155bc4aef952a07f101ea2802[6]      = I0a93f095f9efb1542116a295c0db9c8b +  ~Id4451722e8e2393d627dcd0175dc9903 +1;
assign Ia894c8a3585def468e93aa51039d405c[0]      = I989ba39f188a44475a83e65a4960d2af +  ~Ic10356f9069e3651b9c045c906e63512 +1;
assign Ia894c8a3585def468e93aa51039d405c[1]      = I989ba39f188a44475a83e65a4960d2af +  ~Ic3a431f39c678b7175ed30fde1fa6424 +1;
assign Ia894c8a3585def468e93aa51039d405c[2]      = I989ba39f188a44475a83e65a4960d2af +  ~Ib01cfd833a63500e03333f263805db3d +1;
assign Ia894c8a3585def468e93aa51039d405c[3]      = I989ba39f188a44475a83e65a4960d2af +  ~I0b7b4c0a8503c751229edfe0237cc903 +1;
assign Ia894c8a3585def468e93aa51039d405c[4]      = I989ba39f188a44475a83e65a4960d2af +  ~Iace01234164c8a9f7c98eeb83268745b +1;
assign Ia894c8a3585def468e93aa51039d405c[5]      = I989ba39f188a44475a83e65a4960d2af +  ~Iace8b3b3a4c16763132b5aaa6b24212d +1;
assign Ia894c8a3585def468e93aa51039d405c[6]      = I989ba39f188a44475a83e65a4960d2af +  ~I80a89644e278e96b1cd1c4b7f764dc34 +1;
assign Iaf1c895fc85487f017d3c084e125551c[0]      = I9bcc1d9b3dd258fa7b6042f0185d48cb +  ~Ia92d2276a8a23521ad1b88df7c27bc2e +1;
assign Iaf1c895fc85487f017d3c084e125551c[1]      = I9bcc1d9b3dd258fa7b6042f0185d48cb +  ~I39bbec42c442d1e8c818f46ad9c096a8 +1;
assign Iaf1c895fc85487f017d3c084e125551c[2]      = I9bcc1d9b3dd258fa7b6042f0185d48cb +  ~I88f1b5c12759a5efb2d2ded8483c9ed2 +1;
assign Iaf1c895fc85487f017d3c084e125551c[3]      = I9bcc1d9b3dd258fa7b6042f0185d48cb +  ~Iaf4ae293c576af16f5f43a8b86c1aa3d +1;
assign Iaf1c895fc85487f017d3c084e125551c[4]      = I9bcc1d9b3dd258fa7b6042f0185d48cb +  ~I68b575fcbc5321d4d26a22bcdbb506f6 +1;
assign Iaf1c895fc85487f017d3c084e125551c[5]      = I9bcc1d9b3dd258fa7b6042f0185d48cb +  ~Idf600b93ee1018ecf969ed7944b6bc7b +1;
assign Iaf1c895fc85487f017d3c084e125551c[6]      = I9bcc1d9b3dd258fa7b6042f0185d48cb +  ~I1cd93172cf5996bc870063aa642188a2 +1;
assign I63d67a9bf5a46800216b38df1eb185eb[0]      = I9ba14715d9f33ef45681ad52f5be9593 +  ~I4af080cb4e5cc525db95e5f401019e8c +1;
assign I63d67a9bf5a46800216b38df1eb185eb[1]      = I9ba14715d9f33ef45681ad52f5be9593 +  ~I6fc8044eb226a14ff1a786ddc96d2414 +1;
assign I63d67a9bf5a46800216b38df1eb185eb[2]      = I9ba14715d9f33ef45681ad52f5be9593 +  ~I27fd0073dbcdee599fbe85cf48806efc +1;
assign I63d67a9bf5a46800216b38df1eb185eb[3]      = I9ba14715d9f33ef45681ad52f5be9593 +  ~Iaee6d725a8b2653eeac6d5acb91f8f36 +1;
assign I63d67a9bf5a46800216b38df1eb185eb[4]      = I9ba14715d9f33ef45681ad52f5be9593 +  ~I4afdeba4fc2a12a6cbe3567a519367fc +1;
assign I63d67a9bf5a46800216b38df1eb185eb[5]      = I9ba14715d9f33ef45681ad52f5be9593 +  ~Ib42816335dd8475dcc78662c4c0786c1 +1;
assign I63d67a9bf5a46800216b38df1eb185eb[6]      = I9ba14715d9f33ef45681ad52f5be9593 +  ~I343c9efe71164c01e9c7d599e032864a +1;
assign I63d67a9bf5a46800216b38df1eb185eb[7]      = I9ba14715d9f33ef45681ad52f5be9593 +  ~I108c269ceec4adcff9afeda01101b838 +1;
assign I63d67a9bf5a46800216b38df1eb185eb[8]      = I9ba14715d9f33ef45681ad52f5be9593 +  ~I761983331fb6e3c6c437b3f1660f0b6b +1;
assign I63d67a9bf5a46800216b38df1eb185eb[9]      = I9ba14715d9f33ef45681ad52f5be9593 +  ~I70d32affde22f9dcb2d77430fca39069 +1;
assign I63d67a9bf5a46800216b38df1eb185eb[10]      = I9ba14715d9f33ef45681ad52f5be9593 +  ~Ic08e85346f61da036a15345a13ac12f0 +1;
assign I63d67a9bf5a46800216b38df1eb185eb[11]      = I9ba14715d9f33ef45681ad52f5be9593 +  ~If5dfdadb3868ed5a495007362f7db648 +1;
assign I63d67a9bf5a46800216b38df1eb185eb[12]      = I9ba14715d9f33ef45681ad52f5be9593 +  ~Ia1ee5579358b564de06c08ca418a9bf4 +1;
assign Ic087eef7b3d2a51f34f317a6b9e49144[0]      = I396a897f79b519f4fa02af39d0274f64 +  ~I9bb81dda8102b829441be46460eb8900 +1;
assign Ic087eef7b3d2a51f34f317a6b9e49144[1]      = I396a897f79b519f4fa02af39d0274f64 +  ~I8eef6ca0a61a21882ea28b3d63735228 +1;
assign Ic087eef7b3d2a51f34f317a6b9e49144[2]      = I396a897f79b519f4fa02af39d0274f64 +  ~I438522d92cce6f7010246424746ca255 +1;
assign Ic087eef7b3d2a51f34f317a6b9e49144[3]      = I396a897f79b519f4fa02af39d0274f64 +  ~I92496f68b44a94565af28a2c28d6fbae +1;
assign Ic087eef7b3d2a51f34f317a6b9e49144[4]      = I396a897f79b519f4fa02af39d0274f64 +  ~I66528f43f614f0edb715564eba3c77c1 +1;
assign Ic087eef7b3d2a51f34f317a6b9e49144[5]      = I396a897f79b519f4fa02af39d0274f64 +  ~I8cab9fba615b94fd4bb6934325be8ab8 +1;
assign Ic087eef7b3d2a51f34f317a6b9e49144[6]      = I396a897f79b519f4fa02af39d0274f64 +  ~I92d9fec22d36b1baac8bd78abfc1bbd5 +1;
assign Ic087eef7b3d2a51f34f317a6b9e49144[7]      = I396a897f79b519f4fa02af39d0274f64 +  ~I4eadce87f47df6d8f0e4acd057de5a09 +1;
assign Ic087eef7b3d2a51f34f317a6b9e49144[8]      = I396a897f79b519f4fa02af39d0274f64 +  ~I73203143fe37933c16fff873c1abf512 +1;
assign Ic087eef7b3d2a51f34f317a6b9e49144[9]      = I396a897f79b519f4fa02af39d0274f64 +  ~Ibed2a63af723a7abf96dacf1951e5266 +1;
assign Ic087eef7b3d2a51f34f317a6b9e49144[10]      = I396a897f79b519f4fa02af39d0274f64 +  ~Id667c80003b5541de9f84d3b8709c828 +1;
assign Ic087eef7b3d2a51f34f317a6b9e49144[11]      = I396a897f79b519f4fa02af39d0274f64 +  ~I02cbb4255db2b21ea32140f9e9ddb36b +1;
assign Ic087eef7b3d2a51f34f317a6b9e49144[12]      = I396a897f79b519f4fa02af39d0274f64 +  ~I65354f2069de0c25bbe7cd50fbe892aa +1;
assign I6d360540762be9eab571c0bfe0500f67[0]      = I197c0cd576e16ee2197a28c86397f801 +  ~Ic279867ebf3055980f3d813d5dc8dec6 +1;
assign I6d360540762be9eab571c0bfe0500f67[1]      = I197c0cd576e16ee2197a28c86397f801 +  ~I5c05da8a222ad5effb9815cbf3ec25f3 +1;
assign I6d360540762be9eab571c0bfe0500f67[2]      = I197c0cd576e16ee2197a28c86397f801 +  ~Ib8bf21f32c0e8b9cfa42a53807bfe3a3 +1;
assign I6d360540762be9eab571c0bfe0500f67[3]      = I197c0cd576e16ee2197a28c86397f801 +  ~I7208256bb198bfce1be71390b01bc028 +1;
assign I6d360540762be9eab571c0bfe0500f67[4]      = I197c0cd576e16ee2197a28c86397f801 +  ~I49f2a06ceb3a59773c65b19f54ff362b +1;
assign I6d360540762be9eab571c0bfe0500f67[5]      = I197c0cd576e16ee2197a28c86397f801 +  ~I86e495dc894d2aace15c1aff89798bf7 +1;
assign I6d360540762be9eab571c0bfe0500f67[6]      = I197c0cd576e16ee2197a28c86397f801 +  ~I0d53bb5344cabe5fa5ce3ecf7122a260 +1;
assign I6d360540762be9eab571c0bfe0500f67[7]      = I197c0cd576e16ee2197a28c86397f801 +  ~Ib2f5f5fc77ea8b529f2471c54388f2d1 +1;
assign I6d360540762be9eab571c0bfe0500f67[8]      = I197c0cd576e16ee2197a28c86397f801 +  ~Idcada1bfb3c0d1f2a09aab58a2071a57 +1;
assign I6d360540762be9eab571c0bfe0500f67[9]      = I197c0cd576e16ee2197a28c86397f801 +  ~I814b62120953991f9da055f118967e05 +1;
assign I6d360540762be9eab571c0bfe0500f67[10]      = I197c0cd576e16ee2197a28c86397f801 +  ~I123a212546a8ac394051425db4924812 +1;
assign I6d360540762be9eab571c0bfe0500f67[11]      = I197c0cd576e16ee2197a28c86397f801 +  ~Ie95f1a7e0effcec0aa423dc803056a13 +1;
assign I6d360540762be9eab571c0bfe0500f67[12]      = I197c0cd576e16ee2197a28c86397f801 +  ~I106deaff50b8480eac31ddbae2ec7c61 +1;
assign Ieb702849c7e744c5d04be8f86a00a4fa[0]      = I094a178e55425f27ac1ff6195217396b +  ~I68528be9951f5b8805411711cd11ea59 +1;
assign Ieb702849c7e744c5d04be8f86a00a4fa[1]      = I094a178e55425f27ac1ff6195217396b +  ~I0f034a8f077b0ab231727b6298e366d8 +1;
assign Ieb702849c7e744c5d04be8f86a00a4fa[2]      = I094a178e55425f27ac1ff6195217396b +  ~If9c12f8662333fb54a45cfa1bc5da487 +1;
assign Ieb702849c7e744c5d04be8f86a00a4fa[3]      = I094a178e55425f27ac1ff6195217396b +  ~Ie1681d905517daafcc7584725cd6014c +1;
assign Ieb702849c7e744c5d04be8f86a00a4fa[4]      = I094a178e55425f27ac1ff6195217396b +  ~I2ff3edcdb6158f1e3c9a555aeefc0850 +1;
assign Ieb702849c7e744c5d04be8f86a00a4fa[5]      = I094a178e55425f27ac1ff6195217396b +  ~I43b380be6df7df0d354223d0a0d6d6b6 +1;
assign Ieb702849c7e744c5d04be8f86a00a4fa[6]      = I094a178e55425f27ac1ff6195217396b +  ~I23eb1dc4d1c992f804dd04a2d823c778 +1;
assign Ieb702849c7e744c5d04be8f86a00a4fa[7]      = I094a178e55425f27ac1ff6195217396b +  ~I7f90f96c0260560ad5e6dc7448b2670a +1;
assign Ieb702849c7e744c5d04be8f86a00a4fa[8]      = I094a178e55425f27ac1ff6195217396b +  ~I07b417cdcc99eaea3413f563e26ddc73 +1;
assign Ieb702849c7e744c5d04be8f86a00a4fa[9]      = I094a178e55425f27ac1ff6195217396b +  ~I2f3ab9654e515a54e22e73d6c130ccc3 +1;
assign Ieb702849c7e744c5d04be8f86a00a4fa[10]      = I094a178e55425f27ac1ff6195217396b +  ~Iebdc41368d57498a04fa73e30b10a966 +1;
assign Ieb702849c7e744c5d04be8f86a00a4fa[11]      = I094a178e55425f27ac1ff6195217396b +  ~I5b4305bef5b4350c1d7ae143667afddd +1;
assign Ieb702849c7e744c5d04be8f86a00a4fa[12]      = I094a178e55425f27ac1ff6195217396b +  ~I2795d21d343b83a69146314a2407cfa2 +1;
assign I8519162455bacafeb7f45c170c0b5e7e[0]      = I3177408f7d08b431be99297fb10586e6 +  ~Ic6386d7d8813731d612e24b715740275 +1;
assign I8519162455bacafeb7f45c170c0b5e7e[1]      = I3177408f7d08b431be99297fb10586e6 +  ~I4c366a57920ff090a98a2cb8b9caa00b +1;
assign I8519162455bacafeb7f45c170c0b5e7e[2]      = I3177408f7d08b431be99297fb10586e6 +  ~I14cf5d43fc9864820a8a25efcc5c6d86 +1;
assign I8519162455bacafeb7f45c170c0b5e7e[3]      = I3177408f7d08b431be99297fb10586e6 +  ~I33b99994abbb5ecf8eed4de39033e4f8 +1;
assign I8519162455bacafeb7f45c170c0b5e7e[4]      = I3177408f7d08b431be99297fb10586e6 +  ~I7c3291f0250d13ca94802b0b071a95c6 +1;
assign I8519162455bacafeb7f45c170c0b5e7e[5]      = I3177408f7d08b431be99297fb10586e6 +  ~I2c926fd9d306e9ae13364e07c4b0395b +1;
assign I0d7c184fb7627c9c50a0026ac5052448[0]      = Id4948c876d48bdbf317d32f135e645b4 +  ~Ib23edc35fa5bbfe0415fcf0861a22d9b +1;
assign I0d7c184fb7627c9c50a0026ac5052448[1]      = Id4948c876d48bdbf317d32f135e645b4 +  ~I3e0e682047f7cc36142e668828cbff1e +1;
assign I0d7c184fb7627c9c50a0026ac5052448[2]      = Id4948c876d48bdbf317d32f135e645b4 +  ~I99fb9030e8361e57818c07511479a9b8 +1;
assign I0d7c184fb7627c9c50a0026ac5052448[3]      = Id4948c876d48bdbf317d32f135e645b4 +  ~Ic87c3d7762a18772972552162e1d1a8c +1;
assign I0d7c184fb7627c9c50a0026ac5052448[4]      = Id4948c876d48bdbf317d32f135e645b4 +  ~I7e393e6c1d1bc44daaab120d55f5dd59 +1;
assign I0d7c184fb7627c9c50a0026ac5052448[5]      = Id4948c876d48bdbf317d32f135e645b4 +  ~I448f126fd3932d5065abbe7bb2d92c56 +1;
assign If5cd4834f1cb99b40cd4084fea388070[0]      = Ice5ff01d4fb4583898498651a0ac0171 +  ~Ifc8c6df8904b97674f2970ebc95b523c +1;
assign If5cd4834f1cb99b40cd4084fea388070[1]      = Ice5ff01d4fb4583898498651a0ac0171 +  ~Icd0622a90782b9c451950e7ab0399567 +1;
assign If5cd4834f1cb99b40cd4084fea388070[2]      = Ice5ff01d4fb4583898498651a0ac0171 +  ~I6493b3c087d4685a6b3f98c73dc2ff49 +1;
assign If5cd4834f1cb99b40cd4084fea388070[3]      = Ice5ff01d4fb4583898498651a0ac0171 +  ~I20c2057240417146df144b518b43d052 +1;
assign If5cd4834f1cb99b40cd4084fea388070[4]      = Ice5ff01d4fb4583898498651a0ac0171 +  ~Ied029d0bdea3bf134744c99426fa72dc +1;
assign If5cd4834f1cb99b40cd4084fea388070[5]      = Ice5ff01d4fb4583898498651a0ac0171 +  ~Icb82c9ff4cb58159a1c3115c6fdd5f8c +1;
assign Ia3aa64fb9d2eb1168da1f7e178c05c4e[0]      = I0fb33a5ced3d15622c9aefa188052e24 +  ~Ia3450e134e4086c35acbdee1e6042396 +1;
assign Ia3aa64fb9d2eb1168da1f7e178c05c4e[1]      = I0fb33a5ced3d15622c9aefa188052e24 +  ~I5a0f27df5158309f32f0df31e8ae3ae3 +1;
assign Ia3aa64fb9d2eb1168da1f7e178c05c4e[2]      = I0fb33a5ced3d15622c9aefa188052e24 +  ~I17d9e19854cef197fd3267618617efc3 +1;
assign Ia3aa64fb9d2eb1168da1f7e178c05c4e[3]      = I0fb33a5ced3d15622c9aefa188052e24 +  ~I2993acb61f1abe529f8a60c94a438550 +1;
assign Ia3aa64fb9d2eb1168da1f7e178c05c4e[4]      = I0fb33a5ced3d15622c9aefa188052e24 +  ~Ic8be2c94235fb40f78da33179ce4873a +1;
assign Ia3aa64fb9d2eb1168da1f7e178c05c4e[5]      = I0fb33a5ced3d15622c9aefa188052e24 +  ~Ib3367565e4456da15e7c2315dccdb5e4 +1;
assign I58c319fa3e05e8f7ca440775482ba8fe[0]      = I0074e1c3ca0ff903a9201ac5fe7ca841 +  ~I15a1671def323cd294591564ae6ef8b1 +1;
assign I58c319fa3e05e8f7ca440775482ba8fe[1]      = I0074e1c3ca0ff903a9201ac5fe7ca841 +  ~Ic512effb493a06ece58a2af155135004 +1;
assign I58c319fa3e05e8f7ca440775482ba8fe[2]      = I0074e1c3ca0ff903a9201ac5fe7ca841 +  ~I2c72248cbe49ec0a0febac2437b8a6dc +1;
assign I58c319fa3e05e8f7ca440775482ba8fe[3]      = I0074e1c3ca0ff903a9201ac5fe7ca841 +  ~I964e17c41a134c080e9c43412a514f3f +1;
assign I58c319fa3e05e8f7ca440775482ba8fe[4]      = I0074e1c3ca0ff903a9201ac5fe7ca841 +  ~I94f1724740defe5bb7e40041d0e266a0 +1;
assign I58c319fa3e05e8f7ca440775482ba8fe[5]      = I0074e1c3ca0ff903a9201ac5fe7ca841 +  ~Ic19486b6ab0373b9c0ad8f7597782d8f +1;
assign I58c319fa3e05e8f7ca440775482ba8fe[6]      = I0074e1c3ca0ff903a9201ac5fe7ca841 +  ~I31243de90dc2a1656ca9d5e03bdd78da +1;
assign I58c319fa3e05e8f7ca440775482ba8fe[7]      = I0074e1c3ca0ff903a9201ac5fe7ca841 +  ~I242a30bdc8699d8ff550b25dd53d6c59 +1;
assign I23f3a4487998f2384d9323f9103f7aca[0]      = If65f587e987a51c093e8dd4df532e26c +  ~I9d15f76bb68b214057566cba4b511214 +1;
assign I23f3a4487998f2384d9323f9103f7aca[1]      = If65f587e987a51c093e8dd4df532e26c +  ~I9cc16a00912e7dfc05fb505a9db23cd8 +1;
assign I23f3a4487998f2384d9323f9103f7aca[2]      = If65f587e987a51c093e8dd4df532e26c +  ~Iacf9640cbf486411d6ceb8fe1a2fd5c9 +1;
assign I23f3a4487998f2384d9323f9103f7aca[3]      = If65f587e987a51c093e8dd4df532e26c +  ~I9015033ab0caf3fa41dae4de43f24a82 +1;
assign I23f3a4487998f2384d9323f9103f7aca[4]      = If65f587e987a51c093e8dd4df532e26c +  ~Ia630e59cbce82a570ae3890a6c0221e5 +1;
assign I23f3a4487998f2384d9323f9103f7aca[5]      = If65f587e987a51c093e8dd4df532e26c +  ~I4904ab14b19fa1b6befc218bc7be3842 +1;
assign I23f3a4487998f2384d9323f9103f7aca[6]      = If65f587e987a51c093e8dd4df532e26c +  ~I282d2eb4e74e034694e33273b9cb19d5 +1;
assign I23f3a4487998f2384d9323f9103f7aca[7]      = If65f587e987a51c093e8dd4df532e26c +  ~I3f33901c407a87e10d86c13c83dd52eb +1;
assign I081087845b5c62dc79fd5b9882339572[0]      = I33d7e77d08590f0dfb1867e741dd8b6b +  ~I43f41bf07836cee48069e9890c1de2a0 +1;
assign I081087845b5c62dc79fd5b9882339572[1]      = I33d7e77d08590f0dfb1867e741dd8b6b +  ~Id88480a0a350bb5fcf01ed5fff0bbd4c +1;
assign I081087845b5c62dc79fd5b9882339572[2]      = I33d7e77d08590f0dfb1867e741dd8b6b +  ~I1d9b9ff357667a362f0442f19986f451 +1;
assign I081087845b5c62dc79fd5b9882339572[3]      = I33d7e77d08590f0dfb1867e741dd8b6b +  ~Ice73589836da9028def6efb24a04dbbd +1;
assign I081087845b5c62dc79fd5b9882339572[4]      = I33d7e77d08590f0dfb1867e741dd8b6b +  ~Idb72c046c5996fbbd80b706666ffbd92 +1;
assign I081087845b5c62dc79fd5b9882339572[5]      = I33d7e77d08590f0dfb1867e741dd8b6b +  ~Ie5757e7b1647ab7d43cdbcf98cbb77fc +1;
assign I081087845b5c62dc79fd5b9882339572[6]      = I33d7e77d08590f0dfb1867e741dd8b6b +  ~I6072331f838d82329a07a4ffa340c7b6 +1;
assign I081087845b5c62dc79fd5b9882339572[7]      = I33d7e77d08590f0dfb1867e741dd8b6b +  ~Idf6875955525d80dc660ce956f4a84e7 +1;
assign I8aa441e2ed6f41bca12ddbeaac9f5c3d[0]      = I678c22563e0273403b046df4261f21cf +  ~Ia96955d9c0a8a587e0afab37c8415d8c +1;
assign I8aa441e2ed6f41bca12ddbeaac9f5c3d[1]      = I678c22563e0273403b046df4261f21cf +  ~Ifec374bce7f5507438f550df22d61a01 +1;
assign I8aa441e2ed6f41bca12ddbeaac9f5c3d[2]      = I678c22563e0273403b046df4261f21cf +  ~Ief67e897e57b96e2ec200e82bbc7caeb +1;
assign I8aa441e2ed6f41bca12ddbeaac9f5c3d[3]      = I678c22563e0273403b046df4261f21cf +  ~Ide604e9bbe35cb55892a4602e18b2527 +1;
assign I8aa441e2ed6f41bca12ddbeaac9f5c3d[4]      = I678c22563e0273403b046df4261f21cf +  ~I262f2390e77ec486ccd3a6ed05816e2d +1;
assign I8aa441e2ed6f41bca12ddbeaac9f5c3d[5]      = I678c22563e0273403b046df4261f21cf +  ~I280e20c20c0b4f26278b3de9b2ff84e4 +1;
assign I8aa441e2ed6f41bca12ddbeaac9f5c3d[6]      = I678c22563e0273403b046df4261f21cf +  ~Ib3a0307176d424a4733720416d71069d +1;
assign I8aa441e2ed6f41bca12ddbeaac9f5c3d[7]      = I678c22563e0273403b046df4261f21cf +  ~I76060709de3ea188748849f043c59ac0 +1;
assign I4bc30140a67bbc7b19449fcf946a17aa[0]      = Icca700c12ae2e8155ca6b41e692e8a8c +  ~I8be20605d26d218911e80a883a90d085 +1;
assign I4bc30140a67bbc7b19449fcf946a17aa[1]      = Icca700c12ae2e8155ca6b41e692e8a8c +  ~Ieafa9d74d4a61d28ac4a913db460bf33 +1;
assign I4bc30140a67bbc7b19449fcf946a17aa[2]      = Icca700c12ae2e8155ca6b41e692e8a8c +  ~I6fd1b4395af175eff85b3bfeef4c329b +1;
assign I4bc30140a67bbc7b19449fcf946a17aa[3]      = Icca700c12ae2e8155ca6b41e692e8a8c +  ~I39e6d3fb468aa40ea73535e81556ea65 +1;
assign I4bc30140a67bbc7b19449fcf946a17aa[4]      = Icca700c12ae2e8155ca6b41e692e8a8c +  ~Iae449b74e50e0907feae9e60f2329426 +1;
assign I4bc30140a67bbc7b19449fcf946a17aa[5]      = Icca700c12ae2e8155ca6b41e692e8a8c +  ~Iebf769a6bdaf214c1006c55c608d4eda +1;
assign I4bc30140a67bbc7b19449fcf946a17aa[6]      = Icca700c12ae2e8155ca6b41e692e8a8c +  ~Ia030c08757123aae947f86ab8bfb6d94 +1;
assign I4bc30140a67bbc7b19449fcf946a17aa[7]      = Icca700c12ae2e8155ca6b41e692e8a8c +  ~I8c35c5b343b552c22000e194c517ca12 +1;
assign I4bc30140a67bbc7b19449fcf946a17aa[8]      = Icca700c12ae2e8155ca6b41e692e8a8c +  ~Ibf80bb564263ea85bd886a8617f09bb2 +1;
assign I943f523a14e49f42d9c6ceb3ad1dd841[0]      = I5ed74e81d2497681af5a0ca13fe23088 +  ~Ib8dfd9b8badef282ca00a4f793c3c868 +1;
assign I943f523a14e49f42d9c6ceb3ad1dd841[1]      = I5ed74e81d2497681af5a0ca13fe23088 +  ~I596ad7e132f272cb196b74faa8c75aa4 +1;
assign I943f523a14e49f42d9c6ceb3ad1dd841[2]      = I5ed74e81d2497681af5a0ca13fe23088 +  ~Idc629414f6d0236ce0714cfaae23f065 +1;
assign I943f523a14e49f42d9c6ceb3ad1dd841[3]      = I5ed74e81d2497681af5a0ca13fe23088 +  ~I157fdf8775206858c08682db3039b084 +1;
assign I943f523a14e49f42d9c6ceb3ad1dd841[4]      = I5ed74e81d2497681af5a0ca13fe23088 +  ~Iacbb4daf5ce5c7eb1a2afe30d0cb5382 +1;
assign I943f523a14e49f42d9c6ceb3ad1dd841[5]      = I5ed74e81d2497681af5a0ca13fe23088 +  ~I4e08021c0235fafb60200aab97827a8f +1;
assign I943f523a14e49f42d9c6ceb3ad1dd841[6]      = I5ed74e81d2497681af5a0ca13fe23088 +  ~I730634ea15ac94d241f3ad2d6393a227 +1;
assign I943f523a14e49f42d9c6ceb3ad1dd841[7]      = I5ed74e81d2497681af5a0ca13fe23088 +  ~Iee367c535d9c39f872d2ec043e7e7b33 +1;
assign I943f523a14e49f42d9c6ceb3ad1dd841[8]      = I5ed74e81d2497681af5a0ca13fe23088 +  ~I68bb1f26f878862f288c1f57049cf58b +1;
assign I10ab80965b99680e93ea304f6e261094[0]      = Ic7fa6b8cdfcf7d83d4e101d9c8b7b34f +  ~Ia9b5d9ede006c56a6d83905529c77b7b +1;
assign I10ab80965b99680e93ea304f6e261094[1]      = Ic7fa6b8cdfcf7d83d4e101d9c8b7b34f +  ~I1487170cb1f3370ad45efc801cefc8ab +1;
assign I10ab80965b99680e93ea304f6e261094[2]      = Ic7fa6b8cdfcf7d83d4e101d9c8b7b34f +  ~Id88568dd34fbee42c9cb8cc15ac5c31d +1;
assign I10ab80965b99680e93ea304f6e261094[3]      = Ic7fa6b8cdfcf7d83d4e101d9c8b7b34f +  ~Ia30539545e66c4cfc16828140149180a +1;
assign I10ab80965b99680e93ea304f6e261094[4]      = Ic7fa6b8cdfcf7d83d4e101d9c8b7b34f +  ~Icbfbb37bad6344005dd233b3605a784f +1;
assign I10ab80965b99680e93ea304f6e261094[5]      = Ic7fa6b8cdfcf7d83d4e101d9c8b7b34f +  ~I91a6408a11fab36a8ba3dbd3f895a803 +1;
assign I10ab80965b99680e93ea304f6e261094[6]      = Ic7fa6b8cdfcf7d83d4e101d9c8b7b34f +  ~I47b878f27c30f79a37e97e022307e9e9 +1;
assign I10ab80965b99680e93ea304f6e261094[7]      = Ic7fa6b8cdfcf7d83d4e101d9c8b7b34f +  ~Ie76b0739aec66f8860870e66e87a6445 +1;
assign I10ab80965b99680e93ea304f6e261094[8]      = Ic7fa6b8cdfcf7d83d4e101d9c8b7b34f +  ~I50383e3d7c172eedfa00aa50a9faac4c +1;
assign Ibfef15cf57c5850241c05384f18da5ea[0]      = I26010e26e22d8a2ea831e86fae34a24e +  ~Ifeaa99e03bda8ded058f98387de3d49d +1;
assign Ibfef15cf57c5850241c05384f18da5ea[1]      = I26010e26e22d8a2ea831e86fae34a24e +  ~I4255ac1af4367c321567c4e46b06ab25 +1;
assign Ibfef15cf57c5850241c05384f18da5ea[2]      = I26010e26e22d8a2ea831e86fae34a24e +  ~Ia445bdc7def7d8c1eec31ab892c25c41 +1;
assign Ibfef15cf57c5850241c05384f18da5ea[3]      = I26010e26e22d8a2ea831e86fae34a24e +  ~Ic3b4752136ac08e343933ccc3a4ec47c +1;
assign Ibfef15cf57c5850241c05384f18da5ea[4]      = I26010e26e22d8a2ea831e86fae34a24e +  ~Ica6707efd6d44ba6bbb87c0593a3d828 +1;
assign Ibfef15cf57c5850241c05384f18da5ea[5]      = I26010e26e22d8a2ea831e86fae34a24e +  ~I739267bcc50c54b8a685cb3c6afc5cc1 +1;
assign Ibfef15cf57c5850241c05384f18da5ea[6]      = I26010e26e22d8a2ea831e86fae34a24e +  ~I9160d11439c5140c0109b5190eb82e6b +1;
assign Ibfef15cf57c5850241c05384f18da5ea[7]      = I26010e26e22d8a2ea831e86fae34a24e +  ~I6ff7b86cd7f63f9243646f1be10b2577 +1;
assign Ibfef15cf57c5850241c05384f18da5ea[8]      = I26010e26e22d8a2ea831e86fae34a24e +  ~I165653ab165cfafe2b74cd441331f9e1 +1;
assign I0aa8bcd235f4c4f32c3075d5f39bc20f[0]      = I578efe5c2c504f12c8f2466a7f734215 +  ~I08a8cd6965c23af6650568b654831b20 +1;
assign I0aa8bcd235f4c4f32c3075d5f39bc20f[1]      = I578efe5c2c504f12c8f2466a7f734215 +  ~I9b6a674dbcbfcf65f1ae0deb8fc3566d +1;
assign I0aa8bcd235f4c4f32c3075d5f39bc20f[2]      = I578efe5c2c504f12c8f2466a7f734215 +  ~Ie3a336de822ac7baf8486b1618ef1126 +1;
assign I0aa8bcd235f4c4f32c3075d5f39bc20f[3]      = I578efe5c2c504f12c8f2466a7f734215 +  ~I5fc3c26d6c5aa893dfd5caa0f677233a +1;
assign I0aa8bcd235f4c4f32c3075d5f39bc20f[4]      = I578efe5c2c504f12c8f2466a7f734215 +  ~Ie22b94121b58f17af14c75bfb27f96dd +1;
assign I0aa8bcd235f4c4f32c3075d5f39bc20f[5]      = I578efe5c2c504f12c8f2466a7f734215 +  ~I0d9f8c99194d9d6e187b4ad02fcce8b4 +1;
assign I0aa8bcd235f4c4f32c3075d5f39bc20f[6]      = I578efe5c2c504f12c8f2466a7f734215 +  ~I71e101962e766a4d1484b3235359a4b5 +1;
assign I0aa8bcd235f4c4f32c3075d5f39bc20f[7]      = I578efe5c2c504f12c8f2466a7f734215 +  ~If2539da6722562bbf31786fd0036666a +1;
assign I0aa8bcd235f4c4f32c3075d5f39bc20f[8]      = I578efe5c2c504f12c8f2466a7f734215 +  ~I22c8ccd4a9018ad1c129aa058bf579d8 +1;
assign I0aa8bcd235f4c4f32c3075d5f39bc20f[9]      = I578efe5c2c504f12c8f2466a7f734215 +  ~I83330fef69470d2f5def8e6d7d9c50d2 +1;
assign I0aa8bcd235f4c4f32c3075d5f39bc20f[10]      = I578efe5c2c504f12c8f2466a7f734215 +  ~I0539d598bbe3d50940329a282c801328 +1;
assign I0aa8bcd235f4c4f32c3075d5f39bc20f[11]      = I578efe5c2c504f12c8f2466a7f734215 +  ~I202f88fdc946494d55fc8831c2e8a34c +1;
assign I0aa8bcd235f4c4f32c3075d5f39bc20f[12]      = I578efe5c2c504f12c8f2466a7f734215 +  ~I3ee10f6a7785a236db317515fdd23a2d +1;
assign I0aa8bcd235f4c4f32c3075d5f39bc20f[13]      = I578efe5c2c504f12c8f2466a7f734215 +  ~I453fdf4fbb5af5bd28a20d7643da9eb2 +1;
assign I0aa8bcd235f4c4f32c3075d5f39bc20f[14]      = I578efe5c2c504f12c8f2466a7f734215 +  ~Ic4a6c02880a9aead7353332708e3f388 +1;
assign I0aa8bcd235f4c4f32c3075d5f39bc20f[15]      = I578efe5c2c504f12c8f2466a7f734215 +  ~I7fb3b66cb48521f8715f66bf5642cdb2 +1;
assign Ic5e951c3193081b1880ccf868e740e92[0]      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~I2fd872df07f50688486c0d602cfc5549 +1;
assign Ic5e951c3193081b1880ccf868e740e92[1]      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~Iccefa45795486757515d95e5908b306a +1;
assign Ic5e951c3193081b1880ccf868e740e92[2]      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~Ib1357cb20f471f1670ac2448f964f8eb +1;
assign Ic5e951c3193081b1880ccf868e740e92[3]      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~Iab953a8974a1eb619dc0f074c003b5f9 +1;
assign Ic5e951c3193081b1880ccf868e740e92[4]      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~I6e37582849c2c98fd15ad92d22c222da +1;
assign Ic5e951c3193081b1880ccf868e740e92[5]      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~If004de0cac6e5f7701a1fce48c6936d5 +1;
assign Ic5e951c3193081b1880ccf868e740e92[6]      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~Ic1efa395cc1fd2c5a1d1559fb169a5a0 +1;
assign Ic5e951c3193081b1880ccf868e740e92[7]      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~I8e96c69e7d872be23229353808c34953 +1;
assign Ic5e951c3193081b1880ccf868e740e92[8]      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~Ib6aded6c73a8cc3cb964b0ae895b859e +1;
assign Ic5e951c3193081b1880ccf868e740e92[9]      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~I939368b76d98b43826c68c7f468a5632 +1;
assign Ic5e951c3193081b1880ccf868e740e92[10]      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~I544f6263f16cd5e0b7cf28c511a8f6e3 +1;
assign Ic5e951c3193081b1880ccf868e740e92[11]      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~I484545c4d2c869d79eb17f51e11070a3 +1;
assign Ic5e951c3193081b1880ccf868e740e92[12]      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~I39289e6385a9bc378a9b8dd440249a7f +1;
assign Ic5e951c3193081b1880ccf868e740e92[13]      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~Ie9cce5746a83479a567bbaeac6dbf497 +1;
assign Ic5e951c3193081b1880ccf868e740e92[14]      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~Ic044d7419cc43736d278c2df33b4a3cc +1;
assign Ic5e951c3193081b1880ccf868e740e92[15]      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~I6714551e8885ef5e4490673fe1b2dad1 +1;
assign Ie8edae9436451bc0a4dbdbf531401682[0]      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~Ie9ab3c88ac62369e3d92d110165a94a8 +1;
assign Ie8edae9436451bc0a4dbdbf531401682[1]      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~If38feb4f76f761dce6145731ad235d7f +1;
assign Ie8edae9436451bc0a4dbdbf531401682[2]      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~I6359856a1843d8c8b65dc478bccb3acd +1;
assign Ie8edae9436451bc0a4dbdbf531401682[3]      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~If6f3d91c3c7a43622b9a522492cd83d3 +1;
assign Ie8edae9436451bc0a4dbdbf531401682[4]      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~Id023a6298e65da1f4da3831f5136afc2 +1;
assign Ie8edae9436451bc0a4dbdbf531401682[5]      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~I6b24690f394792edb0d82b3b9e110851 +1;
assign Ie8edae9436451bc0a4dbdbf531401682[6]      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~I5b55c285f7e3e78447fee68532ab9f7f +1;
assign Ie8edae9436451bc0a4dbdbf531401682[7]      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~I32701d9e4b96853c53f0ab651a6a4ba2 +1;
assign Ie8edae9436451bc0a4dbdbf531401682[8]      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~I82f266e5792cdb6e7ebd264e246161f5 +1;
assign Ie8edae9436451bc0a4dbdbf531401682[9]      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~Ibfacfe5b83819afe7fbd4bffa2d6d4e2 +1;
assign Ie8edae9436451bc0a4dbdbf531401682[10]      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~Ib8e68a77ad8b9e7cf415bee17645c3f9 +1;
assign Ie8edae9436451bc0a4dbdbf531401682[11]      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~I644ee0055a55f54ab3544bb532e39c61 +1;
assign Ie8edae9436451bc0a4dbdbf531401682[12]      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~Ic5467e42aa377c6ffd8f70673808774f +1;
assign Ie8edae9436451bc0a4dbdbf531401682[13]      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~Ic57eb4a034247a4c952d8224ea9f2bac +1;
assign Ie8edae9436451bc0a4dbdbf531401682[14]      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~Ia642db613c0ec1ca4e69afde7a14a839 +1;
assign Ie8edae9436451bc0a4dbdbf531401682[15]      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~I432aa7cb844286c442356954f8814260 +1;
assign I84a56b9dce9dfafc97fbdc2ad3b2ae68[0]      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~If520c1cd27f9d4bc52d0d029f693b660 +1;
assign I84a56b9dce9dfafc97fbdc2ad3b2ae68[1]      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~Ie87075ac979410cc11099a356966b8a2 +1;
assign I84a56b9dce9dfafc97fbdc2ad3b2ae68[2]      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~I6fab46b1766878b26b53f352fee98223 +1;
assign I84a56b9dce9dfafc97fbdc2ad3b2ae68[3]      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~Ieaf14683f40374c4531326d228cb43c3 +1;
assign I84a56b9dce9dfafc97fbdc2ad3b2ae68[4]      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~I5149125aaaad943d891df6a3c2be93a0 +1;
assign I84a56b9dce9dfafc97fbdc2ad3b2ae68[5]      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~I770dff588ee1f52f58bea1921cb23383 +1;
assign I84a56b9dce9dfafc97fbdc2ad3b2ae68[6]      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~I8f0a90e761111a613d2488285534a500 +1;
assign I84a56b9dce9dfafc97fbdc2ad3b2ae68[7]      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~I765a8825e42180a6c63f7b33703bb483 +1;
assign I84a56b9dce9dfafc97fbdc2ad3b2ae68[8]      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~I512cc8f6519aa08aee18225b56d47c9f +1;
assign I84a56b9dce9dfafc97fbdc2ad3b2ae68[9]      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~If08370fd0e8af818c6db20f43e74034d +1;
assign I84a56b9dce9dfafc97fbdc2ad3b2ae68[10]      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~I0ff382edfc8051459657ffa3899f5f73 +1;
assign I84a56b9dce9dfafc97fbdc2ad3b2ae68[11]      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~I9d2864024148337277523ef7fa2e1600 +1;
assign I84a56b9dce9dfafc97fbdc2ad3b2ae68[12]      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~I1c85a2d1df6749a194072eb731506bfe +1;
assign I84a56b9dce9dfafc97fbdc2ad3b2ae68[13]      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~I3e3ce8b4ead150a6eae2e5c701c7b598 +1;
assign I84a56b9dce9dfafc97fbdc2ad3b2ae68[14]      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~I45bc13ae0e0554a79c62cd9c6aa8f2a5 +1;
assign I84a56b9dce9dfafc97fbdc2ad3b2ae68[15]      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~I92678f5b52c9c55556ff7f17f0f607b7 +1;
assign I8afac763670df6f56525d3192e04e784[0]      = I0e872d4c07169cac84549178fa144274 +  ~Ib4bdc9069d0c08655f5e87f705943eda +1;
assign I8afac763670df6f56525d3192e04e784[1]      = I0e872d4c07169cac84549178fa144274 +  ~Idbf9094c94c931f16fba468b9dd59a25 +1;
assign I8afac763670df6f56525d3192e04e784[2]      = I0e872d4c07169cac84549178fa144274 +  ~I1c3c4ce44610e04c5eef2fcbc2ea5114 +1;
assign I8afac763670df6f56525d3192e04e784[3]      = I0e872d4c07169cac84549178fa144274 +  ~Ie84be0ae8311d906eff08f7f5b214943 +1;
assign I8afac763670df6f56525d3192e04e784[4]      = I0e872d4c07169cac84549178fa144274 +  ~Ic90b98708faa8c8b75d4bd9a52c292f7 +1;
assign I8afac763670df6f56525d3192e04e784[5]      = I0e872d4c07169cac84549178fa144274 +  ~I8eba6f14f42701d22859fbea94bd1871 +1;
assign I8afac763670df6f56525d3192e04e784[6]      = I0e872d4c07169cac84549178fa144274 +  ~I6d83efa9f988328f487e9232bf2633a2 +1;
assign I8afac763670df6f56525d3192e04e784[7]      = I0e872d4c07169cac84549178fa144274 +  ~Ic23e01562c8a753fd70c343297be288a +1;
assign I8afac763670df6f56525d3192e04e784[8]      = I0e872d4c07169cac84549178fa144274 +  ~I5669856f88f5e2c98f64df696db76414 +1;
assign I8cd574c061a4f1bb0da529d2a892324b[0]      = I6f4ef0f404ae046519b8436171d51e09 +  ~Ic3a608b850709286ea0ad2f67425d9ac +1;
assign I8cd574c061a4f1bb0da529d2a892324b[1]      = I6f4ef0f404ae046519b8436171d51e09 +  ~I5267fa34449e6eebe891017fc32d0749 +1;
assign I8cd574c061a4f1bb0da529d2a892324b[2]      = I6f4ef0f404ae046519b8436171d51e09 +  ~I599d01cfe6e54d8e45d64446c446818d +1;
assign I8cd574c061a4f1bb0da529d2a892324b[3]      = I6f4ef0f404ae046519b8436171d51e09 +  ~I8f94dbafaac589ac9f14b56d4556ff96 +1;
assign I8cd574c061a4f1bb0da529d2a892324b[4]      = I6f4ef0f404ae046519b8436171d51e09 +  ~I754563caea429d3d0e22df5d193b84eb +1;
assign I8cd574c061a4f1bb0da529d2a892324b[5]      = I6f4ef0f404ae046519b8436171d51e09 +  ~If7f373506cac70f8ba1222db135c27e8 +1;
assign I8cd574c061a4f1bb0da529d2a892324b[6]      = I6f4ef0f404ae046519b8436171d51e09 +  ~I69f563e7b7ad483893ac9c4684349769 +1;
assign I8cd574c061a4f1bb0da529d2a892324b[7]      = I6f4ef0f404ae046519b8436171d51e09 +  ~Ia0a02781c674fe5d769206448d475245 +1;
assign I8cd574c061a4f1bb0da529d2a892324b[8]      = I6f4ef0f404ae046519b8436171d51e09 +  ~I1b7a401bc11741e6f011fb9895b5c797 +1;
assign I919a7f8471a46de33447530b4f3b591d[0]      = I4d04e66ad9103a685fbe088b74517452 +  ~Ieb528d666fdb708279184bb59eac25d9 +1;
assign I919a7f8471a46de33447530b4f3b591d[1]      = I4d04e66ad9103a685fbe088b74517452 +  ~Ic3ff7ce12c836bf0693252b9a7a7cfe8 +1;
assign I919a7f8471a46de33447530b4f3b591d[2]      = I4d04e66ad9103a685fbe088b74517452 +  ~I19bba6a58ad3ef959b33701f82761984 +1;
assign I919a7f8471a46de33447530b4f3b591d[3]      = I4d04e66ad9103a685fbe088b74517452 +  ~I8acc93b34974c1e708b0e1591f7b2d3d +1;
assign I919a7f8471a46de33447530b4f3b591d[4]      = I4d04e66ad9103a685fbe088b74517452 +  ~Ib60d4ac0fcadcdfce5a14fb92f58423f +1;
assign I919a7f8471a46de33447530b4f3b591d[5]      = I4d04e66ad9103a685fbe088b74517452 +  ~I039f05d5be891a37e04556f1eae674d2 +1;
assign I919a7f8471a46de33447530b4f3b591d[6]      = I4d04e66ad9103a685fbe088b74517452 +  ~Id0f75e19b94541ed5c5c352d13390d2d +1;
assign I919a7f8471a46de33447530b4f3b591d[7]      = I4d04e66ad9103a685fbe088b74517452 +  ~Ife1190f76c2e251704c2960c23330a48 +1;
assign I919a7f8471a46de33447530b4f3b591d[8]      = I4d04e66ad9103a685fbe088b74517452 +  ~Id3e0c98bff2636e216b4d3a0ffd51054 +1;
assign Ib1f53b5c820345ccdba27ab5be3fa49f[0]      = I988e525020c1e43d238fad41dab4e6ea +  ~If4d3b31b87c0f723241d35ce7e854eba +1;
assign Ib1f53b5c820345ccdba27ab5be3fa49f[1]      = I988e525020c1e43d238fad41dab4e6ea +  ~I72369dedfe36cb22269033cc305b730c +1;
assign Ib1f53b5c820345ccdba27ab5be3fa49f[2]      = I988e525020c1e43d238fad41dab4e6ea +  ~Iec71fe7fcebccf1ae0d10a5d187fcc44 +1;
assign Ib1f53b5c820345ccdba27ab5be3fa49f[3]      = I988e525020c1e43d238fad41dab4e6ea +  ~Ie11da10808c4ca84f399535df6261307 +1;
assign Ib1f53b5c820345ccdba27ab5be3fa49f[4]      = I988e525020c1e43d238fad41dab4e6ea +  ~I280fa9d114e227cd649bf0e55e845651 +1;
assign Ib1f53b5c820345ccdba27ab5be3fa49f[5]      = I988e525020c1e43d238fad41dab4e6ea +  ~I94c4e11670b4233fa072517a8f19c901 +1;
assign Ib1f53b5c820345ccdba27ab5be3fa49f[6]      = I988e525020c1e43d238fad41dab4e6ea +  ~I4dca2dd40a7127ce44f83b430a34c738 +1;
assign Ib1f53b5c820345ccdba27ab5be3fa49f[7]      = I988e525020c1e43d238fad41dab4e6ea +  ~I1a24e98165afa62bd14986911a36fb6e +1;
assign Ib1f53b5c820345ccdba27ab5be3fa49f[8]      = I988e525020c1e43d238fad41dab4e6ea +  ~Ife1164cad7cda4aa9a08d94dfe86add6 +1;
assign I384c493c3195d97eea0a9faaec860f78[0]      = I90d92887cb2526a2956d5e8c9fad760c +  ~I8d8d95ff26f33f69a182b32ccde23905 +1;
assign I384c493c3195d97eea0a9faaec860f78[1]      = I90d92887cb2526a2956d5e8c9fad760c +  ~I2508854bcbab37bd09c9465c377c06aa +1;
assign I384c493c3195d97eea0a9faaec860f78[2]      = I90d92887cb2526a2956d5e8c9fad760c +  ~I140078292f7209eccacd53a8bab18016 +1;
assign I384c493c3195d97eea0a9faaec860f78[3]      = I90d92887cb2526a2956d5e8c9fad760c +  ~I141fb1cbe09f9abe282cffd4de815d25 +1;
assign I384c493c3195d97eea0a9faaec860f78[4]      = I90d92887cb2526a2956d5e8c9fad760c +  ~If79d1d378f7c6fd29fc3335ec5f5c51d +1;
assign I384c493c3195d97eea0a9faaec860f78[5]      = I90d92887cb2526a2956d5e8c9fad760c +  ~I4a41999cea9357a85c73a0af509eeac9 +1;
assign I384c493c3195d97eea0a9faaec860f78[6]      = I90d92887cb2526a2956d5e8c9fad760c +  ~I8e517c401d62dbb10dcc96ab536f6afb +1;
assign I384c493c3195d97eea0a9faaec860f78[7]      = I90d92887cb2526a2956d5e8c9fad760c +  ~I8ad3627f171eadcc960a688ac0afcbc0 +1;
assign I384c493c3195d97eea0a9faaec860f78[8]      = I90d92887cb2526a2956d5e8c9fad760c +  ~I85c4d3d6c8408c6f38741257ed177ca6 +1;
assign I384c493c3195d97eea0a9faaec860f78[9]      = I90d92887cb2526a2956d5e8c9fad760c +  ~Id66c47fd69c175a4393e975a269cf053 +1;
assign I384c493c3195d97eea0a9faaec860f78[10]      = I90d92887cb2526a2956d5e8c9fad760c +  ~I37dca40506d61bdeab1255ed4892ca20 +1;
assign I384c493c3195d97eea0a9faaec860f78[11]      = I90d92887cb2526a2956d5e8c9fad760c +  ~I340c98b886123c541a1b8d9fc8a6d48c +1;
assign Ida1ee79b7a153e40e91549c2180d8425[0]      = I00fe3792cde1eeab36e576fd6634c4fa +  ~I2dc64c3b06588542b027f997437bee63 +1;
assign Ida1ee79b7a153e40e91549c2180d8425[1]      = I00fe3792cde1eeab36e576fd6634c4fa +  ~Id92a37c091100e9df08e24498ecb4022 +1;
assign Ida1ee79b7a153e40e91549c2180d8425[2]      = I00fe3792cde1eeab36e576fd6634c4fa +  ~I74a4b9365391fd20c34588002ad40547 +1;
assign Ida1ee79b7a153e40e91549c2180d8425[3]      = I00fe3792cde1eeab36e576fd6634c4fa +  ~I461195b7ae78743e09ee50486ad6ebe5 +1;
assign Ida1ee79b7a153e40e91549c2180d8425[4]      = I00fe3792cde1eeab36e576fd6634c4fa +  ~I356d747600182675699a2d2634d4c5ce +1;
assign Ida1ee79b7a153e40e91549c2180d8425[5]      = I00fe3792cde1eeab36e576fd6634c4fa +  ~I87d6a5d30c3e4202cf51f33c7a770c51 +1;
assign Ida1ee79b7a153e40e91549c2180d8425[6]      = I00fe3792cde1eeab36e576fd6634c4fa +  ~I960768a84aec9d5b8bc7c1c523024a25 +1;
assign Ida1ee79b7a153e40e91549c2180d8425[7]      = I00fe3792cde1eeab36e576fd6634c4fa +  ~I09b5273bb15d48a7fd78559930fa6d1c +1;
assign Ida1ee79b7a153e40e91549c2180d8425[8]      = I00fe3792cde1eeab36e576fd6634c4fa +  ~I5814a85c45fd0f7be21ed325235fe4b7 +1;
assign Ida1ee79b7a153e40e91549c2180d8425[9]      = I00fe3792cde1eeab36e576fd6634c4fa +  ~Ib06b60cf9933dd8952206c5f3ccced8e +1;
assign Ida1ee79b7a153e40e91549c2180d8425[10]      = I00fe3792cde1eeab36e576fd6634c4fa +  ~I67347c413b5efd8ff9e0d5bc7ab2a047 +1;
assign Ida1ee79b7a153e40e91549c2180d8425[11]      = I00fe3792cde1eeab36e576fd6634c4fa +  ~I72b1bb104bf2843f161448baf7aab44b +1;
assign Ib6bfc051a54fef77204b41e38cdfc6a8[0]      = I6e586c5ac59a28b30c377e51287bf04d +  ~Ib23d889edb5a6d9f27de977d3b1a2616 +1;
assign Ib6bfc051a54fef77204b41e38cdfc6a8[1]      = I6e586c5ac59a28b30c377e51287bf04d +  ~Ifaff9dd032cf96487be819c59b03000a +1;
assign Ib6bfc051a54fef77204b41e38cdfc6a8[2]      = I6e586c5ac59a28b30c377e51287bf04d +  ~I028ce03be0618b816e0ecdf43d4cd6e6 +1;
assign Ib6bfc051a54fef77204b41e38cdfc6a8[3]      = I6e586c5ac59a28b30c377e51287bf04d +  ~I6ae2523095237282533e0b5f1c26b488 +1;
assign Ib6bfc051a54fef77204b41e38cdfc6a8[4]      = I6e586c5ac59a28b30c377e51287bf04d +  ~I5aba6218461e8d571be03a3ef041ebaa +1;
assign Ib6bfc051a54fef77204b41e38cdfc6a8[5]      = I6e586c5ac59a28b30c377e51287bf04d +  ~I6ca8a1fa2c72b1c61d11dc7d1ba5f37b +1;
assign Ib6bfc051a54fef77204b41e38cdfc6a8[6]      = I6e586c5ac59a28b30c377e51287bf04d +  ~I3ec5819176ad4b0895a9118d90ab22b5 +1;
assign Ib6bfc051a54fef77204b41e38cdfc6a8[7]      = I6e586c5ac59a28b30c377e51287bf04d +  ~I49b64469d298012dbb131d879bff38d6 +1;
assign Ib6bfc051a54fef77204b41e38cdfc6a8[8]      = I6e586c5ac59a28b30c377e51287bf04d +  ~I95361d5f524ccb9feb42811af5c482e2 +1;
assign Ib6bfc051a54fef77204b41e38cdfc6a8[9]      = I6e586c5ac59a28b30c377e51287bf04d +  ~I9c4b34b5fb1d59c132bcaeb6258675df +1;
assign Ib6bfc051a54fef77204b41e38cdfc6a8[10]      = I6e586c5ac59a28b30c377e51287bf04d +  ~I613d4b1e3b9e812b785c9cf14fefdfe6 +1;
assign Ib6bfc051a54fef77204b41e38cdfc6a8[11]      = I6e586c5ac59a28b30c377e51287bf04d +  ~I848ed394bd4f0b199d11c0ff458394a7 +1;
assign Ie6d740bc0451311c5f93f4954812613d[0]      = Ib5dc74106d8841d25a793010fdac599a +  ~Ie65a0634454381e24bb3223a333e3ad0 +1;
assign Ie6d740bc0451311c5f93f4954812613d[1]      = Ib5dc74106d8841d25a793010fdac599a +  ~Iad166146f7df5e8068fc6efe4d3e4141 +1;
assign Ie6d740bc0451311c5f93f4954812613d[2]      = Ib5dc74106d8841d25a793010fdac599a +  ~I63e45abd4d27219bddcef06108b72021 +1;
assign Ie6d740bc0451311c5f93f4954812613d[3]      = Ib5dc74106d8841d25a793010fdac599a +  ~Id1bacd13718f7c29c26b63c239d04dd8 +1;
assign Ie6d740bc0451311c5f93f4954812613d[4]      = Ib5dc74106d8841d25a793010fdac599a +  ~Ia3104c69fb4f7abfb5efa3874169a7ad +1;
assign Ie6d740bc0451311c5f93f4954812613d[5]      = Ib5dc74106d8841d25a793010fdac599a +  ~Ie1b7257c99831ec5864f65958ecf14fb +1;
assign Ie6d740bc0451311c5f93f4954812613d[6]      = Ib5dc74106d8841d25a793010fdac599a +  ~I4accbad1b451ed2b622e15ef9ae16d13 +1;
assign Ie6d740bc0451311c5f93f4954812613d[7]      = Ib5dc74106d8841d25a793010fdac599a +  ~I5ce8b2f633011e89356243a1a71edeb6 +1;
assign Ie6d740bc0451311c5f93f4954812613d[8]      = Ib5dc74106d8841d25a793010fdac599a +  ~I3e5139f24e3d082eb31b0e61ea9fa1aa +1;
assign Ie6d740bc0451311c5f93f4954812613d[9]      = Ib5dc74106d8841d25a793010fdac599a +  ~I61cc8a0f49e393721a62a776e4793deb +1;
assign Ie6d740bc0451311c5f93f4954812613d[10]      = Ib5dc74106d8841d25a793010fdac599a +  ~Ie631e40caade823a196370fc3358f042 +1;
assign Ie6d740bc0451311c5f93f4954812613d[11]      = Ib5dc74106d8841d25a793010fdac599a +  ~I4c971e714427664c59c6371e14781bae +1;
assign Ia6ac09257dfd071a132e96619a662f57[0]      = I3eaf142d2734d2d0decef084dc037b50 +  ~I36ca732e811d67cd742d24fd4cae887b +1;
assign Id2e5704c73c707a217875dbf2743e6f3[0]      = I2d171ad83e27a3745d204849a6f46954 +  ~I354fdd241d5d07f0d8380fe8924e0a8c +1;
assign If152a76f9c612e979151b8f51262efc1[0]      = I977f1083f5e4f6f8ac38e2c5aecf1b79 +  ~Id38b705f5d2863a020a475ffffc8afd6 +1;
assign Ifdb6febe29caf3ce300d9cea4954927a[0]      = I9bcd673a4293e14fd20b48fa20492df7 +  ~Id6e5d67e7bb7c4b999459374ea80459a +1;
assign Icfb2b3a2e096f55ba29dd2f9b5761852[0]      = Icb7422ea46b22b9330c123b40fe343fe +  ~I05341013abd4206eb66fcddfd63bfe26 +1;
assign I06c6597547e69bb46e1bede7b7b7f24a[0]      = Ic414cdba230d7ea73972b0eda1ec6b1b +  ~I15da71a21f5842cb65b543d9bc3e267b +1;
assign I325f629c52919e62b3c0075481267744[0]      = Ie4e1e00503dba189b0f871c3c0810d76 +  ~Iccf255fb3422c558465e45226068a16d +1;
assign I56dc657b33a933d2e5d3ac517a9d1fef[0]      = I721c43ab62b42a18c3f5228fc0a73262 +  ~I1c2674b2e6b269ed539827412c5199a5 +1;
assign Ie17d5d171cb71e3748dd0b6c800263ca[0]      = I1f7cb03cf806b247be1cace4d75de942 +  ~I6a3f405bb4a0c4448d9b9d3dd95d036c +1;
assign I9cabb772f5988b877afae0c3b65f340a[0]      = I775cc766b069022bc00220050feee4e4 +  ~Ib528bb7a64cce4f694081d151fa6fa86 +1;
assign Ie29294b754845c1c5602dade95c9e762[0]      = I08b78f774ed494fa7f119977bd92679e +  ~Iaa40bd3abf668a21e0f87c7bda7b3f69 +1;
assign Ibfc5db8e8f393324f06568278da33b4e[0]      = Ic7dc7f94af108ca7c8003a2d07e1e168 +  ~I919d36a7f6ad42c4bbc23222beb73106 +1;
assign I44aace203d154a4d0fc8f10f2cdc5626[0]      = Ibe1327961152cc2d26b3f19476a6e2c9 +  ~I648d2a279dd1f587b1e45eeb35f2fa90 +1;
assign I75526eea62d190615e13ac2731e07074[0]      = I5ba97de444af4e8c9744c3b707502edc +  ~I194a64bef92ecf6714141eaa5d41c9d4 +1;
assign I67bc090d5c81788569b837217febf22d[0]      = I3e4f1314042010b5d7384693b580da7b +  ~Id332e7f482524adeac7f7cdafcf5ca46 +1;
assign I28d725840d5db12ad4940ef965775cc4[0]      = I4a47ce6e21c1a274578397e480c184c9 +  ~I226383d68f89db716cfd8d08b837865a +1;
assign Ia9e617fb96d7ae3706736fafa5dce67c[0]      = Id184731beb200ad6a53ce273b963bb3e +  ~I2bdf5d319ba9089a4da34b108f5c5ae5 +1;
assign Ie033e6fdf59cdfd67ff238b68924dfb5[0]      = I3317f2f6eef9a8ef1fe1ff68b47c5d03 +  ~Ia91800792941ec7cc60415c3f844e4ed +1;
assign I6190c7e2fd99fcb3394fc330e0b08678[0]      = Ia6b9fa10c79e6f3847f89b35afb4cc59 +  ~Id7c507d96098ee7a955af8a48ee5d72a +1;
assign I91f50b160f3a0bc73c84123d977fa4ab[0]      = I91e98b804ef82eea53c5e8eccfec827f +  ~Ie15e4c1bcdb0e18085d4b320ac6a925c +1;
assign Ic05ea9ae53b9396b54c4484a56c7ec79[0]      = I5f1e0d0c6b50f70a6f5584124e095501 +  ~I5485d9edcafc6202f6e5f0969979802f +1;
assign Icf4d6deb47e202e607a07639d064ca55[0]      = Id61fcc605b4b581f5d42024c2610c8b7 +  ~I7fe364f9f537cbef782e7007848a1c10 +1;
assign I85ee05cc8e67b77acbd3ddc7fdfd6bca[0]      = Id64738b7668931553151dbadd5605b71 +  ~I52dcf5bace9cadcf8a895aaa6a8c1da8 +1;
assign I803822a38e626e789a50bade0961edab[0]      = I3bdfb451eb96d256da542864d39024df +  ~I13a9eec6175e695ab8bc4516cf57d6ec +1;
assign If93330fbf9bc863d2837ffc2a0466e70[0]      = Ia740d8ccd8230b28d078b2ea3e58d6ba +  ~Iee73a7c685a4cee03f33d3ef379b1c8a +1;
assign I8ac880ea1c849c493c66a82534400d8c[0]      = I574050722f82569d34bc2cfae1eedaa9 +  ~I740dc91716e3906ad078e2c7cc3c925a +1;
assign I7cf96d4e28b02fd623d8c76161410eb6[0]      = Ic8f7ec6ee09fb9ee2467e3cea30a44a3 +  ~I514d2dc697e9b39ba027c418a6df6cb9 +1;
assign I637636f1d78f96c75bf5c3841419e9fe[0]      = I2b77d922a74fdcef0d57debc789bd539 +  ~I782726e317a2aada9e755bcbc4b0d3fa +1;
assign Icc7d8812ba512a84d2905f1182e69d0a[0]      = Ia1d8127af4944b23475bd7deac91d60e +  ~I11eb26cf0f0b3a334e8f7317bf8d9eb0 +1;
assign Iba60ce25380dc39b44ba505a04453614[0]      = I247abcede9914633c0a33fc402bf58ae +  ~I26cb63ba20245b2c332b09e25c4409aa +1;
assign I9a6a2b184e5122aaa964c2bc818c255d[0]      = I1f413d3e081c6aea012b122fc94f73d5 +  ~Idd7691d31f8d0c09ee988116d574ec59 +1;
assign I4dea7825b6a0eab3aebeb7c4889cdae9[0]      = I1b812fb764d3b48511c0d15a7efaea29 +  ~Iecc02842a2d2b9b9e8187f2d39e62e05 +1;
assign I4809ebf07d855a2e48f92df77ac08b89[0]      = I88882bd8a9f8718411564221ad85b223 +  ~I5551342f1751fc64f32744a46b9649be +1;
assign Ie0a958d83a20d204b3e7a9b4235c4b19[0]      = I232f24e2798488ee66003f3b8cc294c0 +  ~Iff7c29299f005c1cd5a16b64601e727e +1;
assign I8280db7b6ab8c525afd18dc79c0715fb[0]      = I856284e951773518eb6c4232ea7f3d40 +  ~I17a5446e942bcc1dc2c96930e0a87a70 +1;
assign Ifd4e06675d2b57e0064369490c20b8ba[0]      = I82cbeaf5b3e4796b2aaf33dcbd119f4f +  ~I719b67f84e07e90dfd29a8cd5d94cf39 +1;
assign I887915cd3be831277d41e47417ae42e7[0]      = Iaa7791bbc193412e5fe25000ceec23d6 +  ~I2c835dfb3596b8bf057a7cc21122c81f +1;
assign Ic3af54bfe225c905cd146c6ccd3e34e6[0]      = I44bdc0baed3d51ef54ce2728618ad339 +  ~Ib71b3d357c98dcdfae5c777ca3082275 +1;
assign Ida4ab0033193d0b40f4ab5d8b74d7625[0]      = Ib6bc7e75ce750a26113cbb8895c2f024 +  ~I086bf19f620c8a8f6888e775cb1ed7f4 +1;
assign Ic0c2d77062c77982f91941bd99eea68a[0]      = Ib4188380f7e96d5afb99f5045674193d +  ~I802c554d5b04af6b949677819a4966ed +1;
assign I783f9d09de5fce4d69c179fb398a58ae[0]      = I5bba219c5024301e420e9a5acbdc5845 +  ~Iceefb06cb3715e1b41e6f7d89420e5ba +1;
assign I0af2bc8f858473a4b6f9467d5635f2ed[0]      = I1bb52988c9ba03e16b1b69335d3d7e7c +  ~I56948bc48c0220893d68004615a6ebaa +1;
assign Id882b47b85085b9603449499ecfcdb49[0]      = I1b9990aaeae716f66b0f89fb02be0a74 +  ~Iec1368f034655d61354ab5b5e94d7d89 +1;
assign I5b2752f489336c41887046ed4673a717[0]      = Iceec2cf6aba9138648a3340390f39fe9 +  ~I1e43c0aeeb8a2461d208eba24967af30 +1;
assign I75b2328b94afd38404e28c46d7358b22[0]      = Iad7842f3d4672f42c1064c28d4c8ec4e +  ~Ia6eb85b127cf9c1a437611556296b967 +1;
assign I7a642ae71b9f5454a31702d6c3197c79[0]      = Ie5a53cf9343fdcdb5788667c45fadc83 +  ~Ieba89aa901e61218074af53a2484a74b +1;
assign I0f8357de84a9c9e19d35ddd0715b7be4[0]      = I30e06d190906bc9eb6f1c3156c47f9f1 +  ~I8b3b875c6c07bd97ba598a5139156fa4 +1;
assign I76599476765ec5b54c1ed75efddc909d[0]      = Ieaaaced47e22029ad2945eac9cc45e6c +  ~I7b33ddad346077928620344542b9481e +1;
assign I9e277097d3f55ad75b5b0e819d6d3651[0]      = I08dc6f8e837b1f6b80bd3fc742290dab +  ~I11d967a5c5d14c88b5587d4cfed1d05f +1;
assign Ibade670ce04ec07f3b5174fcfc67fabb[0]      = I8eb6a9c907c5909dad6cda98022d70b8 +  ~I27458d76b3ac6520fb379405c6b2956f +1;
assign I19a9636de4b8153208ebef0cfbf811ea[0]      = Ia5067b1b458af82c3c2cd50653099854 +  ~I2525111a2fb5f10d64bbd16e148653b8 +1;
assign Ieb302f84fbd92b0fa4a5747cb1764926[0]      = I198c6753cf12d423c709d1512e66fa9b +  ~I7b7cbcd1c6d2a2eeaaff474536a69eed +1;
assign If88f7bba0fc9ca004e41cf047f6e6410[0]      = Ib600dd8a39fda48d28e1289d44d49a84 +  ~Id2a7f0781d18dccc7c4e0b383b7cddfa +1;
assign I5989aa844d0d73de1a11b8902002efee[0]      = Iabf09191227584c76d7fbc634b706d12 +  ~If8bc141d98ebe1be7fa81cde5c65868e +1;
assign Ia683e321a3334e9668b39f5fea591cd4[0]      = I4869ba08cab90a6dcbc454b0001a7a20 +  ~I8645e1326c66f5efef4b9c923599d1a3 +1;
assign Ic16cfcc11cd03b06afab4b96ab13a350[0]      = If97974406672507f8c9a1c507c4b6951 +  ~I0426ef66185128dd1ef4dbb68dcda585 +1;
assign Icb19ea7dbeb8d826bf85e1e8518e7558[0]      = I4210341f99ac7cb08245137999739114 +  ~Iddd954df5bae9b4240e0512f746669a9 +1;
assign Ie1c0888b2c811ca399501f4669dd8267[0]      = Ic24f4dbd99c8f4d88c8450d4fef762b8 +  ~I29e940970d87e8e09b26ab1b0b8f2286 +1;
assign I65008ba6af7af0ee93fd085692ff4705[0]      = I68dffa1a13eb6ab54615347729c1d6af +  ~I488f6d9676aa85a55d030bf12e8997a7 +1;
assign I0818a864ca9a381fd4b8492410037437[0]      = I10153d5548b184b9ac2cecdba4ec4b1a +  ~I99d761b75ade1fb2e8afbb1a77752609 +1;
assign I11e799346dda7e851c5d48f116216d5a[0]      = I104b7f0512440cffc0fcce25e477f537 +  ~Iac4e3d20178049f9c59abf374752dccc +1;
assign I1bea6ddcb374caef97e35af1eb33d878[0]      = I18b6758319272eebbe76e1eee5ae55b2 +  ~I618d33f26badabfa578908903a613bce +1;
assign Iae87b81938ba6be7fcfb902e35b55ff2[0]      = I780263b10b98f9bb0eaf66c045d8d37c +  ~I822d7973afe090b2764335f1b72dfd0e +1;
assign I2cf76e56c5212c0921ac6725ca41be3c[0]      = I37b772442e55cbcd44ba892a0608d662 +  ~I12c1035353e553b3b6a13bb174ce6020 +1;
assign I21cf97f59f8387bdd451934e800a501d[0]      = I0ac256a6659ff5c6673fd110a8bf578f +  ~Ia6d61947d36fc128c689808c82db80f6 +1;
assign I9c91a8ca3a41b5df249ad6e0cd9b6601[0]      = If134e1d27e736005e5a390e7a2ea1f4b +  ~Ie9b042f686381739b9ff219041f1e0ce +1;
assign I02e4ad55fc6e12cd60370ae782bbd36b[0]      = I7b37b8f908cd82683832536e02faab0d +  ~I0c4268c01aed70ce4fc71531bf4bb862 +1;
assign I5192b23d7d4742e17ffcf58679d96734[0]      = I08b4bf60c9c7e7229bd1952cc88bc7b3 +  ~Ia34e42f8de91fa4861b0c6cac5dcfc29 +1;
assign I0aaea02d5fbc4cfe6478060df6a92441[0]      = I267d637eb63fef9f4723f7978fad88f0 +  ~Ib7c5850b4f7cc77be2048d114a2128d9 +1;
assign I64476c4b13b6612ab90845870c8fcec6[0]      = I4fb56a70e5ffa71f58f715da36368e04 +  ~I32bb50faa2b246b2d3b462a79be597c5 +1;
assign I46cb13c147e8087f9f93618f946d0f75[0]      = I5e9e2acb258baf96ac4b525bba54a462 +  ~Idc6d40a49f05c5422758cee50f787eb1 +1;
assign Ida1dc39acb508dea4487357625f65a62[0]      = Ic40f61443a4d8f87769067fc39381cb3 +  ~Ide1d7dc22a4b271ef764df14ac22366a +1;
assign Ief0a83a4d2ab6337a9a842850ed9c8d2[0]      = Ieb36710c9a3726f33407436d62639c8d +  ~I7ace6778ac86b3e05939a3fcc716136f +1;
assign Iabc0481ca8b87650597db2ab82d9526a[0]      = Ic804af393da2e4b9c8ef25d4a3b4e8d5 +  ~I044e01e8d2df46e03f00a0af2beb0bf5 +1;
assign I273daf63e8da53e5e9b99de802715b44[0]      = I52e4c446693c29a42bb3b665f72d382d +  ~I45a7ddcda2662e36b7617dfe64514346 +1;
assign I9bec797aec01899ccab507296d7f4d53[0]      = Idbf02cf10add496d30fa44bbb18458c6 +  ~Idada779a1ac7b844867571d77054b657 +1;
assign Id769ce05d2596a106b4e750d272b6d86[0]      = Ida095585ad26e215f1c1bf989912da89 +  ~Ieeba01b18a244ab8c0ac263c138fabcc +1;
assign Ifcd0ef96ba3a7a7ef8ab4f64c5671f80[0]      = I19f1ffa05c7c9a0df5e7014044024c7b +  ~Ie4c9797a955778694dd8615219cb51e7 +1;
assign I2789f24264b92b82f7e9f34a5ccaa489[0]      = I4d68a2fe778fa93faac38b138138291f +  ~I28a5ed4c239e64c76bb6e566b50cfd23 +1;
assign Ic9f02e5a9bad9928c784d38980f709ff[0]      = I54393ada6f76ac82c31f2668e228e29d +  ~I79a705ee1e414fe4a5fb14e9b3ce9597 +1;
assign I5729f3c3121489f404f8964abb3e842a[0]      = If5b9ef84f09680f3593250b13a852c1c +  ~I04f90a907f10a7fa1ae3591b48094d5c +1;
assign If076d265cc6b8f7baf4059ea5fa7525d[0]      = Ibb759bc4179e5b7aa759d850c7cfa467 +  ~I31d25b1b49e65216e90b39aa27acd6be +1;
assign I7acc5316ae2768ce90598a82ad196eca[0]      = I05e8b5f8b83f07b609b5ebf272bb2229 +  ~I1f6540c5f037d861dee2c0091cba01ec +1;
assign Idc81e8df0b1b36ee2885c180c992a8db[0]      = If6ac15373ec1146d38e7aeb71c3ece64 +  ~I9632bb500b7faaaaeb649d74c21cbe8c +1;
assign I2f587d7d70873b05956908ded54c36f9[0]      = I2ab3675e1eede757af80716ba980a4e6 +  ~Idd0217a35c3adc8abc7bb581a5df7a2d +1;
assign I7f013f76d9fcc1b14984188e7af2ec0d[0]      = I388c271687ab31b57421ad57192273ed +  ~Ic05b46168884322644db4e331d37d759 +1;
assign Ica4903599938b7e1996702a51a7e9ec8[0]      = I6121679cec8caa51dc5ff0d1a61f9821 +  ~I53c88dc237bb2cd02d50fd7f0a168a48 +1;
assign I53484a61ff8b4273d872779c33b292d5[0]      = Ia0649b990bf5716cfab230127cd5d47f +  ~I7450d4ab3ef0227e93a02bfd620d047b +1;
assign Iae00c13f4457b91d9a252b5b2aa67780[0]      = I867a0626ca22108b16267d95c0aadf4f +  ~I2b16e5b4e279bb29c3c675b72083e5fe +1;
assign I208b29bdae3040b547e8e40ffdc96d34[0]      = I1af54bcb73d7c6b93e55450871207976 +  ~I70c92e8ada46476d15ef4b3c620d2601 +1;
assign Ic6378ae3bd73ac1ddfb25e7d7882c671[0]      = I91883553543d0425e9c6dd726dce3d27 +  ~Ib193b07804d6d5f111b06bda487bfa5f +1;
assign I81f95de60a5dd186e51f9f4bf0b624da[0]      = Ie95405659701278e3f87bf1f823a037b +  ~I885433b0ab16c6d87abe45af13c9e529 +1;
assign Ic05bdf0bf00ca3ba90c6ee7728b2d49b[0]      = Ia42392e2104b50c0908aad82738a5ee7 +  ~I198c055930cb89d0390c336eda8fed4f +1;
assign Ic74ef5ce41d9db0920015b60cd80dada[0]      = I68ad63230a51b9b9e3daffb307ea970d +  ~I688a2c72e69b217d2673e8da75146a83 +1;
assign If54ee451267f16296945fca60801b6da[0]      = I7a052d63944ccf42e598efe3a95b88f8 +  ~I3b6fde4ed14cd68af1468ae1d4cc1a22 +1;
assign I22af03550c9ffd5ee75db6b34f444612[0]      = I2b3c6d69f79c8d51e4d1614c62c44fcc +  ~I5d3df1e7563630311f56143ee6d97a8e +1;
assign I76d5529e20b89a706595f65abe004da2[0]      = Ifcef0e92f50e3920bf1208af5d64c632 +  ~I90a7ea789d3bf7f9126c786474a56da0 +1;
assign Iebca060c7873173db59d0e1a244a5f62[0]      = I111340a19625901a3c1b95fd0bd1570e +  ~I5029424c9d9fe923eeb858b1e62cd758 +1;
assign I39ebf0c6f66596aeb1c56eaf50bc6b55[0]      = I11aec4fa85c30f6fe1fd9fa72542ef6c +  ~I1e805c70d50c2765b4a03ad2982dc421 +1;
assign I685db637ba885fcd9a37a9457b56c827[0]      = I80cc333c181c16a96b7bd6501c27c2b3 +  ~Iba58175a7fd5c5da650222193caff0b3 +1;
assign If659617a922c1800e53f789111d7f946[0]      = Idc6354325a6280ae9890da33c06c33ec +  ~I7401a0501ba69c5559fbf00c77e58dc5 +1;
assign I3cde77dbb4b236619f7d00d6212d8f46[0]      = Ibb04cf82acc4ac16599ad3ddb0c2ada2 +  ~Idd9f7ea657ea9cdcb45a7e4b573b9d50 +1;
assign Ic1f7f01098e573cdab8482bd3f0dfe0c[0]      = I3ed096dfd8a14f4acb4d53a70cf8aceb +  ~I53f275395dd6be17961a5edc3e8da7f2 +1;
assign Ic229657d83879de9bd470c1739254faa[0]      = I0fa07f95e96326cb0599c0c3f76e2b48 +  ~Icab010d78cd66b02e089c74f04bf4e75 +1;
assign I3e69a3b20cf7ac74e77887b37fc3a5d7[0]      = I87d98fbc97d9a78c2e7d6a6280e7a49a +  ~I376a48b7e0195a5aacc76a0ad8bd14b2 +1;
assign Ief74f9042bd0058f17af181156b58456[0]      = Ib7ddc4dca877f7cf5697a02c3d1915ba +  ~I241622b0367dde514f96ece55c8c3964 +1;
assign Ide1209ba9c80b0f69b0f17a1320b7a33[0]      = I3612ef280891f6017fad205d0484bde7 +  ~If94a1abfb972f63629d07e64dc23863c +1;
assign Ib8c08ba5cf3c7bd8233532cc8ecb4825[0]      = I561547649aeb5b4c3f10d9506db1f3cf +  ~I07b9b1f4fa01b16cc69356057d3b6154 +1;
assign I812e31439ca7c94df3d6bf578b60beaf[0]      = I84cc76c0079b86da7b994844c3ccb875 +  ~I2288a6ad3b748b716249f4adc42d52c4 +1;
assign Ie93978ee93511b6ed29aad9aed8ee903[0]      = Iec013c508d0c6401d7eb856e7eb60446 +  ~I022df337bcc05ac5648b8ae2e42f3a76 +1;
assign If0c12a1750d279b90738aacac5b35e04[0]      = Ifd8979aac6b6b24aa560b46b18240e92 +  ~I60d9a7f95fb8623753002ecaf9a4efcc +1;
assign I0501ec6e9230839738818ae2b19a5b65[0]      = If12394e78dc913b01890b56650856a44 +  ~I23a74ea5e7174d95e6d16a5e85ac236b +1;
assign I9e9c3529814bb741e0e425dba9ba0abf[0]      = I94d18aa10695f3f22b23246884b72822 +  ~Ie697d28d757df82b3901564bda43251c +1;
assign I3898f311fc81d9bbcda50e18e7f978e1[0]      = Ic90b38835dd7e760dd54067b196f8470 +  ~I8572aedc94f7243ce5eacb332c81eae2 +1;
assign I4bf59374718f169f17fea6adb9d9c7e1[0]      = If3691ea51f6efe9b165a31964854d2fe +  ~I6734123aaf6320da75638b212812732f +1;
assign Ide127cda229e55eca7ef703c0d794e6e[0]      = Ic2ce582555add38a14f5006d3c87eb15 +  ~I7f6dc6f0f403c58f9aaaa70c2383a666 +1;
assign I482955b75319360d2646b1f712acdbde[0]      = I58cc950ee2cbe56b7c5a619be3792511 +  ~I66391978843c39b6acbdb4847a01050a +1;
assign I158984c3dfe52e5107e4aa64548c1ab5[0]      = I0d8e329ec5873db96df1ec309445a096 +  ~I4f756e4125c8af5c412944b273e01cb0 +1;
assign Ibdfb487053f2567b45db76d12e9eb75a[0]      = I106325488e2ecfdba1cf9e5201e6bc8c +  ~Id2c9f7ac95de07148c54803f69347f56 +1;
assign I1fc2b706279a62a29d90f261f211c3a9[0]      = Iff73a0085541a511d3912b64686a82c5 +  ~I5061e13a179d27e1ba5f89ce8ee0fd4a +1;
assign I988227c12ad87b2ced8fd8fd89eb138d[0]      = Icdab59de68f2870504598c9ea18f1d2c +  ~I0f7c32fc1548fb49b8041f55c157498a +1;
assign Id537c7ec3b2e195d892f7fb1a63dcf46[0]      = I75604d727e82c977741f90113719183a +  ~I89ffab735ee30423c82e079ed98216c5 +1;
assign I92a93c16158990f624973e9cc487fc00[0]      = I6f50c4d0d2639857b2dcca300c2d7b04 +  ~I9494921d8487ee0b314f75cf0380fd2f +1;
assign Iab0879a7d17f0fbf2c2ed147e41d3f32[0]      = I5cd013a2be2e761c10c6a957632517de +  ~If2b3e7d1541cbd8ffc2b4cfc3ad13a57 +1;
assign I762ebc964e606e803121e347086668e4[0]      = Iafeedddd02428bd2610c576e68d4ae25 +  ~Idf3d79da44f2d686f5bd43c3c1427430 +1;
assign I032010a0a18eaf23274cdff5c99442bc[0]      = I912d6325e34180e0f668f0f024e63581 +  ~If8125ad3c9e7f0a2b84106064d320996 +1;
assign I24956c032de466de716b6ab57dd8a265[0]      = Id1e05294dfd02df499ad0c08bb5c191b +  ~Ic9018b88fa91fb638bbab0613795ae13 +1;
assign If816e24bfd42448c3c0fb03b6e9e9404[0]      = Id3bb9b100ee4302473b49ac14615e9b0 +  ~Iad4ea0196eb32f9a152c9e6fe5059e46 +1;
assign I0903046199323180f148f13aedaa0ab3[0]      = Ief32db1cfc443119b6202b0cc7bf70a2 +  ~Ia8ff29ed728e7f2ae4213f00328b495d +1;
assign I25ec8dfa866fe300e67a01944f893bf6[0]      = Iad7dbe9909b5eed3261adf92d3813acc +  ~I70717726200ec02929f679ef05496455 +1;
assign I77ac8c7c5ea03d948931590d57c8d649[0]      = Ie7daf0789c35caaadbba06cafabd2b70 +  ~Iaf1e4c7dae6ad89567836877c08f57d2 +1;
assign Ief5d16bc74276d3aec10a56fe8234b8a[0]      = I2bd1f9b75d9ab94af9ddceb7528935e8 +  ~Icd09aa81e9b43528af73e23b2f0f80cb +1;
assign I6bec62410ca887855fafaa4be4c09d72[0]      = Ic3d9f5c6677758810e4865779ec303e3 +  ~I6ebb2b94f0f80425f8401ae823d92a1d +1;
assign I290223476b30aa41df98af3016119109[0]      = I00af04882a25e2832d913a67d4d86d7b +  ~I4a2c3204a6a9936d4a215b46c0ffd045 +1;
assign I07e3ae59ec05fa46d6ca3398a42e287c[0]      = Ic9db631df0a1a9108c10c3e0eca7bf15 +  ~Ib02c0694762c4815448b2c8d3df767c2 +1;
assign I7b019b5e5991ad8497a048367d83341f[0]      = I749f9ed1fb2dddd40ebc28f638e02935 +  ~I98cee6efbbe565d3a4de16703189782f +1;
assign I80f8ed713e4b0281f94804a0b66fadcf[0]      = Ia45b2a24df24bd5e3c95885c8928686c +  ~Ibf981c01a9d44cbea3c6d8ead92bc2ab +1;
assign I8cd2472defb068d6e3af7070c97c25ef[0]      = I7427464fde340780aba7f9847b4ad564 +  ~I864c33e8ea204d20a9baef4584f22d4e +1;
assign I3689f559a9636f9dd4558e99424d6c80[0]      = I33fd1ae225e2b881b2b41e0358675e22 +  ~I6ad3228e0e2e1f19648d73e83ba5a229 +1;
assign I77c454b260ff3c291b59ac8679966ab1[0]      = I2e21a35d1cf560936fd19b944a208b6b +  ~Ie099210a99a4899c53baf39559592690 +1;
assign Iddb9b8c346479631362bfc4aa039b746[0]      = I249522a3d42cc75d7a6b9ede1222ee76 +  ~Ieeec71d9df4613555fade2ced7b3baf1 +1;
assign I3db9cdf51e4437b6e979f8c1a0be96df[0]      = I68b4c43d9f40ae4bfd70d2983594392c +  ~I4931884e3544af182bcda9061091a42d +1;
assign I2a2352cab4f2edc64f156ef7b5e5595b[0]      = I63145e0fec15c7e7c0de105f348bfd31 +  ~Ib3fb10da528d450251764a9b9ede0dba +1;
assign Iee3314c9bfca7066dcbb138d5f46d1f8[0]      = I8af625de86c04016c3424d116fddab5b +  ~Icdc9e676957b2223d60c413331fa982f +1;
assign I4883185d078ac45e5eb2d6dbcd2c875b[0]      = I54c9c10527f83b4ee4e1e22f1e4044ed +  ~I381f6051282c062ccf53866830344cd4 +1;
assign Ie6242ba25d061a37a41d7ca41370e919[0]      = I972559e47c7f83bd9000ca1cfc14d8e0 +  ~Icfc21935c007fbbceb2a67ebe1a68a0b +1;
assign I99d9fb1f21a8aba32da690b3bbb786df[0]      = Ib97a7f941eb7ce2a867503a04ff86a67 +  ~I120d597a80158374726e064fb0f099fb +1;
assign I1328d62797b528de9c98372d828d4af0[0]      = I5979b55f607c71017537f2b48b40cbea +  ~I2520aa556aadf851f58f0b1820498730 +1;
assign Id71c488586e019260c79018420d61673[0]      = I6a56760b621f238843b091279c69897f +  ~I6203f49a08107f7185ebadeecf2c16b0 +1;
assign I6f2d4122c89e56e6640df3cec76c3c48[0]      = Icec45bf76c241d37c9a50a5cd092da9d +  ~Ia706fb593b63cebbee0321c154cb859b +1;
assign I37d02ddb7b52ae3495a3a182a3d4708a[0]      = I2f6d3f61f2890e584d3063a09587e99b +  ~Ia4b5f2b07556629673fc6576bc49a5dc +1;
assign I30b006cb2cf34c967066041123ac3698[0]      = I7c396ea2e959d84fd9a6964617cb29c6 +  ~Ic532c6b85b156f821e0742f47239a65c +1;

// Ie4894ca167b08880bfc35862f18575eb Ied2b5c0139cec8ad2873829dc1117d50 I05531b19bb846b18c09f979eeb429ad3 I92354deea988f3beb25bfba90735c6ac valid Ied2b5c0139cec8ad2873829dc1117d50 I6d3acefe6d7dfb94a5d66dcaa1bbbb76
       assign tmp_bit[0]  =   (I748f85f6680918a2e992df339b4b6558[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[1]  =   (Ib0f57837099e3fdf1b908d78bcda4a43[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[2]  =   (If75e99660e3997f53f7b903bc366f47f[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[3]  =   (I3253481bee7dbfc0f3eac94c3252ee4e[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[4]  =   (Ia80693da8182ee2c3708b6ec21d397d2[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[5]  =   (I7fa3f2648baacebf9e4b59c179601fa6[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[6]  =   (Id7699f8f89380c315303644fdebacb32[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[7]  =   (Ibf3e1ead3776901898d4b154aeb61267[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[8]  =   (Ie486617fc1d6354c7f347692cdbd894d[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[9]  =   (I7ba403c6745e7d026282ad704e065702[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[10]  =   (I93cb3974b8594665b2e7ce5593fde69b[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[11]  =   (Id6a9ab06d58c3a01e1fe04fcf61406fd[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[12]  =   (I261bd53528b82128acabd405389c8d60[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[13]  =   (If7fa833bf1b1438e7a5bc783ee745252[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[14]  =   (Ibb103853fc21f8f3d466ca16557ccd3e[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[15]  =   (I37446eb66ccfd268cb418655b8160fe1[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[16]  =   (Id17f6250f8c7f1d7f75fd27f92698da3[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[17]  =   (I9957b02e8d0d888e6950eb553d9084d7[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[18]  =   (Ic71258b745437bc8463fb4f847c55e27[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[19]  =   (I24bb5c315eacf0f4e8c86f6582389e39[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[20]  =   (I607f203694ff76930cfee4103cb73c30[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[21]  =   (Ica8e4c56ebb37e189ca8e6b3daafdb80[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[22]  =   (I7089386c94261e0febf3b4f7dc1aec30[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[23]  =   (Ia1e4f20f32f7371cb0078d6e80fe8b7e[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[24]  =   (I790cbca796af58b1726d0a4680cc164f[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[25]  =   (I0a93f095f9efb1542116a295c0db9c8b[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[26]  =   (I989ba39f188a44475a83e65a4960d2af[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[27]  =   (I9bcc1d9b3dd258fa7b6042f0185d48cb[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[28]  =   (I9ba14715d9f33ef45681ad52f5be9593[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[29]  =   (I396a897f79b519f4fa02af39d0274f64[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[30]  =   (I197c0cd576e16ee2197a28c86397f801[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[31]  =   (I094a178e55425f27ac1ff6195217396b[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[32]  =   (I3177408f7d08b431be99297fb10586e6[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[33]  =   (Id4948c876d48bdbf317d32f135e645b4[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[34]  =   (Ice5ff01d4fb4583898498651a0ac0171[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[35]  =   (I0fb33a5ced3d15622c9aefa188052e24[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[36]  =   (I0074e1c3ca0ff903a9201ac5fe7ca841[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[37]  =   (If65f587e987a51c093e8dd4df532e26c[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[38]  =   (I33d7e77d08590f0dfb1867e741dd8b6b[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[39]  =   (I678c22563e0273403b046df4261f21cf[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[40]  =   (Icca700c12ae2e8155ca6b41e692e8a8c[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[41]  =   (I5ed74e81d2497681af5a0ca13fe23088[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[42]  =   (Ic7fa6b8cdfcf7d83d4e101d9c8b7b34f[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[43]  =   (I26010e26e22d8a2ea831e86fae34a24e[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[44]  =   (I578efe5c2c504f12c8f2466a7f734215[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[45]  =   (Ida86d05f907d23ff9fed06927c2ec9d9[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[46]  =   (I9d9f8c7a23d9750ec44e706bf763df76[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[47]  =   (I0b41b002a32b8e9e2fe68e819f228fb7[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[48]  =   (I0e872d4c07169cac84549178fa144274[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[49]  =   (I6f4ef0f404ae046519b8436171d51e09[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[50]  =   (I4d04e66ad9103a685fbe088b74517452[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[51]  =   (I988e525020c1e43d238fad41dab4e6ea[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[52]  =   (I90d92887cb2526a2956d5e8c9fad760c[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[53]  =   (I00fe3792cde1eeab36e576fd6634c4fa[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[54]  =   (I6e586c5ac59a28b30c377e51287bf04d[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[55]  =   (Ib5dc74106d8841d25a793010fdac599a[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[56]  =   (I3eaf142d2734d2d0decef084dc037b50[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[57]  =   (I2d171ad83e27a3745d204849a6f46954[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[58]  =   (I977f1083f5e4f6f8ac38e2c5aecf1b79[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[59]  =   (I9bcd673a4293e14fd20b48fa20492df7[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[60]  =   (Icb7422ea46b22b9330c123b40fe343fe[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[61]  =   (Ic414cdba230d7ea73972b0eda1ec6b1b[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[62]  =   (Ie4e1e00503dba189b0f871c3c0810d76[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[63]  =   (I721c43ab62b42a18c3f5228fc0a73262[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[64]  =   (I1f7cb03cf806b247be1cace4d75de942[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[65]  =   (I775cc766b069022bc00220050feee4e4[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[66]  =   (I08b78f774ed494fa7f119977bd92679e[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[67]  =   (Ic7dc7f94af108ca7c8003a2d07e1e168[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[68]  =   (Ibe1327961152cc2d26b3f19476a6e2c9[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[69]  =   (I5ba97de444af4e8c9744c3b707502edc[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[70]  =   (I3e4f1314042010b5d7384693b580da7b[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[71]  =   (I4a47ce6e21c1a274578397e480c184c9[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[72]  =   (Id184731beb200ad6a53ce273b963bb3e[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[73]  =   (I3317f2f6eef9a8ef1fe1ff68b47c5d03[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[74]  =   (Ia6b9fa10c79e6f3847f89b35afb4cc59[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[75]  =   (I91e98b804ef82eea53c5e8eccfec827f[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[76]  =   (I5f1e0d0c6b50f70a6f5584124e095501[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[77]  =   (Id61fcc605b4b581f5d42024c2610c8b7[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[78]  =   (Id64738b7668931553151dbadd5605b71[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[79]  =   (I3bdfb451eb96d256da542864d39024df[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[80]  =   (Ia740d8ccd8230b28d078b2ea3e58d6ba[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[81]  =   (I574050722f82569d34bc2cfae1eedaa9[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[82]  =   (Ic8f7ec6ee09fb9ee2467e3cea30a44a3[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[83]  =   (I2b77d922a74fdcef0d57debc789bd539[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[84]  =   (Ia1d8127af4944b23475bd7deac91d60e[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[85]  =   (I247abcede9914633c0a33fc402bf58ae[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[86]  =   (I1f413d3e081c6aea012b122fc94f73d5[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[87]  =   (I1b812fb764d3b48511c0d15a7efaea29[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[88]  =   (I88882bd8a9f8718411564221ad85b223[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[89]  =   (I232f24e2798488ee66003f3b8cc294c0[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[90]  =   (I856284e951773518eb6c4232ea7f3d40[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[91]  =   (I82cbeaf5b3e4796b2aaf33dcbd119f4f[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[92]  =   (Iaa7791bbc193412e5fe25000ceec23d6[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[93]  =   (I44bdc0baed3d51ef54ce2728618ad339[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[94]  =   (Ib6bc7e75ce750a26113cbb8895c2f024[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[95]  =   (Ib4188380f7e96d5afb99f5045674193d[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[96]  =   (I5bba219c5024301e420e9a5acbdc5845[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[97]  =   (I1bb52988c9ba03e16b1b69335d3d7e7c[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[98]  =   (I1b9990aaeae716f66b0f89fb02be0a74[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[99]  =   (Iceec2cf6aba9138648a3340390f39fe9[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[100]  =   (Iad7842f3d4672f42c1064c28d4c8ec4e[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[101]  =   (Ie5a53cf9343fdcdb5788667c45fadc83[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[102]  =   (I30e06d190906bc9eb6f1c3156c47f9f1[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[103]  =   (Ieaaaced47e22029ad2945eac9cc45e6c[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[104]  =   (I08dc6f8e837b1f6b80bd3fc742290dab[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[105]  =   (I8eb6a9c907c5909dad6cda98022d70b8[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[106]  =   (Ia5067b1b458af82c3c2cd50653099854[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[107]  =   (I198c6753cf12d423c709d1512e66fa9b[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[108]  =   (Ib600dd8a39fda48d28e1289d44d49a84[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[109]  =   (Iabf09191227584c76d7fbc634b706d12[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[110]  =   (I4869ba08cab90a6dcbc454b0001a7a20[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[111]  =   (If97974406672507f8c9a1c507c4b6951[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[112]  =   (I4210341f99ac7cb08245137999739114[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[113]  =   (Ic24f4dbd99c8f4d88c8450d4fef762b8[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[114]  =   (I68dffa1a13eb6ab54615347729c1d6af[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[115]  =   (I10153d5548b184b9ac2cecdba4ec4b1a[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[116]  =   (I104b7f0512440cffc0fcce25e477f537[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[117]  =   (I18b6758319272eebbe76e1eee5ae55b2[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[118]  =   (I780263b10b98f9bb0eaf66c045d8d37c[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[119]  =   (I37b772442e55cbcd44ba892a0608d662[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[120]  =   (I0ac256a6659ff5c6673fd110a8bf578f[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[121]  =   (If134e1d27e736005e5a390e7a2ea1f4b[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[122]  =   (I7b37b8f908cd82683832536e02faab0d[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[123]  =   (I08b4bf60c9c7e7229bd1952cc88bc7b3[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[124]  =   (I267d637eb63fef9f4723f7978fad88f0[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[125]  =   (I4fb56a70e5ffa71f58f715da36368e04[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[126]  =   (I5e9e2acb258baf96ac4b525bba54a462[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[127]  =   (Ic40f61443a4d8f87769067fc39381cb3[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[128]  =   (Ieb36710c9a3726f33407436d62639c8d[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[129]  =   (Ic804af393da2e4b9c8ef25d4a3b4e8d5[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[130]  =   (I52e4c446693c29a42bb3b665f72d382d[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[131]  =   (Idbf02cf10add496d30fa44bbb18458c6[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[132]  =   (Ida095585ad26e215f1c1bf989912da89[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[133]  =   (I19f1ffa05c7c9a0df5e7014044024c7b[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[134]  =   (I4d68a2fe778fa93faac38b138138291f[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[135]  =   (I54393ada6f76ac82c31f2668e228e29d[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[136]  =   (If5b9ef84f09680f3593250b13a852c1c[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[137]  =   (Ibb759bc4179e5b7aa759d850c7cfa467[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[138]  =   (I05e8b5f8b83f07b609b5ebf272bb2229[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[139]  =   (If6ac15373ec1146d38e7aeb71c3ece64[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[140]  =   (I2ab3675e1eede757af80716ba980a4e6[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[141]  =   (I388c271687ab31b57421ad57192273ed[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[142]  =   (I6121679cec8caa51dc5ff0d1a61f9821[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[143]  =   (Ia0649b990bf5716cfab230127cd5d47f[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[144]  =   (I867a0626ca22108b16267d95c0aadf4f[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[145]  =   (I1af54bcb73d7c6b93e55450871207976[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[146]  =   (I91883553543d0425e9c6dd726dce3d27[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[147]  =   (Ie95405659701278e3f87bf1f823a037b[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[148]  =   (Ia42392e2104b50c0908aad82738a5ee7[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[149]  =   (I68ad63230a51b9b9e3daffb307ea970d[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[150]  =   (I7a052d63944ccf42e598efe3a95b88f8[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[151]  =   (I2b3c6d69f79c8d51e4d1614c62c44fcc[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[152]  =   (Ifcef0e92f50e3920bf1208af5d64c632[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[153]  =   (I111340a19625901a3c1b95fd0bd1570e[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[154]  =   (I11aec4fa85c30f6fe1fd9fa72542ef6c[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[155]  =   (I80cc333c181c16a96b7bd6501c27c2b3[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[156]  =   (Idc6354325a6280ae9890da33c06c33ec[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[157]  =   (Ibb04cf82acc4ac16599ad3ddb0c2ada2[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[158]  =   (I3ed096dfd8a14f4acb4d53a70cf8aceb[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[159]  =   (I0fa07f95e96326cb0599c0c3f76e2b48[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[160]  =   (I87d98fbc97d9a78c2e7d6a6280e7a49a[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[161]  =   (Ib7ddc4dca877f7cf5697a02c3d1915ba[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[162]  =   (I3612ef280891f6017fad205d0484bde7[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[163]  =   (I561547649aeb5b4c3f10d9506db1f3cf[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[164]  =   (I84cc76c0079b86da7b994844c3ccb875[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[165]  =   (Iec013c508d0c6401d7eb856e7eb60446[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[166]  =   (Ifd8979aac6b6b24aa560b46b18240e92[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[167]  =   (If12394e78dc913b01890b56650856a44[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[168]  =   (I94d18aa10695f3f22b23246884b72822[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[169]  =   (Ic90b38835dd7e760dd54067b196f8470[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[170]  =   (If3691ea51f6efe9b165a31964854d2fe[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[171]  =   (Ic2ce582555add38a14f5006d3c87eb15[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[172]  =   (I58cc950ee2cbe56b7c5a619be3792511[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[173]  =   (I0d8e329ec5873db96df1ec309445a096[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[174]  =   (I106325488e2ecfdba1cf9e5201e6bc8c[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[175]  =   (Iff73a0085541a511d3912b64686a82c5[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[176]  =   (Icdab59de68f2870504598c9ea18f1d2c[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[177]  =   (I75604d727e82c977741f90113719183a[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[178]  =   (I6f50c4d0d2639857b2dcca300c2d7b04[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[179]  =   (I5cd013a2be2e761c10c6a957632517de[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[180]  =   (Iafeedddd02428bd2610c576e68d4ae25[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[181]  =   (I912d6325e34180e0f668f0f024e63581[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[182]  =   (Id1e05294dfd02df499ad0c08bb5c191b[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[183]  =   (Id3bb9b100ee4302473b49ac14615e9b0[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[184]  =   (Ief32db1cfc443119b6202b0cc7bf70a2[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[185]  =   (Iad7dbe9909b5eed3261adf92d3813acc[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[186]  =   (Ie7daf0789c35caaadbba06cafabd2b70[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[187]  =   (I2bd1f9b75d9ab94af9ddceb7528935e8[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[188]  =   (Ic3d9f5c6677758810e4865779ec303e3[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[189]  =   (I00af04882a25e2832d913a67d4d86d7b[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[190]  =   (Ic9db631df0a1a9108c10c3e0eca7bf15[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[191]  =   (I749f9ed1fb2dddd40ebc28f638e02935[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[192]  =   (Ia45b2a24df24bd5e3c95885c8928686c[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[193]  =   (I7427464fde340780aba7f9847b4ad564[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[194]  =   (I33fd1ae225e2b881b2b41e0358675e22[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[195]  =   (I2e21a35d1cf560936fd19b944a208b6b[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[196]  =   (I249522a3d42cc75d7a6b9ede1222ee76[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[197]  =   (I68b4c43d9f40ae4bfd70d2983594392c[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[198]  =   (I63145e0fec15c7e7c0de105f348bfd31[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[199]  =   (I8af625de86c04016c3424d116fddab5b[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[200]  =   (I54c9c10527f83b4ee4e1e22f1e4044ed[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[201]  =   (I972559e47c7f83bd9000ca1cfc14d8e0[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[202]  =   (Ib97a7f941eb7ce2a867503a04ff86a67[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[203]  =   (I5979b55f607c71017537f2b48b40cbea[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[204]  =   (I6a56760b621f238843b091279c69897f[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[205]  =   (Icec45bf76c241d37c9a50a5cd092da9d[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[206]  =   (I2f6d3f61f2890e584d3063a09587e99b[SIGN_MAX_SUM_WDTH_LONG]);
       assign tmp_bit[207]  =   (I7c396ea2e959d84fd9a6964617cb29c6[SIGN_MAX_SUM_WDTH_LONG]);







always_comb begin
            I43864225be03ea8e9379eb28dfa6c599 = I29b4fdd4c13c96461c76660df767ea73(I95878a848ec38c4f334bc1915576e6d6[0]);
            I31cb0c699cffcd2fedfbed0e1b86490e = I29b4fdd4c13c96461c76660df767ea73(I95878a848ec38c4f334bc1915576e6d6[1]);
            Ibed5004d869a01005768ba694c2234d6 = I29b4fdd4c13c96461c76660df767ea73(I95878a848ec38c4f334bc1915576e6d6[2]);
            Ia4b2db3d48f946b0bfd0be0e32d7518d = I29b4fdd4c13c96461c76660df767ea73(I95878a848ec38c4f334bc1915576e6d6[3]);
            I4d908bbe633c193cd9fc93dd33c60bd2 = I29b4fdd4c13c96461c76660df767ea73(I95878a848ec38c4f334bc1915576e6d6[4]);
            Ib14733d3585dbf7f196cfc068e9508f0 = I29b4fdd4c13c96461c76660df767ea73(I95878a848ec38c4f334bc1915576e6d6[5]);
            Idfcf7f3240d92bfc87d44833bc00ff9d = I29b4fdd4c13c96461c76660df767ea73(I95878a848ec38c4f334bc1915576e6d6[6]);
            I1cff7306aaf303bb3342ea3d72048908 = I29b4fdd4c13c96461c76660df767ea73(I95878a848ec38c4f334bc1915576e6d6[7]);
            I26bdcc44692db066911c8d5b0a1aae0c = I29b4fdd4c13c96461c76660df767ea73(I95878a848ec38c4f334bc1915576e6d6[8]);
            Id144785da9b171f1e2d0e9182d693e31 = I29b4fdd4c13c96461c76660df767ea73(I95878a848ec38c4f334bc1915576e6d6[9]);
            I6b7a8ba12de5b44817ec99faebe54617 = I29b4fdd4c13c96461c76660df767ea73(I95878a848ec38c4f334bc1915576e6d6[10]);
            I4a403449a9ba75243369032e1cca1a0d = I29b4fdd4c13c96461c76660df767ea73(I95878a848ec38c4f334bc1915576e6d6[11]);
            If85d9a95c1c02ce2da1dc3486b53eb81 = I29b4fdd4c13c96461c76660df767ea73(I95878a848ec38c4f334bc1915576e6d6[12]);
            I8e470b68bf35c647af42b6e46201e570 = I29b4fdd4c13c96461c76660df767ea73(I95878a848ec38c4f334bc1915576e6d6[13]);
            I484ec87270fcc959a486ebce40a9a03c = I29b4fdd4c13c96461c76660df767ea73(I95878a848ec38c4f334bc1915576e6d6[14]);
            I079932780612fbce79cbe9b58bb6c2b5 = I29b4fdd4c13c96461c76660df767ea73(I95878a848ec38c4f334bc1915576e6d6[15]);
            Ibb157b97546cb19fa7c1c0a7c79b1d38 = I29b4fdd4c13c96461c76660df767ea73(I95878a848ec38c4f334bc1915576e6d6[16]);
            I45cb51c25c426c296f97a5d23a08c063 = I29b4fdd4c13c96461c76660df767ea73(I95878a848ec38c4f334bc1915576e6d6[17]);
            Iff1d4b06901796098f91e87a3c30f7a5 = I29b4fdd4c13c96461c76660df767ea73(I95878a848ec38c4f334bc1915576e6d6[18]);
            I16db9cab1981451a02dab21e2ca221b4 = I29b4fdd4c13c96461c76660df767ea73(I95878a848ec38c4f334bc1915576e6d6[19]);
            I72756ea6a4997bc4afd4bfde1dfb2d26 = I29b4fdd4c13c96461c76660df767ea73(I95878a848ec38c4f334bc1915576e6d6[20]);
            I2882ae2eb6d79a5b96d1ed937dcfd8bf = I29b4fdd4c13c96461c76660df767ea73(I95878a848ec38c4f334bc1915576e6d6[21]);
            I1a632a3e06ad738d5865acc77e204f48 = I29b4fdd4c13c96461c76660df767ea73(I3eb1902edf9266038f39c281d134c26c[0]);
            I4d4ec5540257040d10182ed478a71918 = I29b4fdd4c13c96461c76660df767ea73(I3eb1902edf9266038f39c281d134c26c[1]);
            I8da7e01f56dc9a70eb6b3f110dc005c2 = I29b4fdd4c13c96461c76660df767ea73(I3eb1902edf9266038f39c281d134c26c[2]);
            Icc5d7bcbd7fcdb5092e6d8e18f6de6ec = I29b4fdd4c13c96461c76660df767ea73(I3eb1902edf9266038f39c281d134c26c[3]);
            I83cec264bd378f1dc23f87e439e7310e = I29b4fdd4c13c96461c76660df767ea73(I3eb1902edf9266038f39c281d134c26c[4]);
            Ied7e494fb288f78d110ed06662f1926a = I29b4fdd4c13c96461c76660df767ea73(I3eb1902edf9266038f39c281d134c26c[5]);
            Idd5b362dab4f93bba0c39af78c4c5981 = I29b4fdd4c13c96461c76660df767ea73(I3eb1902edf9266038f39c281d134c26c[6]);
            Id033e7adfcfb0420cc592a1fb6c297b6 = I29b4fdd4c13c96461c76660df767ea73(I3eb1902edf9266038f39c281d134c26c[7]);
            Iaee91a5e94c3f174682f72a1ebfd0021 = I29b4fdd4c13c96461c76660df767ea73(I3eb1902edf9266038f39c281d134c26c[8]);
            I0cd8a6e719305ee3fbe8228081993957 = I29b4fdd4c13c96461c76660df767ea73(I3eb1902edf9266038f39c281d134c26c[9]);
            I9b8cfdb69b76453a3ac687a1e098417f = I29b4fdd4c13c96461c76660df767ea73(I3eb1902edf9266038f39c281d134c26c[10]);
            Ic2159627df2efa5e677fa6f4498bdd31 = I29b4fdd4c13c96461c76660df767ea73(I3eb1902edf9266038f39c281d134c26c[11]);
            I59fba74472ded0a985cb237104ac127f = I29b4fdd4c13c96461c76660df767ea73(I3eb1902edf9266038f39c281d134c26c[12]);
            Ia526539cc0f844b802d412b7a17cb6a6 = I29b4fdd4c13c96461c76660df767ea73(I3eb1902edf9266038f39c281d134c26c[13]);
            I5d80b7c7d102d2c2bfa73a68c73376be = I29b4fdd4c13c96461c76660df767ea73(I3eb1902edf9266038f39c281d134c26c[14]);
            Ia92defa0ca87c7c30fbe901da40a575e = I29b4fdd4c13c96461c76660df767ea73(I3eb1902edf9266038f39c281d134c26c[15]);
            I8fb1602dcdcd2912ea8aec42e2b7848f = I29b4fdd4c13c96461c76660df767ea73(I3eb1902edf9266038f39c281d134c26c[16]);
            I0cedca0e2c589104d6f3318505910594 = I29b4fdd4c13c96461c76660df767ea73(I3eb1902edf9266038f39c281d134c26c[17]);
            I54c260db5c1b2c76527c8fc1cee229fe = I29b4fdd4c13c96461c76660df767ea73(I3eb1902edf9266038f39c281d134c26c[18]);
            I3d700e050cb7f22b0e381f3c72a20124 = I29b4fdd4c13c96461c76660df767ea73(I3eb1902edf9266038f39c281d134c26c[19]);
            I63c0c8bef1dea4e499a16ce01e781951 = I29b4fdd4c13c96461c76660df767ea73(I3eb1902edf9266038f39c281d134c26c[20]);
            Ia8abcb8cf8d9ecc17c27ff015aa0b71f = I29b4fdd4c13c96461c76660df767ea73(I3eb1902edf9266038f39c281d134c26c[21]);
            I3f59174b3764a0b0741462024be9fb92 = I29b4fdd4c13c96461c76660df767ea73(Ie791b43e8d5c9d1669743ea4d6e3139c[0]);
            If0c2d002c315b21e11ae776bb48c9338 = I29b4fdd4c13c96461c76660df767ea73(Ie791b43e8d5c9d1669743ea4d6e3139c[1]);
            I18e548b082364c75686f2b7ad2ef46ab = I29b4fdd4c13c96461c76660df767ea73(Ie791b43e8d5c9d1669743ea4d6e3139c[2]);
            I5e0d6b44474a226ab2ce916a6d46072a = I29b4fdd4c13c96461c76660df767ea73(Ie791b43e8d5c9d1669743ea4d6e3139c[3]);
            I0c53d8d6a5b92960e29fc31cf456c23b = I29b4fdd4c13c96461c76660df767ea73(Ie791b43e8d5c9d1669743ea4d6e3139c[4]);
            Ib16c6096ce80e2f15a5ccea145e28510 = I29b4fdd4c13c96461c76660df767ea73(Ie791b43e8d5c9d1669743ea4d6e3139c[5]);
            I0e7ca2d6470b9bfc6a1ca6143b468507 = I29b4fdd4c13c96461c76660df767ea73(Ie791b43e8d5c9d1669743ea4d6e3139c[6]);
            I4ba05e74c2f63e2f4c59268775d549aa = I29b4fdd4c13c96461c76660df767ea73(Ie791b43e8d5c9d1669743ea4d6e3139c[7]);
            Iaed26e1c4a2578d16b111d15d31339d2 = I29b4fdd4c13c96461c76660df767ea73(Ie791b43e8d5c9d1669743ea4d6e3139c[8]);
            Ic566fe27ccaf2220101cbc49fc187a6b = I29b4fdd4c13c96461c76660df767ea73(Ie791b43e8d5c9d1669743ea4d6e3139c[9]);
            Ibf9f6d7baed9e761b69fb41442761ac6 = I29b4fdd4c13c96461c76660df767ea73(Ie791b43e8d5c9d1669743ea4d6e3139c[10]);
            Id5b4ee69444e5b499476c05a7f1d6e60 = I29b4fdd4c13c96461c76660df767ea73(Ie791b43e8d5c9d1669743ea4d6e3139c[11]);
            Id6105518ade80c89d4f20222a2382efb = I29b4fdd4c13c96461c76660df767ea73(Ie791b43e8d5c9d1669743ea4d6e3139c[12]);
            I26cf25e680483bf4e556d74efec35ee7 = I29b4fdd4c13c96461c76660df767ea73(Ie791b43e8d5c9d1669743ea4d6e3139c[13]);
            I8636f5c91b567780d3324e4b8a320fc2 = I29b4fdd4c13c96461c76660df767ea73(Ie791b43e8d5c9d1669743ea4d6e3139c[14]);
            I914bef0326cf82d350344317eb1359be = I29b4fdd4c13c96461c76660df767ea73(Ie791b43e8d5c9d1669743ea4d6e3139c[15]);
            I7de222bc26e38b8b6543819701740302 = I29b4fdd4c13c96461c76660df767ea73(Ie791b43e8d5c9d1669743ea4d6e3139c[16]);
            Ie3361a270ebc41698ef4651bb3548a49 = I29b4fdd4c13c96461c76660df767ea73(Ie791b43e8d5c9d1669743ea4d6e3139c[17]);
            I1240c9410b897a4d0504affca5ba139e = I29b4fdd4c13c96461c76660df767ea73(Ie791b43e8d5c9d1669743ea4d6e3139c[18]);
            If17b4f86674bc5fb212a1f7751fb043a = I29b4fdd4c13c96461c76660df767ea73(Ie791b43e8d5c9d1669743ea4d6e3139c[19]);
            I275f6334127640b2de3f0f87f54fd74c = I29b4fdd4c13c96461c76660df767ea73(Ie791b43e8d5c9d1669743ea4d6e3139c[20]);
            Iec844d10736440b96f9d6c651e604efd = I29b4fdd4c13c96461c76660df767ea73(Ie791b43e8d5c9d1669743ea4d6e3139c[21]);
            Ie04ce30f26a4ef1ee5b34474368dbac7 = I29b4fdd4c13c96461c76660df767ea73(I5b892f00b2642ca102f7755ab512d067[0]);
            Ibfee0b4ad5cdf16e88fcf469c5e031e9 = I29b4fdd4c13c96461c76660df767ea73(I5b892f00b2642ca102f7755ab512d067[1]);
            I3a4a965f22487553dec2a3e8e7836264 = I29b4fdd4c13c96461c76660df767ea73(I5b892f00b2642ca102f7755ab512d067[2]);
            I2a2d014f94d7a3b9fb3024a3e9107a73 = I29b4fdd4c13c96461c76660df767ea73(I5b892f00b2642ca102f7755ab512d067[3]);
            I5bab5ae46114c487f67b8e779d7461df = I29b4fdd4c13c96461c76660df767ea73(I5b892f00b2642ca102f7755ab512d067[4]);
            I45373bff54eccf8137da2931d841934e = I29b4fdd4c13c96461c76660df767ea73(I5b892f00b2642ca102f7755ab512d067[5]);
            Ib9322ec1d3866ba3cb42e96b5ff5cfb2 = I29b4fdd4c13c96461c76660df767ea73(I5b892f00b2642ca102f7755ab512d067[6]);
            I0a9cb91319cc0d0c1c4d0020cce321d7 = I29b4fdd4c13c96461c76660df767ea73(I5b892f00b2642ca102f7755ab512d067[7]);
            I299b37fd45c6ee2031fb2c74caac73be = I29b4fdd4c13c96461c76660df767ea73(I5b892f00b2642ca102f7755ab512d067[8]);
            Ic2f450f7ab60ba57dfc1406c92c0f077 = I29b4fdd4c13c96461c76660df767ea73(I5b892f00b2642ca102f7755ab512d067[9]);
            Ieca5b21b91e150c9d509964bdcea500d = I29b4fdd4c13c96461c76660df767ea73(I5b892f00b2642ca102f7755ab512d067[10]);
            I48b39ee498563e23c3a4be079b6100d8 = I29b4fdd4c13c96461c76660df767ea73(I5b892f00b2642ca102f7755ab512d067[11]);
            Iac8cb32c2d86b975f51a2ed605002e51 = I29b4fdd4c13c96461c76660df767ea73(I5b892f00b2642ca102f7755ab512d067[12]);
            Ic989dc794ce4356856b3916ab1889589 = I29b4fdd4c13c96461c76660df767ea73(I5b892f00b2642ca102f7755ab512d067[13]);
            Ie380b37a78242e6d45b659d568887457 = I29b4fdd4c13c96461c76660df767ea73(I5b892f00b2642ca102f7755ab512d067[14]);
            Ie43a7f8082f91c2955076a6373028b55 = I29b4fdd4c13c96461c76660df767ea73(I5b892f00b2642ca102f7755ab512d067[15]);
            Iea765ae5e9c65b3186445b15c56f69e5 = I29b4fdd4c13c96461c76660df767ea73(I5b892f00b2642ca102f7755ab512d067[16]);
            I74b55d2f94073ba8f948e4b02386867c = I29b4fdd4c13c96461c76660df767ea73(I5b892f00b2642ca102f7755ab512d067[17]);
            I015630502f5cb4eb27b2a673e810f1dc = I29b4fdd4c13c96461c76660df767ea73(I5b892f00b2642ca102f7755ab512d067[18]);
            I5085f161323433d8d38be2e4511b0c46 = I29b4fdd4c13c96461c76660df767ea73(I5b892f00b2642ca102f7755ab512d067[19]);
            Ie9fd8f7dc0c3849c0437a2a3d8607b4c = I29b4fdd4c13c96461c76660df767ea73(I5b892f00b2642ca102f7755ab512d067[20]);
            I9306d9ef7934ffe5902306b9783c351e = I29b4fdd4c13c96461c76660df767ea73(I5b892f00b2642ca102f7755ab512d067[21]);
            I70e68beb262fbdeba621b3794adf9f84 = I29b4fdd4c13c96461c76660df767ea73(I8f906015dba99b4a73dcf767cbd948ee[0]);
            Ie7bf11bab3d601fd0a6e3eb415e263c8 = I29b4fdd4c13c96461c76660df767ea73(I8f906015dba99b4a73dcf767cbd948ee[1]);
            Ica3d4ebff001fb6ee69a66eb898eb5bd = I29b4fdd4c13c96461c76660df767ea73(I8f906015dba99b4a73dcf767cbd948ee[2]);
            I27951ef3d612004abdc639662807426b = I29b4fdd4c13c96461c76660df767ea73(I8f906015dba99b4a73dcf767cbd948ee[3]);
            Ice4f4ba8bb3381c8846941d5d5fe4534 = I29b4fdd4c13c96461c76660df767ea73(I8f906015dba99b4a73dcf767cbd948ee[4]);
            I223151b6414d9979d71023053dd3f5e2 = I29b4fdd4c13c96461c76660df767ea73(I8f906015dba99b4a73dcf767cbd948ee[5]);
            I73d2731c1b1ae5ef73ce0eb9c8995912 = I29b4fdd4c13c96461c76660df767ea73(I8f906015dba99b4a73dcf767cbd948ee[6]);
            I5ca15c7da1f49580ddedd9ff8ba822c0 = I29b4fdd4c13c96461c76660df767ea73(I8f906015dba99b4a73dcf767cbd948ee[7]);
            I8289bfc08a5d8979ec26825bcb6e3d18 = I29b4fdd4c13c96461c76660df767ea73(I8f906015dba99b4a73dcf767cbd948ee[8]);
            Ie3c88bc240576aa220f0f110b13bfdd3 = I29b4fdd4c13c96461c76660df767ea73(I8f906015dba99b4a73dcf767cbd948ee[9]);
            I583c6d23506c7d7b84403bfe977ec1ec = I29b4fdd4c13c96461c76660df767ea73(I8f906015dba99b4a73dcf767cbd948ee[10]);
            I768afe193d9d79b136736abc6846d945 = I29b4fdd4c13c96461c76660df767ea73(I8f906015dba99b4a73dcf767cbd948ee[11]);
            I277d7065150714e33d8ba64875d18190 = I29b4fdd4c13c96461c76660df767ea73(I8f906015dba99b4a73dcf767cbd948ee[12]);
            Ia5c77c9be26d62b026f24ee5a5e25fb8 = I29b4fdd4c13c96461c76660df767ea73(I8f906015dba99b4a73dcf767cbd948ee[13]);
            I88a325547ccfe4eabf90792abd60e356 = I29b4fdd4c13c96461c76660df767ea73(I8f906015dba99b4a73dcf767cbd948ee[14]);
            I21842d06e25948ef461d1fd03485f86c = I29b4fdd4c13c96461c76660df767ea73(I8f906015dba99b4a73dcf767cbd948ee[15]);
            Id65f22fa8fc9c47bfd00c796b63c9fa4 = I29b4fdd4c13c96461c76660df767ea73(I8f906015dba99b4a73dcf767cbd948ee[16]);
            I288ff69a7395e74f7de8da5a6a7f9062 = I29b4fdd4c13c96461c76660df767ea73(I8f906015dba99b4a73dcf767cbd948ee[17]);
            I2ba94ef71f97b9ba731b306d4a5fd02c = I29b4fdd4c13c96461c76660df767ea73(I8f906015dba99b4a73dcf767cbd948ee[18]);
            I26ae9e570a101c6f8237d7941285b924 = I29b4fdd4c13c96461c76660df767ea73(I8f906015dba99b4a73dcf767cbd948ee[19]);
            Icb92c7c10f0bfc5d287228f98d8a235c = I29b4fdd4c13c96461c76660df767ea73(I8f906015dba99b4a73dcf767cbd948ee[20]);
            Iba4972a3b71a3101ab23190ed905dc17 = I29b4fdd4c13c96461c76660df767ea73(I8f906015dba99b4a73dcf767cbd948ee[21]);
            I33703f538ec70268e6c00ad6eef6c4e0 = I29b4fdd4c13c96461c76660df767ea73(I8f906015dba99b4a73dcf767cbd948ee[22]);
            I71b93abe4b20e6a17ff17e0f33ac2ca5 = I29b4fdd4c13c96461c76660df767ea73(I9ab4bbe4191d0f284defcdce6b885054[0]);
            I91c2f3cdd7cc98a60090ec6e46d52ae7 = I29b4fdd4c13c96461c76660df767ea73(I9ab4bbe4191d0f284defcdce6b885054[1]);
            I4254f2987cd014ed703ae18e9963e585 = I29b4fdd4c13c96461c76660df767ea73(I9ab4bbe4191d0f284defcdce6b885054[2]);
            I9068cca0de6ecff56ca542d0998fcab2 = I29b4fdd4c13c96461c76660df767ea73(I9ab4bbe4191d0f284defcdce6b885054[3]);
            Ib3ec015a3d43d46e0b7142b21a81cfee = I29b4fdd4c13c96461c76660df767ea73(I9ab4bbe4191d0f284defcdce6b885054[4]);
            I8cb171677016e4309034dc5d83981a48 = I29b4fdd4c13c96461c76660df767ea73(I9ab4bbe4191d0f284defcdce6b885054[5]);
            I2a4b3573ae7c3b38ec34591f20c1d076 = I29b4fdd4c13c96461c76660df767ea73(I9ab4bbe4191d0f284defcdce6b885054[6]);
            I276c2ce5d3a1b7551c2790971071b094 = I29b4fdd4c13c96461c76660df767ea73(I9ab4bbe4191d0f284defcdce6b885054[7]);
            I9dff504e40aaddefedbb7b0f822c844a = I29b4fdd4c13c96461c76660df767ea73(I9ab4bbe4191d0f284defcdce6b885054[8]);
            I4ed5da534afbfe9ecbc10ef4cc649a55 = I29b4fdd4c13c96461c76660df767ea73(I9ab4bbe4191d0f284defcdce6b885054[9]);
            I618363a8ac413dd0ee52eb658940eaed = I29b4fdd4c13c96461c76660df767ea73(I9ab4bbe4191d0f284defcdce6b885054[10]);
            I54166b387c02e12374d6febc425bfb7a = I29b4fdd4c13c96461c76660df767ea73(I9ab4bbe4191d0f284defcdce6b885054[11]);
            I0b6cdfa1dbfa774fc9a12d856e61cddb = I29b4fdd4c13c96461c76660df767ea73(I9ab4bbe4191d0f284defcdce6b885054[12]);
            Ic4af6c9097257c9b22a57ce4b79b40fe = I29b4fdd4c13c96461c76660df767ea73(I9ab4bbe4191d0f284defcdce6b885054[13]);
            Iae21bdea20a6266d3f69aa680b6b2817 = I29b4fdd4c13c96461c76660df767ea73(I9ab4bbe4191d0f284defcdce6b885054[14]);
            I37e360420c7dd061de93a6647513676d = I29b4fdd4c13c96461c76660df767ea73(I9ab4bbe4191d0f284defcdce6b885054[15]);
            Ia81c31ea4f4786136b539c9766987596 = I29b4fdd4c13c96461c76660df767ea73(I9ab4bbe4191d0f284defcdce6b885054[16]);
            I5a4f0749acdc34fd0786e4b3d062f88b = I29b4fdd4c13c96461c76660df767ea73(I9ab4bbe4191d0f284defcdce6b885054[17]);
            I5529d6db17b6184c45cc4487e5a2c24a = I29b4fdd4c13c96461c76660df767ea73(I9ab4bbe4191d0f284defcdce6b885054[18]);
            Iabe5aea929c668c9b9728d073ffb00c8 = I29b4fdd4c13c96461c76660df767ea73(I9ab4bbe4191d0f284defcdce6b885054[19]);
            I4fb3fe065daa2708e55c812e57c19fb6 = I29b4fdd4c13c96461c76660df767ea73(I9ab4bbe4191d0f284defcdce6b885054[20]);
            I4bd98e902e805426fdd4606fcb5a5214 = I29b4fdd4c13c96461c76660df767ea73(I9ab4bbe4191d0f284defcdce6b885054[21]);
            Ia5e26c2417aba1005971749f4ab2f367 = I29b4fdd4c13c96461c76660df767ea73(I9ab4bbe4191d0f284defcdce6b885054[22]);
            I0e112f1d4e9c934a118f79f3856744a9 = I29b4fdd4c13c96461c76660df767ea73(Ic8a3b3e2aacd0eb24cbc429e9bb734ee[0]);
            I005e8b590924f9486cb23191d35c9797 = I29b4fdd4c13c96461c76660df767ea73(Ic8a3b3e2aacd0eb24cbc429e9bb734ee[1]);
            I8c5f98353b5b082dc3cf056469945a08 = I29b4fdd4c13c96461c76660df767ea73(Ic8a3b3e2aacd0eb24cbc429e9bb734ee[2]);
            I9aa11f30712f1779339b985212a7979c = I29b4fdd4c13c96461c76660df767ea73(Ic8a3b3e2aacd0eb24cbc429e9bb734ee[3]);
            I65928407b1d5447dbc815cd2d2e7b37d = I29b4fdd4c13c96461c76660df767ea73(Ic8a3b3e2aacd0eb24cbc429e9bb734ee[4]);
            If5b3850da967f6f3d7a71d680341ad1c = I29b4fdd4c13c96461c76660df767ea73(Ic8a3b3e2aacd0eb24cbc429e9bb734ee[5]);
            I0aa5522190c741b7df4c4d7d34e46987 = I29b4fdd4c13c96461c76660df767ea73(Ic8a3b3e2aacd0eb24cbc429e9bb734ee[6]);
            Iff777b2c4a3939e330c4cbb36cbe1ac5 = I29b4fdd4c13c96461c76660df767ea73(Ic8a3b3e2aacd0eb24cbc429e9bb734ee[7]);
            I2d839c10960739097d449efab58b9fd4 = I29b4fdd4c13c96461c76660df767ea73(Ic8a3b3e2aacd0eb24cbc429e9bb734ee[8]);
            Ice8765807beffd3acf59fa137ee0baac = I29b4fdd4c13c96461c76660df767ea73(Ic8a3b3e2aacd0eb24cbc429e9bb734ee[9]);
            I529eaa7e5eeb6d0a1aba78df5d5a2fa0 = I29b4fdd4c13c96461c76660df767ea73(Ic8a3b3e2aacd0eb24cbc429e9bb734ee[10]);
            Icb2805685607d5fedd0300c9d800f863 = I29b4fdd4c13c96461c76660df767ea73(Ic8a3b3e2aacd0eb24cbc429e9bb734ee[11]);
            Idadf072247b351cf51d718f797c3b375 = I29b4fdd4c13c96461c76660df767ea73(Ic8a3b3e2aacd0eb24cbc429e9bb734ee[12]);
            I6fcb3b133a6a654b69f41468a713d922 = I29b4fdd4c13c96461c76660df767ea73(Ic8a3b3e2aacd0eb24cbc429e9bb734ee[13]);
            I77e1f5f504a794edbb89c66cf1ffcf66 = I29b4fdd4c13c96461c76660df767ea73(Ic8a3b3e2aacd0eb24cbc429e9bb734ee[14]);
            I185085cbf8da6df921ba32442b28bcca = I29b4fdd4c13c96461c76660df767ea73(Ic8a3b3e2aacd0eb24cbc429e9bb734ee[15]);
            Ibcb80df5bed66f8498561e3f3ffa4ec4 = I29b4fdd4c13c96461c76660df767ea73(Ic8a3b3e2aacd0eb24cbc429e9bb734ee[16]);
            I2cf5304a672431888916e08b3c15f0c7 = I29b4fdd4c13c96461c76660df767ea73(Ic8a3b3e2aacd0eb24cbc429e9bb734ee[17]);
            Icf266f710358631b7119ef526acb301c = I29b4fdd4c13c96461c76660df767ea73(Ic8a3b3e2aacd0eb24cbc429e9bb734ee[18]);
            Ia209e5b03deaf4fcb8ae12b731a49e0a = I29b4fdd4c13c96461c76660df767ea73(Ic8a3b3e2aacd0eb24cbc429e9bb734ee[19]);
            Iffb7fe9c74dfc01a43e99a099c4e7e04 = I29b4fdd4c13c96461c76660df767ea73(Ic8a3b3e2aacd0eb24cbc429e9bb734ee[20]);
            I43f52bcba1bd2e8ee5fac03320e4f19f = I29b4fdd4c13c96461c76660df767ea73(Ic8a3b3e2aacd0eb24cbc429e9bb734ee[21]);
            I9fdfe73e77c384d33196c0f2d2a2fde2 = I29b4fdd4c13c96461c76660df767ea73(Ic8a3b3e2aacd0eb24cbc429e9bb734ee[22]);
            I546657528d591e8bb44c32fed7707af5 = I29b4fdd4c13c96461c76660df767ea73(I6ff6fafd1a3364131b269724ad273ba5[0]);
            I6e4ae763dc4e8aa8afc4599de96c75d3 = I29b4fdd4c13c96461c76660df767ea73(I6ff6fafd1a3364131b269724ad273ba5[1]);
            Id8c36004ae8e550569a491f6b514945a = I29b4fdd4c13c96461c76660df767ea73(I6ff6fafd1a3364131b269724ad273ba5[2]);
            I111ac0aadbdd3e4479ca0786491a7b08 = I29b4fdd4c13c96461c76660df767ea73(I6ff6fafd1a3364131b269724ad273ba5[3]);
            Ib83242b57ab050b0e5f9bdf91fa118fb = I29b4fdd4c13c96461c76660df767ea73(I6ff6fafd1a3364131b269724ad273ba5[4]);
            I7be8b2f8a9fe8e13001c2a1fce4a8a3f = I29b4fdd4c13c96461c76660df767ea73(I6ff6fafd1a3364131b269724ad273ba5[5]);
            If4d030e5858f325debc6f37abf4a7d6c = I29b4fdd4c13c96461c76660df767ea73(I6ff6fafd1a3364131b269724ad273ba5[6]);
            I627e4bdc8061c69e3fcac17535b9f1e0 = I29b4fdd4c13c96461c76660df767ea73(I6ff6fafd1a3364131b269724ad273ba5[7]);
            Ia443284a35e0873de59b3ae55b7f809d = I29b4fdd4c13c96461c76660df767ea73(I6ff6fafd1a3364131b269724ad273ba5[8]);
            Ibafedcf9f2990ed9c1efa973a0b1d81d = I29b4fdd4c13c96461c76660df767ea73(I6ff6fafd1a3364131b269724ad273ba5[9]);
            I439c7c302b535bfd7db655c3c607d71f = I29b4fdd4c13c96461c76660df767ea73(I6ff6fafd1a3364131b269724ad273ba5[10]);
            I2133d362ba45ceb3dceaa84e95ace1e6 = I29b4fdd4c13c96461c76660df767ea73(I6ff6fafd1a3364131b269724ad273ba5[11]);
            I67534b68fee8f76ac0c5e64cd02aba42 = I29b4fdd4c13c96461c76660df767ea73(I6ff6fafd1a3364131b269724ad273ba5[12]);
            I8613cac4ccd4f956e8a0ae7b627f5be2 = I29b4fdd4c13c96461c76660df767ea73(I6ff6fafd1a3364131b269724ad273ba5[13]);
            I8493e2dac01f009db1d2d5504b49d135 = I29b4fdd4c13c96461c76660df767ea73(I6ff6fafd1a3364131b269724ad273ba5[14]);
            I5c278aad08b7c4b0237d68f88fcb3f3a = I29b4fdd4c13c96461c76660df767ea73(I6ff6fafd1a3364131b269724ad273ba5[15]);
            Iba75ff0f3b67c7e28cf627706733d528 = I29b4fdd4c13c96461c76660df767ea73(I6ff6fafd1a3364131b269724ad273ba5[16]);
            I9164fa2a9a33da6612ea692cf3fa7d2f = I29b4fdd4c13c96461c76660df767ea73(I6ff6fafd1a3364131b269724ad273ba5[17]);
            I0f3c4fb63ef1e88168b4d28175a0b68c = I29b4fdd4c13c96461c76660df767ea73(I6ff6fafd1a3364131b269724ad273ba5[18]);
            I99d236d41be79090ca7ba1fb6faaec4c = I29b4fdd4c13c96461c76660df767ea73(I6ff6fafd1a3364131b269724ad273ba5[19]);
            I487b9b236d118786e475ccc5e4e56a6d = I29b4fdd4c13c96461c76660df767ea73(I6ff6fafd1a3364131b269724ad273ba5[20]);
            I6cb09ac924c3b3b44443263e08c3315c = I29b4fdd4c13c96461c76660df767ea73(I6ff6fafd1a3364131b269724ad273ba5[21]);
            Id924dafd31fd0af0b28c7e6b7e95ec37 = I29b4fdd4c13c96461c76660df767ea73(I6ff6fafd1a3364131b269724ad273ba5[22]);
            I9184110e3e9b8614460fc0abe5fff2d9 = I29b4fdd4c13c96461c76660df767ea73(I154fcd3171f1231e825ee603d53ecfe8[0]);
            If8865fee7dbf593b34ea54692d947f10 = I29b4fdd4c13c96461c76660df767ea73(I154fcd3171f1231e825ee603d53ecfe8[1]);
            I4854ff71aa885da3d07acaaa24740d7c = I29b4fdd4c13c96461c76660df767ea73(I154fcd3171f1231e825ee603d53ecfe8[2]);
            Ie8befb003fe83e774e8d1d01d4e2f4ad = I29b4fdd4c13c96461c76660df767ea73(I154fcd3171f1231e825ee603d53ecfe8[3]);
            Ie7e196fbb66ba6bee51ef0064ca519c2 = I29b4fdd4c13c96461c76660df767ea73(I154fcd3171f1231e825ee603d53ecfe8[4]);
            I685699f60c76b00df87c9c53e9a8e448 = I29b4fdd4c13c96461c76660df767ea73(I154fcd3171f1231e825ee603d53ecfe8[5]);
            Ib6c0e635e659f54724737f0cffd1b0fc = I29b4fdd4c13c96461c76660df767ea73(I154fcd3171f1231e825ee603d53ecfe8[6]);
            I3a8bcfdab631a268d21c87b98e9d1c49 = I29b4fdd4c13c96461c76660df767ea73(I154fcd3171f1231e825ee603d53ecfe8[7]);
            I3faeba79f7af7a006ab5cd256352e2db = I29b4fdd4c13c96461c76660df767ea73(I154fcd3171f1231e825ee603d53ecfe8[8]);
            I02e672436ade3ee620c72c0d9ceee664 = I29b4fdd4c13c96461c76660df767ea73(I154fcd3171f1231e825ee603d53ecfe8[9]);
            I65708fb59e90bb79b8107da619fe63eb = I29b4fdd4c13c96461c76660df767ea73(I489e70342dbba4a551097e3064dc9835[0]);
            I840a1a7c0bf49f4f42499b33f32fa02d = I29b4fdd4c13c96461c76660df767ea73(I489e70342dbba4a551097e3064dc9835[1]);
            If7543e2f5a158b1f3f3a4078ec54cab5 = I29b4fdd4c13c96461c76660df767ea73(I489e70342dbba4a551097e3064dc9835[2]);
            I98a2aa729628adde0b6047869bd12743 = I29b4fdd4c13c96461c76660df767ea73(I489e70342dbba4a551097e3064dc9835[3]);
            Ibfb57f2b507c27759a3556759f23977b = I29b4fdd4c13c96461c76660df767ea73(I489e70342dbba4a551097e3064dc9835[4]);
            Ib20dec1346f227042c749ec1abfa4d39 = I29b4fdd4c13c96461c76660df767ea73(I489e70342dbba4a551097e3064dc9835[5]);
            Ifba318d4faf308168c5eac8fe92395b4 = I29b4fdd4c13c96461c76660df767ea73(I489e70342dbba4a551097e3064dc9835[6]);
            I95b923444062b4a98918c685c65996d0 = I29b4fdd4c13c96461c76660df767ea73(I489e70342dbba4a551097e3064dc9835[7]);
            I45a6ef43e6e42594444adcbda26700ab = I29b4fdd4c13c96461c76660df767ea73(I489e70342dbba4a551097e3064dc9835[8]);
            I508cea40d87bec2672f980d145c89b55 = I29b4fdd4c13c96461c76660df767ea73(I489e70342dbba4a551097e3064dc9835[9]);
            I0ace1d51fdee91f8f3826a945c4e66a4 = I29b4fdd4c13c96461c76660df767ea73(I0b0a1f577a212bd9024c8b9a44c92e00[0]);
            I99ff3922e018c409dc8ce5f3503e3c56 = I29b4fdd4c13c96461c76660df767ea73(I0b0a1f577a212bd9024c8b9a44c92e00[1]);
            I6a3824a6598bbaa138e1e763ad85f5f7 = I29b4fdd4c13c96461c76660df767ea73(I0b0a1f577a212bd9024c8b9a44c92e00[2]);
            I283107989a436e2c720123b8d9e335c2 = I29b4fdd4c13c96461c76660df767ea73(I0b0a1f577a212bd9024c8b9a44c92e00[3]);
            I7b12345fe53174cadef6811fb8869b42 = I29b4fdd4c13c96461c76660df767ea73(I0b0a1f577a212bd9024c8b9a44c92e00[4]);
            Iac6fcccf3a0cfe04edc0d998b60c2681 = I29b4fdd4c13c96461c76660df767ea73(I0b0a1f577a212bd9024c8b9a44c92e00[5]);
            Ic9678deca4bf44a7b99f853334f6a05c = I29b4fdd4c13c96461c76660df767ea73(I0b0a1f577a212bd9024c8b9a44c92e00[6]);
            Ie40c90fdb38b3e4046ba89295ed77d7c = I29b4fdd4c13c96461c76660df767ea73(I0b0a1f577a212bd9024c8b9a44c92e00[7]);
            Iea4a7766d3b9d5d030ade1739859ef0d = I29b4fdd4c13c96461c76660df767ea73(I0b0a1f577a212bd9024c8b9a44c92e00[8]);
            I844b9a89ffb7a5e48979fdea546e244a = I29b4fdd4c13c96461c76660df767ea73(I0b0a1f577a212bd9024c8b9a44c92e00[9]);
            I656852be6f5b3542862e0f68d48be518 = I29b4fdd4c13c96461c76660df767ea73(I40d311bab75b73e3788c50115a205270[0]);
            Id6551b6b053952162b90792ab73a1a49 = I29b4fdd4c13c96461c76660df767ea73(I40d311bab75b73e3788c50115a205270[1]);
            Ib7fde6a2ec1ff0a3af10bccf3012e63f = I29b4fdd4c13c96461c76660df767ea73(I40d311bab75b73e3788c50115a205270[2]);
            I989091b3586964ab598f166a89279d16 = I29b4fdd4c13c96461c76660df767ea73(I40d311bab75b73e3788c50115a205270[3]);
            I9785922874bba479ce4a9bf1759e2933 = I29b4fdd4c13c96461c76660df767ea73(I40d311bab75b73e3788c50115a205270[4]);
            Ifbaae8b3da03911a4c96d4efdb9283c5 = I29b4fdd4c13c96461c76660df767ea73(I40d311bab75b73e3788c50115a205270[5]);
            I77a54091bc2c3d9006ecb3471b94d8c8 = I29b4fdd4c13c96461c76660df767ea73(I40d311bab75b73e3788c50115a205270[6]);
            I9859b94cda465ceaaa5674eb19e94824 = I29b4fdd4c13c96461c76660df767ea73(I40d311bab75b73e3788c50115a205270[7]);
            I5a7746e9fbb8c009f83ae57423296cdf = I29b4fdd4c13c96461c76660df767ea73(I40d311bab75b73e3788c50115a205270[8]);
            Ibddcc2e26fba20dfe2a2d399be2bc45b = I29b4fdd4c13c96461c76660df767ea73(I40d311bab75b73e3788c50115a205270[9]);
            I8dbe6497a8deabcc60783bfe7548d0fb = I29b4fdd4c13c96461c76660df767ea73(I5fa015a360308bffc46921d119b60c1b[0]);
            Ifef870b405335975988b58b2273d4e1a = I29b4fdd4c13c96461c76660df767ea73(I5fa015a360308bffc46921d119b60c1b[1]);
            Ic1f6842b4f246d624d91daa6ada10ca9 = I29b4fdd4c13c96461c76660df767ea73(I5fa015a360308bffc46921d119b60c1b[2]);
            Ibc8679379ddc43ee4bc508a1f577eb2c = I29b4fdd4c13c96461c76660df767ea73(I5fa015a360308bffc46921d119b60c1b[3]);
            Ibdd9957b7f1a319b797c021933ff75d7 = I29b4fdd4c13c96461c76660df767ea73(I5fa015a360308bffc46921d119b60c1b[4]);
            I041f9455435bfa375395eb330a34993d = I29b4fdd4c13c96461c76660df767ea73(I9e42bc767599ce3cc4e2d886e5ef2e62[0]);
            Ifbe29365e7035c78af9f42902b0d303e = I29b4fdd4c13c96461c76660df767ea73(I9e42bc767599ce3cc4e2d886e5ef2e62[1]);
            Ic8759e2f58848b33082bd1b02acc9c0b = I29b4fdd4c13c96461c76660df767ea73(I9e42bc767599ce3cc4e2d886e5ef2e62[2]);
            Ie2e3d64640c339dc51512979dbd6a173 = I29b4fdd4c13c96461c76660df767ea73(I9e42bc767599ce3cc4e2d886e5ef2e62[3]);
            Ib2c327648cce481482eaf0467e9227d4 = I29b4fdd4c13c96461c76660df767ea73(I9e42bc767599ce3cc4e2d886e5ef2e62[4]);
            I535cad8c919a4330257eb5b4bed61b3a = I29b4fdd4c13c96461c76660df767ea73(Iea43b150eabf3c7781275821eee3e0c1[0]);
            Ib2afdf9534deaae465d99b7e377788bb = I29b4fdd4c13c96461c76660df767ea73(Iea43b150eabf3c7781275821eee3e0c1[1]);
            I6eaffd980e4d77fdbda5e63bad9489d7 = I29b4fdd4c13c96461c76660df767ea73(Iea43b150eabf3c7781275821eee3e0c1[2]);
            I6e4786234b286b12c83e06e93c628534 = I29b4fdd4c13c96461c76660df767ea73(Iea43b150eabf3c7781275821eee3e0c1[3]);
            Idcc745602c4b7b34df9c3d68f9a9d76d = I29b4fdd4c13c96461c76660df767ea73(Iea43b150eabf3c7781275821eee3e0c1[4]);
            I0fc42ce9cc31d781ea3013318c25a571 = I29b4fdd4c13c96461c76660df767ea73(I8012eea3d53fa4e000eb28b121e02ada[0]);
            I4363ca6b3d9ca9863f70958aa7c23777 = I29b4fdd4c13c96461c76660df767ea73(I8012eea3d53fa4e000eb28b121e02ada[1]);
            Ic902e09b33db1b919c102f7971cdef7b = I29b4fdd4c13c96461c76660df767ea73(I8012eea3d53fa4e000eb28b121e02ada[2]);
            Icf4405d4a4063448a2be8ad0354ab1a8 = I29b4fdd4c13c96461c76660df767ea73(I8012eea3d53fa4e000eb28b121e02ada[3]);
            I72108531a608f6d5e51a481c68d7b271 = I29b4fdd4c13c96461c76660df767ea73(I8012eea3d53fa4e000eb28b121e02ada[4]);
            I6922b510e432e06d209095bcc6297e7e = I29b4fdd4c13c96461c76660df767ea73(I49804415d20c0c087f802b25dd609887[0]);
            Ief90f8a8efca2b06eff0d4cba1cbb342 = I29b4fdd4c13c96461c76660df767ea73(I49804415d20c0c087f802b25dd609887[1]);
            Ib5334df42ee8f1574e41cb30b903fae9 = I29b4fdd4c13c96461c76660df767ea73(I49804415d20c0c087f802b25dd609887[2]);
            I535b29f7177b4fc009ee998f1f4f7d7f = I29b4fdd4c13c96461c76660df767ea73(I49804415d20c0c087f802b25dd609887[3]);
            Id0842da8068ee88d99af7acea50e7b77 = I29b4fdd4c13c96461c76660df767ea73(I49804415d20c0c087f802b25dd609887[4]);
            Ib6cdbbb765694d822639b7c8fbfc50c4 = I29b4fdd4c13c96461c76660df767ea73(Id270f05bf5c3fc0bb211d1665d149044[0]);
            Ibdaa6d215d34aa0cc27d5234da6fd991 = I29b4fdd4c13c96461c76660df767ea73(Id270f05bf5c3fc0bb211d1665d149044[1]);
            Id769d4a92f5f6da262ce0521e5509368 = I29b4fdd4c13c96461c76660df767ea73(Id270f05bf5c3fc0bb211d1665d149044[2]);
            Iaf3a0b5ea5d9eda47fcced9260922bc6 = I29b4fdd4c13c96461c76660df767ea73(Id270f05bf5c3fc0bb211d1665d149044[3]);
            I03a8a458ee0942c35001cbfe8e589222 = I29b4fdd4c13c96461c76660df767ea73(Id270f05bf5c3fc0bb211d1665d149044[4]);
            I25eb943ea517a4827efb1e797bfdc4f5 = I29b4fdd4c13c96461c76660df767ea73(If091fe044c792be711325c103b84cf1d[0]);
            Iac4b8906947fc90bfe76cee2f1d4c4ab = I29b4fdd4c13c96461c76660df767ea73(If091fe044c792be711325c103b84cf1d[1]);
            I58a490344f87b4d5bb319e3e85ba9278 = I29b4fdd4c13c96461c76660df767ea73(If091fe044c792be711325c103b84cf1d[2]);
            I9222c4c0eb2b110fd80547d46ba17036 = I29b4fdd4c13c96461c76660df767ea73(If091fe044c792be711325c103b84cf1d[3]);
            Ic1af7410a9d11c5324f3ee5b2e0e9dac = I29b4fdd4c13c96461c76660df767ea73(If091fe044c792be711325c103b84cf1d[4]);
            I9e0a36d0be66b4c02b03e5b75b686226 = I29b4fdd4c13c96461c76660df767ea73(I1550db301291ab131a5536147fb938f6[0]);
            I1eef40a71c8d1e2da9802929a5347e90 = I29b4fdd4c13c96461c76660df767ea73(I1550db301291ab131a5536147fb938f6[1]);
            Ied41909cd443432dafadba42672151c1 = I29b4fdd4c13c96461c76660df767ea73(I1550db301291ab131a5536147fb938f6[2]);
            Ib2c1636a66f6479d6123a038cbc668d5 = I29b4fdd4c13c96461c76660df767ea73(I1550db301291ab131a5536147fb938f6[3]);
            Ica02d19b129c8b1d491ea4747a55113e = I29b4fdd4c13c96461c76660df767ea73(I1550db301291ab131a5536147fb938f6[4]);
            I31bf4597a3b776962f5c820378254065 = I29b4fdd4c13c96461c76660df767ea73(I74d1345ee56f5688f875823a5d7c1f4f[0]);
            I58361fb97f1b5aff0a2751d35c8da672 = I29b4fdd4c13c96461c76660df767ea73(I74d1345ee56f5688f875823a5d7c1f4f[1]);
            I8ab7efc436a0f2cc3efbc299a0ddf914 = I29b4fdd4c13c96461c76660df767ea73(I74d1345ee56f5688f875823a5d7c1f4f[2]);
            I3934ed7170967ff3852944cc39ba1de9 = I29b4fdd4c13c96461c76660df767ea73(I74d1345ee56f5688f875823a5d7c1f4f[3]);
            Ic690477b1672dea4905a5e1c92b47366 = I29b4fdd4c13c96461c76660df767ea73(I74d1345ee56f5688f875823a5d7c1f4f[4]);
            I5eaa11e26f19b94dcb7eaee7f09d24b4 = I29b4fdd4c13c96461c76660df767ea73(I74d1345ee56f5688f875823a5d7c1f4f[5]);
            Iaf1d3be13e6441a7a9ab3f286a7dc21b = I29b4fdd4c13c96461c76660df767ea73(I74d1345ee56f5688f875823a5d7c1f4f[6]);
            I61f5ebea2bbe443b644c95ee559c2234 = I29b4fdd4c13c96461c76660df767ea73(I74d1345ee56f5688f875823a5d7c1f4f[7]);
            I1fbcaf2f6be01b129ebc24dee8a65396 = I29b4fdd4c13c96461c76660df767ea73(I74d1345ee56f5688f875823a5d7c1f4f[8]);
            I1c0df8c2c64b688ae417a238263f33db = I29b4fdd4c13c96461c76660df767ea73(I74d1345ee56f5688f875823a5d7c1f4f[9]);
            I4f169c2c8c0768f2725ed655a03acfc2 = I29b4fdd4c13c96461c76660df767ea73(I74d1345ee56f5688f875823a5d7c1f4f[10]);
            I96f65790e2cacf7b529ce5b88598da00 = I29b4fdd4c13c96461c76660df767ea73(I74d1345ee56f5688f875823a5d7c1f4f[11]);
            I6b5720d71a0b4cd10ea34affa6631a25 = I29b4fdd4c13c96461c76660df767ea73(I74d1345ee56f5688f875823a5d7c1f4f[12]);
            Ifc7eec6765af08463751db128f8818b3 = I29b4fdd4c13c96461c76660df767ea73(I74d1345ee56f5688f875823a5d7c1f4f[13]);
            I8dddcade21ad3bb330c1c25970c32b73 = I29b4fdd4c13c96461c76660df767ea73(I187371a49a27a988920854b2bb61bea5[0]);
            I74a7b85ddacad06ab1c6b0db9b084bd3 = I29b4fdd4c13c96461c76660df767ea73(I187371a49a27a988920854b2bb61bea5[1]);
            I2b0b168ce4fe8aa4a2e7cb69fe532aa3 = I29b4fdd4c13c96461c76660df767ea73(I187371a49a27a988920854b2bb61bea5[2]);
            I3e8d26ea83937cae01aadf1092c59bdf = I29b4fdd4c13c96461c76660df767ea73(I187371a49a27a988920854b2bb61bea5[3]);
            I90a4190941651d885d04deb86a163365 = I29b4fdd4c13c96461c76660df767ea73(I187371a49a27a988920854b2bb61bea5[4]);
            I7d85b73e85379bf3a480e954c05516f3 = I29b4fdd4c13c96461c76660df767ea73(I187371a49a27a988920854b2bb61bea5[5]);
            Id5c9a9b9c34c8f9d56df0aa8d780c9d3 = I29b4fdd4c13c96461c76660df767ea73(I187371a49a27a988920854b2bb61bea5[6]);
            I21255a0ad20a9668c958faf68d53b2bc = I29b4fdd4c13c96461c76660df767ea73(I187371a49a27a988920854b2bb61bea5[7]);
            Ifba1584d599da13b98a3b76b4db10974 = I29b4fdd4c13c96461c76660df767ea73(I187371a49a27a988920854b2bb61bea5[8]);
            Iad0f4602ec545dc6ef12aa34add00ed3 = I29b4fdd4c13c96461c76660df767ea73(I187371a49a27a988920854b2bb61bea5[9]);
            I8bb46c3eb9f54c5d1b28dc6aa0154358 = I29b4fdd4c13c96461c76660df767ea73(I187371a49a27a988920854b2bb61bea5[10]);
            Ic09b4671e867144fe9f54a09e74c5519 = I29b4fdd4c13c96461c76660df767ea73(I187371a49a27a988920854b2bb61bea5[11]);
            I391a2f354262558ff17d7d80b8c39e8c = I29b4fdd4c13c96461c76660df767ea73(I187371a49a27a988920854b2bb61bea5[12]);
            If6b40a030cb120fe017bf9d39e1a35d1 = I29b4fdd4c13c96461c76660df767ea73(I187371a49a27a988920854b2bb61bea5[13]);
            I490996026af34eba5bcd8d553af818eb = I29b4fdd4c13c96461c76660df767ea73(I48c4c6e7414394e3aeff9d17ec25d020[0]);
            Icbc12ab47f586b12402ae5d4361c967d = I29b4fdd4c13c96461c76660df767ea73(I48c4c6e7414394e3aeff9d17ec25d020[1]);
            Iee0e45914c52a357e1e32922299d6937 = I29b4fdd4c13c96461c76660df767ea73(I48c4c6e7414394e3aeff9d17ec25d020[2]);
            Iefe423653d454e21324a6857b52f98ac = I29b4fdd4c13c96461c76660df767ea73(I48c4c6e7414394e3aeff9d17ec25d020[3]);
            I6d6a242cdfadfc97fe656510bef73adc = I29b4fdd4c13c96461c76660df767ea73(I48c4c6e7414394e3aeff9d17ec25d020[4]);
            Ib5c8d91204a2d313c9c23110a53cd0cf = I29b4fdd4c13c96461c76660df767ea73(I48c4c6e7414394e3aeff9d17ec25d020[5]);
            Ic9740baafb1c92e3a25f0a1e7bc46486 = I29b4fdd4c13c96461c76660df767ea73(I48c4c6e7414394e3aeff9d17ec25d020[6]);
            I6f69796a6fe6da57066319ec8210c1a3 = I29b4fdd4c13c96461c76660df767ea73(I48c4c6e7414394e3aeff9d17ec25d020[7]);
            Idb862697f62a6c678072de760e176096 = I29b4fdd4c13c96461c76660df767ea73(I48c4c6e7414394e3aeff9d17ec25d020[8]);
            I06e05a1ed002175a75d02b8b76f52c50 = I29b4fdd4c13c96461c76660df767ea73(I48c4c6e7414394e3aeff9d17ec25d020[9]);
            I1e110e27162231650875dd1152d96e64 = I29b4fdd4c13c96461c76660df767ea73(I48c4c6e7414394e3aeff9d17ec25d020[10]);
            Ic46357bb77f6183329946f7e28294365 = I29b4fdd4c13c96461c76660df767ea73(I48c4c6e7414394e3aeff9d17ec25d020[11]);
            I8741c5cc763512d16cb1186fa3323f45 = I29b4fdd4c13c96461c76660df767ea73(I48c4c6e7414394e3aeff9d17ec25d020[12]);
            I30b5c7aadb5312ce96e833704bb3a320 = I29b4fdd4c13c96461c76660df767ea73(I48c4c6e7414394e3aeff9d17ec25d020[13]);
            If404a00ab81d6ebbc0dbdf4aecdce389 = I29b4fdd4c13c96461c76660df767ea73(I3cba0f4c2ca8c7c200df8e1071ab429d[0]);
            I19875f52f79482b477f1febaa7e97090 = I29b4fdd4c13c96461c76660df767ea73(I3cba0f4c2ca8c7c200df8e1071ab429d[1]);
            Ic7855ca956651bd368cbdde7ec93ba6d = I29b4fdd4c13c96461c76660df767ea73(I3cba0f4c2ca8c7c200df8e1071ab429d[2]);
            Ic57a2627a194099105a2908a41feddfb = I29b4fdd4c13c96461c76660df767ea73(I3cba0f4c2ca8c7c200df8e1071ab429d[3]);
            I4d1ba6ee8fb9505ba3b58b2b7553245b = I29b4fdd4c13c96461c76660df767ea73(I3cba0f4c2ca8c7c200df8e1071ab429d[4]);
            Ieb7b388ff89e352dd239e0ccbe7b9ecc = I29b4fdd4c13c96461c76660df767ea73(I3cba0f4c2ca8c7c200df8e1071ab429d[5]);
            Ib1461f456ebc14f449eee77e386a4c69 = I29b4fdd4c13c96461c76660df767ea73(I3cba0f4c2ca8c7c200df8e1071ab429d[6]);
            I8786eb767f02164cdc32f14f41b5d0e1 = I29b4fdd4c13c96461c76660df767ea73(I3cba0f4c2ca8c7c200df8e1071ab429d[7]);
            Id6fa8ec5d1062fc3e09bdac65ff79f45 = I29b4fdd4c13c96461c76660df767ea73(I3cba0f4c2ca8c7c200df8e1071ab429d[8]);
            I83b77ad1a40dc102f28153f692516eb4 = I29b4fdd4c13c96461c76660df767ea73(I3cba0f4c2ca8c7c200df8e1071ab429d[9]);
            I55e54359961ef6e5a63f1c2eb0ad4aa1 = I29b4fdd4c13c96461c76660df767ea73(I3cba0f4c2ca8c7c200df8e1071ab429d[10]);
            I90001da8c360ccff128f637cd672ad42 = I29b4fdd4c13c96461c76660df767ea73(I3cba0f4c2ca8c7c200df8e1071ab429d[11]);
            Ib38a46dc131d635b81fb7c196110fc4b = I29b4fdd4c13c96461c76660df767ea73(I3cba0f4c2ca8c7c200df8e1071ab429d[12]);
            I926c049036f53f0a0a6ad369de116c57 = I29b4fdd4c13c96461c76660df767ea73(I3cba0f4c2ca8c7c200df8e1071ab429d[13]);
            Iac48d2ccf6c6e0c555e874ae77123f2e = I29b4fdd4c13c96461c76660df767ea73(I35688678e1a83ec39d737d9cdfd44ba3[0]);
            Ic6f40833f5f6284c9015304fd3fc00f0 = I29b4fdd4c13c96461c76660df767ea73(I35688678e1a83ec39d737d9cdfd44ba3[1]);
            I3f2507530dd648814af0964f7da11d35 = I29b4fdd4c13c96461c76660df767ea73(I35688678e1a83ec39d737d9cdfd44ba3[2]);
            Id9edc6ac95a260bf5af3de25f00e9e9c = I29b4fdd4c13c96461c76660df767ea73(I35688678e1a83ec39d737d9cdfd44ba3[3]);
            I28fa295ebd90c2b7255d48ca9ffcfcf3 = I29b4fdd4c13c96461c76660df767ea73(I35688678e1a83ec39d737d9cdfd44ba3[4]);
            Ia308e09137af1cb50167562efb5da628 = I29b4fdd4c13c96461c76660df767ea73(I35688678e1a83ec39d737d9cdfd44ba3[5]);
            I5aa85d9503b0e4ff46bbd63e873053ca = I29b4fdd4c13c96461c76660df767ea73(I35688678e1a83ec39d737d9cdfd44ba3[6]);
            I7ea8fe50c45e213f3257060e2813240b = I29b4fdd4c13c96461c76660df767ea73(I94b86d31e8226723950096e91855b6d3[0]);
            Ic3e6e38a2986c7f14fd0db2246367a1c = I29b4fdd4c13c96461c76660df767ea73(I94b86d31e8226723950096e91855b6d3[1]);
            I581eb136fdd08302e02c1fafb5d5c90b = I29b4fdd4c13c96461c76660df767ea73(I94b86d31e8226723950096e91855b6d3[2]);
            I080832c25509f7003ed50d71210bc7f7 = I29b4fdd4c13c96461c76660df767ea73(I94b86d31e8226723950096e91855b6d3[3]);
            Ib43383830037df764b48c637a28ab6b5 = I29b4fdd4c13c96461c76660df767ea73(I94b86d31e8226723950096e91855b6d3[4]);
            Iddf65ccb4396288264a400ba37cbb655 = I29b4fdd4c13c96461c76660df767ea73(I94b86d31e8226723950096e91855b6d3[5]);
            Ia7673d73f0535906a99d6cb467892104 = I29b4fdd4c13c96461c76660df767ea73(I94b86d31e8226723950096e91855b6d3[6]);
            I8bc3210e86a523accdbeefe7e72ee4fc = I29b4fdd4c13c96461c76660df767ea73(I0ea7c4721ee0c13ad15a9b0fa7b15ad3[0]);
            Ib63574478126e6ee30a388d9648cb548 = I29b4fdd4c13c96461c76660df767ea73(I0ea7c4721ee0c13ad15a9b0fa7b15ad3[1]);
            Ic4501a8a1fb34c30a97e18a0ab189e3a = I29b4fdd4c13c96461c76660df767ea73(I0ea7c4721ee0c13ad15a9b0fa7b15ad3[2]);
            I2b807c16cfc6d65cb2a7f28ffa837974 = I29b4fdd4c13c96461c76660df767ea73(I0ea7c4721ee0c13ad15a9b0fa7b15ad3[3]);
            I0aa93075086164fdbab3814d60633141 = I29b4fdd4c13c96461c76660df767ea73(I0ea7c4721ee0c13ad15a9b0fa7b15ad3[4]);
            I886750aaf8d2040c3f12ff113294f658 = I29b4fdd4c13c96461c76660df767ea73(I0ea7c4721ee0c13ad15a9b0fa7b15ad3[5]);
            I103ec7cf279f527fc6e3648a19a12a8a = I29b4fdd4c13c96461c76660df767ea73(I0ea7c4721ee0c13ad15a9b0fa7b15ad3[6]);
            I9a57f2f03cf8a154c3a7d48ec089306d = I29b4fdd4c13c96461c76660df767ea73(I29dd5fb1c2673cd4daa9cafaf24d8e7c[0]);
            I9d8f8c1792427975a9e7024041f59be9 = I29b4fdd4c13c96461c76660df767ea73(I29dd5fb1c2673cd4daa9cafaf24d8e7c[1]);
            Ie8644d7edbadf19937c399cf275946e5 = I29b4fdd4c13c96461c76660df767ea73(I29dd5fb1c2673cd4daa9cafaf24d8e7c[2]);
            I2b32537c9178028493af165398a60875 = I29b4fdd4c13c96461c76660df767ea73(I29dd5fb1c2673cd4daa9cafaf24d8e7c[3]);
            If06a1563b9d7348de03a98d31bd85b06 = I29b4fdd4c13c96461c76660df767ea73(I29dd5fb1c2673cd4daa9cafaf24d8e7c[4]);
            I58a7c7b05b84d292cd06d68e96ecb9f8 = I29b4fdd4c13c96461c76660df767ea73(I29dd5fb1c2673cd4daa9cafaf24d8e7c[5]);
            I3fdec80112b3fc543b217d1c253406da = I29b4fdd4c13c96461c76660df767ea73(I29dd5fb1c2673cd4daa9cafaf24d8e7c[6]);
            Ia1aedd38250e76763aaee3de2f832b3c = I29b4fdd4c13c96461c76660df767ea73(Iead4c81d836e3befae55049797c30d6b[0]);
            I2087576fbc15119bf5d9e8afa2603b69 = I29b4fdd4c13c96461c76660df767ea73(Iead4c81d836e3befae55049797c30d6b[1]);
            I7a6ab9e700bd94208ab6528af413f3a9 = I29b4fdd4c13c96461c76660df767ea73(Iead4c81d836e3befae55049797c30d6b[2]);
            I4481555c402ba99bee05658ba6017984 = I29b4fdd4c13c96461c76660df767ea73(Iead4c81d836e3befae55049797c30d6b[3]);
            Ib849494e5087777f646ee0947b4f634a = I29b4fdd4c13c96461c76660df767ea73(Iead4c81d836e3befae55049797c30d6b[4]);
            I18d0dd7a10d6533f721a2392d4ad2d02 = I29b4fdd4c13c96461c76660df767ea73(Iead4c81d836e3befae55049797c30d6b[5]);
            Ib8603cb82ceb97c2f35bf8209306a457 = I29b4fdd4c13c96461c76660df767ea73(Iead4c81d836e3befae55049797c30d6b[6]);
            I2418ae211f327ed45cc70c42078180dc = I29b4fdd4c13c96461c76660df767ea73(Iead4c81d836e3befae55049797c30d6b[7]);
            I6521c9167261db6eb37f50b66159ddb7 = I29b4fdd4c13c96461c76660df767ea73(Iead4c81d836e3befae55049797c30d6b[8]);
            I920f95bb52cdc9b07f93afc3a6b5c009 = I29b4fdd4c13c96461c76660df767ea73(Iead4c81d836e3befae55049797c30d6b[9]);
            Iad0ecc5208263d239e4a62c5563f52ab = I29b4fdd4c13c96461c76660df767ea73(Iead4c81d836e3befae55049797c30d6b[10]);
            I0c0be3347a7df9cc39997208b013f17b = I29b4fdd4c13c96461c76660df767ea73(Iead4c81d836e3befae55049797c30d6b[11]);
            I70dc03a46e1ac0da826388abd3bdc503 = I29b4fdd4c13c96461c76660df767ea73(Iead4c81d836e3befae55049797c30d6b[12]);
            I452ba61d5fb5c7ead1824dade4bd7801 = I29b4fdd4c13c96461c76660df767ea73(I23e22f44791c167acaba27c91ef3b497[0]);
            I8b5d10c412daccdcb07645bf239d61bd = I29b4fdd4c13c96461c76660df767ea73(I23e22f44791c167acaba27c91ef3b497[1]);
            I9b1390839ee2b9ba591e3873e967c8e2 = I29b4fdd4c13c96461c76660df767ea73(I23e22f44791c167acaba27c91ef3b497[2]);
            I17e818b67440efaba9a5d19e7467bf85 = I29b4fdd4c13c96461c76660df767ea73(I23e22f44791c167acaba27c91ef3b497[3]);
            Ifa67d343acc6f3ec50c2b01fc26b4374 = I29b4fdd4c13c96461c76660df767ea73(I23e22f44791c167acaba27c91ef3b497[4]);
            If0676ef300628c4097565b13ef2d8854 = I29b4fdd4c13c96461c76660df767ea73(I23e22f44791c167acaba27c91ef3b497[5]);
            I8d26e73fafa909f1e26e329828cf4888 = I29b4fdd4c13c96461c76660df767ea73(I23e22f44791c167acaba27c91ef3b497[6]);
            If29fcea810adbdb1c4d8a4ace1d8081b = I29b4fdd4c13c96461c76660df767ea73(I23e22f44791c167acaba27c91ef3b497[7]);
            I0e3286fca6cd040758950259ab663df7 = I29b4fdd4c13c96461c76660df767ea73(I23e22f44791c167acaba27c91ef3b497[8]);
            I696db0b98e27dcc4657dc7feb23a881b = I29b4fdd4c13c96461c76660df767ea73(I23e22f44791c167acaba27c91ef3b497[9]);
            I06c0921675f464807a63c7965796f0d0 = I29b4fdd4c13c96461c76660df767ea73(I23e22f44791c167acaba27c91ef3b497[10]);
            If36016df78d833c80e1355151c038225 = I29b4fdd4c13c96461c76660df767ea73(I23e22f44791c167acaba27c91ef3b497[11]);
            I0dbf900b4f430b4c1106aa86b640bb37 = I29b4fdd4c13c96461c76660df767ea73(I23e22f44791c167acaba27c91ef3b497[12]);
            Ib8664a2abe9d6326d6e45bb2a7ad59d0 = I29b4fdd4c13c96461c76660df767ea73(Ic91f087829e0b9e0c964229a2dc567bc[0]);
            I91893028c4409cfeceeb7976815b2d31 = I29b4fdd4c13c96461c76660df767ea73(Ic91f087829e0b9e0c964229a2dc567bc[1]);
            I2e14fb1e667e967ab4c116e0c7438aec = I29b4fdd4c13c96461c76660df767ea73(Ic91f087829e0b9e0c964229a2dc567bc[2]);
            I0fb60c4f56f6d7b4007cf0dae39f4573 = I29b4fdd4c13c96461c76660df767ea73(Ic91f087829e0b9e0c964229a2dc567bc[3]);
            I24b4c998d19ae97f7178e37f75c77d06 = I29b4fdd4c13c96461c76660df767ea73(Ic91f087829e0b9e0c964229a2dc567bc[4]);
            Idb73eba1bd4ce25a6109e296f51e7dc4 = I29b4fdd4c13c96461c76660df767ea73(Ic91f087829e0b9e0c964229a2dc567bc[5]);
            Ibc1a16427d8dfa5ee20dac15327a53ea = I29b4fdd4c13c96461c76660df767ea73(Ic91f087829e0b9e0c964229a2dc567bc[6]);
            I0e52c25aa840402d944cbd81f73c1ffe = I29b4fdd4c13c96461c76660df767ea73(Ic91f087829e0b9e0c964229a2dc567bc[7]);
            Id7619819e1297844d92c8bf3a1d61926 = I29b4fdd4c13c96461c76660df767ea73(Ic91f087829e0b9e0c964229a2dc567bc[8]);
            Idfa432a87877e1ce103e56891745b62a = I29b4fdd4c13c96461c76660df767ea73(Ic91f087829e0b9e0c964229a2dc567bc[9]);
            I13b9e098622d90a1074f636d8f351aca = I29b4fdd4c13c96461c76660df767ea73(Ic91f087829e0b9e0c964229a2dc567bc[10]);
            I78e1205de9119fac3ae8f43c72ac71f4 = I29b4fdd4c13c96461c76660df767ea73(Ic91f087829e0b9e0c964229a2dc567bc[11]);
            I5bbbc4eedb7c61516769f429a8498ea7 = I29b4fdd4c13c96461c76660df767ea73(Ic91f087829e0b9e0c964229a2dc567bc[12]);
            Ia1d9dee7a9821283498d17de0cfacb32 = I29b4fdd4c13c96461c76660df767ea73(I0fd9bcdcf8faaaabf94649881419c66f[0]);
            Idd8643af2515f65fd9a1dfe66494ccf2 = I29b4fdd4c13c96461c76660df767ea73(I0fd9bcdcf8faaaabf94649881419c66f[1]);
            I1684820afb9d9cec38cfdfcd6ca8b36a = I29b4fdd4c13c96461c76660df767ea73(I0fd9bcdcf8faaaabf94649881419c66f[2]);
            Ice8a82bdd966719098a8d5f2a826f73d = I29b4fdd4c13c96461c76660df767ea73(I0fd9bcdcf8faaaabf94649881419c66f[3]);
            I338400586daa58006c0a3dcd82ea8f4a = I29b4fdd4c13c96461c76660df767ea73(I0fd9bcdcf8faaaabf94649881419c66f[4]);
            Ie467c5fde1d123da4e9587b5a56748a0 = I29b4fdd4c13c96461c76660df767ea73(I0fd9bcdcf8faaaabf94649881419c66f[5]);
            Ifc52604a4f9f9de392a35f2f9fe885b8 = I29b4fdd4c13c96461c76660df767ea73(I0fd9bcdcf8faaaabf94649881419c66f[6]);
            I20c4e393929b875521e5316f4d8e2d42 = I29b4fdd4c13c96461c76660df767ea73(I0fd9bcdcf8faaaabf94649881419c66f[7]);
            I064499f0315fbeec7b6cb50583388a07 = I29b4fdd4c13c96461c76660df767ea73(I0fd9bcdcf8faaaabf94649881419c66f[8]);
            I894ef04bfa1b7b39ef51b7c82f7686eb = I29b4fdd4c13c96461c76660df767ea73(I0fd9bcdcf8faaaabf94649881419c66f[9]);
            I8d6927b0bcbbb318cf52987c121a07b5 = I29b4fdd4c13c96461c76660df767ea73(I0fd9bcdcf8faaaabf94649881419c66f[10]);
            Ie0ce2826fd13b0e0b23c91e97787691f = I29b4fdd4c13c96461c76660df767ea73(I0fd9bcdcf8faaaabf94649881419c66f[11]);
            I7dbd1aeba00bb8b257990b7bb294211f = I29b4fdd4c13c96461c76660df767ea73(I0fd9bcdcf8faaaabf94649881419c66f[12]);
            Id5ddf5331aba567aaf5b7eb88b31a52e = I29b4fdd4c13c96461c76660df767ea73(I7cbcdd5018de9ceb49554b140e5665e8[0]);
            I0f46a17f14ab18e6338aa3d06678b0a5 = I29b4fdd4c13c96461c76660df767ea73(I7cbcdd5018de9ceb49554b140e5665e8[1]);
            If1ec4241fd12255369f72b3f3310b6e7 = I29b4fdd4c13c96461c76660df767ea73(I7cbcdd5018de9ceb49554b140e5665e8[2]);
            Iedf37dac8b3a5331277ae4f0176968aa = I29b4fdd4c13c96461c76660df767ea73(I7cbcdd5018de9ceb49554b140e5665e8[3]);
            Ia422fbdf8f318ff3ddc049d1374e7939 = I29b4fdd4c13c96461c76660df767ea73(I7cbcdd5018de9ceb49554b140e5665e8[4]);
            I9cbe73d708c561d43d05945552d32dde = I29b4fdd4c13c96461c76660df767ea73(I7cbcdd5018de9ceb49554b140e5665e8[5]);
            I7e36dcae438a712fca2320117b7e3356 = I29b4fdd4c13c96461c76660df767ea73(I5a79c19fd2093d974b574e85245b5617[0]);
            I0f9bc36c9d40290f83489aac3d674924 = I29b4fdd4c13c96461c76660df767ea73(I5a79c19fd2093d974b574e85245b5617[1]);
            I3a09554ca009781e28ef1b3ea70d39ad = I29b4fdd4c13c96461c76660df767ea73(I5a79c19fd2093d974b574e85245b5617[2]);
            I28ea268c5b51ac1d9249e96599bb6b0d = I29b4fdd4c13c96461c76660df767ea73(I5a79c19fd2093d974b574e85245b5617[3]);
            I1d648ed8f07f0743a6d616584270c513 = I29b4fdd4c13c96461c76660df767ea73(I5a79c19fd2093d974b574e85245b5617[4]);
            I82a225237aeb1ceb31e8cd18b1e45c6f = I29b4fdd4c13c96461c76660df767ea73(I5a79c19fd2093d974b574e85245b5617[5]);
            I36ed1a0d0d618f90443fbea17b7c97ec = I29b4fdd4c13c96461c76660df767ea73(Ica937143b618734fa099683949153130[0]);
            I612a41511db375f10f3c2b10d13edb24 = I29b4fdd4c13c96461c76660df767ea73(Ica937143b618734fa099683949153130[1]);
            I19032091a26dfdfffff60818041ec79e = I29b4fdd4c13c96461c76660df767ea73(Ica937143b618734fa099683949153130[2]);
            I6aba8ca0e4b20a6355b43a70f19d9d8c = I29b4fdd4c13c96461c76660df767ea73(Ica937143b618734fa099683949153130[3]);
            I839895c8614ff28df83314c44824900b = I29b4fdd4c13c96461c76660df767ea73(Ica937143b618734fa099683949153130[4]);
            I8cbafa797ef136d7e50c909dc160deb1 = I29b4fdd4c13c96461c76660df767ea73(Ica937143b618734fa099683949153130[5]);
            Ibac0851ce1a3c23f18b072d263afff36 = I29b4fdd4c13c96461c76660df767ea73(I2d4d5d2694718b39e80b89b422d690cc[0]);
            Id58474582f209a3859f65a447fe99191 = I29b4fdd4c13c96461c76660df767ea73(I2d4d5d2694718b39e80b89b422d690cc[1]);
            Ic9e06a355beabfacc053ec48f17f49de = I29b4fdd4c13c96461c76660df767ea73(I2d4d5d2694718b39e80b89b422d690cc[2]);
            I77fd8001d879fc9e9117464fba27902d = I29b4fdd4c13c96461c76660df767ea73(I2d4d5d2694718b39e80b89b422d690cc[3]);
            I2a0dc4ed573a544cb13544e049514903 = I29b4fdd4c13c96461c76660df767ea73(I2d4d5d2694718b39e80b89b422d690cc[4]);
            I71bc7271cc432bb3c5d0b7a416cdfc60 = I29b4fdd4c13c96461c76660df767ea73(I2d4d5d2694718b39e80b89b422d690cc[5]);
            Ib76e892d1a1271844338042381b5690b = I29b4fdd4c13c96461c76660df767ea73(Ic2faea3d4bb97dda16ecc29c27939ca6[0]);
            Icb158c031d434cb419c15e0510511231 = I29b4fdd4c13c96461c76660df767ea73(Ic2faea3d4bb97dda16ecc29c27939ca6[1]);
            I563802213afb6abe2f6e8c6f4d1e5b08 = I29b4fdd4c13c96461c76660df767ea73(Ic2faea3d4bb97dda16ecc29c27939ca6[2]);
            Ia5b779ef95333736b08f63770900e275 = I29b4fdd4c13c96461c76660df767ea73(Ic2faea3d4bb97dda16ecc29c27939ca6[3]);
            Ic1120eb027841908cd64fe5c7274da14 = I29b4fdd4c13c96461c76660df767ea73(Ic2faea3d4bb97dda16ecc29c27939ca6[4]);
            I5160de2c5ce4782d8f8be10dc740694b = I29b4fdd4c13c96461c76660df767ea73(Ic2faea3d4bb97dda16ecc29c27939ca6[5]);
            I5f7b6e6a30348ae86057f7e56f625846 = I29b4fdd4c13c96461c76660df767ea73(Ic2faea3d4bb97dda16ecc29c27939ca6[6]);
            I9de41d0b279b84366640880dbd18c502 = I29b4fdd4c13c96461c76660df767ea73(Ic2faea3d4bb97dda16ecc29c27939ca6[7]);
            Ifec9abca21cf476b70e0befa3926b46a = I29b4fdd4c13c96461c76660df767ea73(I503e83a1146c42d5c1ef011ecb280807[0]);
            Ifc527b6af9486df7f52d7eb9637c671f = I29b4fdd4c13c96461c76660df767ea73(I503e83a1146c42d5c1ef011ecb280807[1]);
            I31d94aae2e3721045fe850d84dd2225a = I29b4fdd4c13c96461c76660df767ea73(I503e83a1146c42d5c1ef011ecb280807[2]);
            If3bdbb4c20efca0c5af78614b4271ed1 = I29b4fdd4c13c96461c76660df767ea73(I503e83a1146c42d5c1ef011ecb280807[3]);
            I4037f1b207aa101f354e59eddd7c9eb4 = I29b4fdd4c13c96461c76660df767ea73(I503e83a1146c42d5c1ef011ecb280807[4]);
            If4d63635a5f99c4dc9e5b57712830c20 = I29b4fdd4c13c96461c76660df767ea73(I503e83a1146c42d5c1ef011ecb280807[5]);
            I1f1f2fefd3381ee48ab0ec9c9301754b = I29b4fdd4c13c96461c76660df767ea73(I503e83a1146c42d5c1ef011ecb280807[6]);
            Iba52b84e6e215842e0ca8e72c42ebce7 = I29b4fdd4c13c96461c76660df767ea73(I503e83a1146c42d5c1ef011ecb280807[7]);
            I597c3f5c14e235f90dc8c796bc3e931d = I29b4fdd4c13c96461c76660df767ea73(Ib9886c1fcd27ceb24afb2d0d7da85c26[0]);
            I397a69dab323c7148b620dd6fe0b0c51 = I29b4fdd4c13c96461c76660df767ea73(Ib9886c1fcd27ceb24afb2d0d7da85c26[1]);
            I401ab1ad994f5018061a3f57d3a51ad1 = I29b4fdd4c13c96461c76660df767ea73(Ib9886c1fcd27ceb24afb2d0d7da85c26[2]);
            I3a47540f34ce47bcfa1da66cc4e6e088 = I29b4fdd4c13c96461c76660df767ea73(Ib9886c1fcd27ceb24afb2d0d7da85c26[3]);
            I18916d0023ca275d84c52af07dcc5ca2 = I29b4fdd4c13c96461c76660df767ea73(Ib9886c1fcd27ceb24afb2d0d7da85c26[4]);
            Ic79072d9e42dbc9974231f1d642b3f12 = I29b4fdd4c13c96461c76660df767ea73(Ib9886c1fcd27ceb24afb2d0d7da85c26[5]);
            I1140fa91b5e22ba0c094c03295781e5a = I29b4fdd4c13c96461c76660df767ea73(Ib9886c1fcd27ceb24afb2d0d7da85c26[6]);
            Id2989aaee3930698cd374e6c9feedf82 = I29b4fdd4c13c96461c76660df767ea73(Ib9886c1fcd27ceb24afb2d0d7da85c26[7]);
            Icda9a86a25dbe516a93b46fe487029e3 = I29b4fdd4c13c96461c76660df767ea73(Icd90612c09423a2817a72f750e585309[0]);
            I53971b75cbd7ebc74b579776a6ea4778 = I29b4fdd4c13c96461c76660df767ea73(Icd90612c09423a2817a72f750e585309[1]);
            I37e5c3118e8536e37bd797aeaa92476c = I29b4fdd4c13c96461c76660df767ea73(Icd90612c09423a2817a72f750e585309[2]);
            I9c68bfa3b888b6a6d41e38e674578284 = I29b4fdd4c13c96461c76660df767ea73(Icd90612c09423a2817a72f750e585309[3]);
            I2c72d6c5fa6968dffa6517cf81219875 = I29b4fdd4c13c96461c76660df767ea73(Icd90612c09423a2817a72f750e585309[4]);
            I9bb4d58b1fe80549451b00c4ed2b3885 = I29b4fdd4c13c96461c76660df767ea73(Icd90612c09423a2817a72f750e585309[5]);
            Ic488e78b5c73251b673301e84c4b5b0b = I29b4fdd4c13c96461c76660df767ea73(Icd90612c09423a2817a72f750e585309[6]);
            I8d07beccef519ab4ce4024d911ac2346 = I29b4fdd4c13c96461c76660df767ea73(Icd90612c09423a2817a72f750e585309[7]);
            I7c191c2c2be09886d0f31e4368797afd = I29b4fdd4c13c96461c76660df767ea73(Ib7b7884d2653893806af34579f7c0760[0]);
            Ia3bfd86e26efbef2cf6bb72be7ac1453 = I29b4fdd4c13c96461c76660df767ea73(Ib7b7884d2653893806af34579f7c0760[1]);
            I4ae59dd2f57bda295e11b077e8668f1a = I29b4fdd4c13c96461c76660df767ea73(Ib7b7884d2653893806af34579f7c0760[2]);
            I3f6fad8bb0fba790fcdb1612b6fa7712 = I29b4fdd4c13c96461c76660df767ea73(Ib7b7884d2653893806af34579f7c0760[3]);
            I58416287b268462d28f55c6c2705e613 = I29b4fdd4c13c96461c76660df767ea73(Ib7b7884d2653893806af34579f7c0760[4]);
            I106d0e71b7378d110b0a624e5cbf0d6e = I29b4fdd4c13c96461c76660df767ea73(Ib7b7884d2653893806af34579f7c0760[5]);
            I59adad4fd84c1fc233dc58f70a12779d = I29b4fdd4c13c96461c76660df767ea73(Ib7b7884d2653893806af34579f7c0760[6]);
            I8e01532a1ab9534b8de0474549d41a2e = I29b4fdd4c13c96461c76660df767ea73(Ib7b7884d2653893806af34579f7c0760[7]);
            I80af3dcb716f3474a7257700aef89b81 = I29b4fdd4c13c96461c76660df767ea73(Ib7b7884d2653893806af34579f7c0760[8]);
            I07d68462362d8453e83570cc793c55db = I29b4fdd4c13c96461c76660df767ea73(Ic3f0ad21d8a446c31afec49309a18133[0]);
            I9a2bba3f62de5f750dc8161a488dc331 = I29b4fdd4c13c96461c76660df767ea73(Ic3f0ad21d8a446c31afec49309a18133[1]);
            I71da7e172b2b967040b6e6d02ef9949e = I29b4fdd4c13c96461c76660df767ea73(Ic3f0ad21d8a446c31afec49309a18133[2]);
            Ib97b2670a6cd88b2327f07f62d887900 = I29b4fdd4c13c96461c76660df767ea73(Ic3f0ad21d8a446c31afec49309a18133[3]);
            Ib2963b82260024e1853d297798d88d3c = I29b4fdd4c13c96461c76660df767ea73(Ic3f0ad21d8a446c31afec49309a18133[4]);
            I0722ec4e9d400f8eaeacd060e42de79c = I29b4fdd4c13c96461c76660df767ea73(Ic3f0ad21d8a446c31afec49309a18133[5]);
            I1972375d51767f0cffa5395a354b3493 = I29b4fdd4c13c96461c76660df767ea73(Ic3f0ad21d8a446c31afec49309a18133[6]);
            Ifb19d75cfa0051107b5fba57bfc002b5 = I29b4fdd4c13c96461c76660df767ea73(Ic3f0ad21d8a446c31afec49309a18133[7]);
            I9d05dc0e39e85c23b62f343a8de12e64 = I29b4fdd4c13c96461c76660df767ea73(Ic3f0ad21d8a446c31afec49309a18133[8]);
            I64ae3cd6f36b8bde29cd3e1fcba7bade = I29b4fdd4c13c96461c76660df767ea73(I2dd65bec7d2bc4778b7fc48a413d2ba7[0]);
            Ia6a78664c080829664158f53ba330312 = I29b4fdd4c13c96461c76660df767ea73(I2dd65bec7d2bc4778b7fc48a413d2ba7[1]);
            I2ba16a10a82c20d54c776a9804ee50e4 = I29b4fdd4c13c96461c76660df767ea73(I2dd65bec7d2bc4778b7fc48a413d2ba7[2]);
            Ie9a316de516ec4fb828a614c67e38b2a = I29b4fdd4c13c96461c76660df767ea73(I2dd65bec7d2bc4778b7fc48a413d2ba7[3]);
            Ie945349d77442536992d9ad52ce84218 = I29b4fdd4c13c96461c76660df767ea73(I2dd65bec7d2bc4778b7fc48a413d2ba7[4]);
            Ic6a7a82d16e6106071934ba79d3698cd = I29b4fdd4c13c96461c76660df767ea73(I2dd65bec7d2bc4778b7fc48a413d2ba7[5]);
            Ide40b1bf9c0b642c49a5685a62af1c93 = I29b4fdd4c13c96461c76660df767ea73(I2dd65bec7d2bc4778b7fc48a413d2ba7[6]);
            I79280400a4c9bed015106e5d006de757 = I29b4fdd4c13c96461c76660df767ea73(I2dd65bec7d2bc4778b7fc48a413d2ba7[7]);
            Ic6e3847f035738243f4c5f71f296da57 = I29b4fdd4c13c96461c76660df767ea73(I2dd65bec7d2bc4778b7fc48a413d2ba7[8]);
            I45b64b2b963963d2d0a8318133941f1d = I29b4fdd4c13c96461c76660df767ea73(I36b5867a3da6f2ed529e791166640d3f[0]);
            I1939152ddbede923cde577984e0aa743 = I29b4fdd4c13c96461c76660df767ea73(I36b5867a3da6f2ed529e791166640d3f[1]);
            Ifbcebda2bb0ce58a0e1764c392a816df = I29b4fdd4c13c96461c76660df767ea73(I36b5867a3da6f2ed529e791166640d3f[2]);
            I6d0d098e6d47dea04d6d7be67b648a0d = I29b4fdd4c13c96461c76660df767ea73(I36b5867a3da6f2ed529e791166640d3f[3]);
            Icaeb9a2ec8ec5822658fa85b88cca04b = I29b4fdd4c13c96461c76660df767ea73(I36b5867a3da6f2ed529e791166640d3f[4]);
            I3cc30aaba3dcd3eda262a19e85e53117 = I29b4fdd4c13c96461c76660df767ea73(I36b5867a3da6f2ed529e791166640d3f[5]);
            Ic0b2f9717b8aacb34325fd5aaf03a366 = I29b4fdd4c13c96461c76660df767ea73(I36b5867a3da6f2ed529e791166640d3f[6]);
            I002869e450d79649d27441ce00bfb575 = I29b4fdd4c13c96461c76660df767ea73(I36b5867a3da6f2ed529e791166640d3f[7]);
            Ie4d20df6b1e7a42f0df9a3cc26b12ac1 = I29b4fdd4c13c96461c76660df767ea73(I36b5867a3da6f2ed529e791166640d3f[8]);
            Idd01d014f0469f893305057ae3f4cb2e = I29b4fdd4c13c96461c76660df767ea73(Iedc20522d3322bbe3f55e2aa611d76df[0]);
            I79444eef1875b6ad1a0675b66392ff9d = I29b4fdd4c13c96461c76660df767ea73(Iedc20522d3322bbe3f55e2aa611d76df[1]);
            I7caf8c7496dd96c1ed08e98b415f5775 = I29b4fdd4c13c96461c76660df767ea73(Iedc20522d3322bbe3f55e2aa611d76df[2]);
            I7fc6e2aecff5bd691872d1e10a39103b = I29b4fdd4c13c96461c76660df767ea73(Iedc20522d3322bbe3f55e2aa611d76df[3]);
            I49321308413cb4dbe5e6c01ba5b9023c = I29b4fdd4c13c96461c76660df767ea73(Iedc20522d3322bbe3f55e2aa611d76df[4]);
            Id27560fb44b4f2fda98d47e9f20d6898 = I29b4fdd4c13c96461c76660df767ea73(Iedc20522d3322bbe3f55e2aa611d76df[5]);
            I745187336b8a5ae4eac66e90539752cf = I29b4fdd4c13c96461c76660df767ea73(Iedc20522d3322bbe3f55e2aa611d76df[6]);
            I772e844c41387e7079259875e0ba3fa0 = I29b4fdd4c13c96461c76660df767ea73(Iedc20522d3322bbe3f55e2aa611d76df[7]);
            I32c35da92922c5b477f8aba837fa6d92 = I29b4fdd4c13c96461c76660df767ea73(Iedc20522d3322bbe3f55e2aa611d76df[8]);
            I3bc01b072987a0c980615abbc2251e5f = I29b4fdd4c13c96461c76660df767ea73(Iedc20522d3322bbe3f55e2aa611d76df[9]);
            If08adda7d796da7c7849e472a73282a3 = I29b4fdd4c13c96461c76660df767ea73(Iedc20522d3322bbe3f55e2aa611d76df[10]);
            Ife3bb8945e14d8746c82b66886293997 = I29b4fdd4c13c96461c76660df767ea73(Iedc20522d3322bbe3f55e2aa611d76df[11]);
            I45ef0ac486fe043f57e8a46aa91461a3 = I29b4fdd4c13c96461c76660df767ea73(Iedc20522d3322bbe3f55e2aa611d76df[12]);
            Ic0ae1191869e636f9e4391efe93309ae = I29b4fdd4c13c96461c76660df767ea73(Iedc20522d3322bbe3f55e2aa611d76df[13]);
            Id92d779518ae724b5fef5221372f8f26 = I29b4fdd4c13c96461c76660df767ea73(Iedc20522d3322bbe3f55e2aa611d76df[14]);
            Id0762ac7710c93249bc11c6ce4ae51a0 = I29b4fdd4c13c96461c76660df767ea73(Iedc20522d3322bbe3f55e2aa611d76df[15]);
            Ife6be241bc50560a14f97650e5cc2959 = I29b4fdd4c13c96461c76660df767ea73(I6821e897aea31f7c237ca1a553bf0cd1[0]);
            I1062442edb2bff727ca6283c8270bf28 = I29b4fdd4c13c96461c76660df767ea73(I6821e897aea31f7c237ca1a553bf0cd1[1]);
            I6c9ae8b8191507f908c27bbde53bf2d5 = I29b4fdd4c13c96461c76660df767ea73(I6821e897aea31f7c237ca1a553bf0cd1[2]);
            Iec936eeebd1f8c95307bd8705e6def81 = I29b4fdd4c13c96461c76660df767ea73(I6821e897aea31f7c237ca1a553bf0cd1[3]);
            I6332af145d560e3f22a4a88106749f98 = I29b4fdd4c13c96461c76660df767ea73(I6821e897aea31f7c237ca1a553bf0cd1[4]);
            I0c121fa3e9e6e0e2e8291a594d6b4ceb = I29b4fdd4c13c96461c76660df767ea73(I6821e897aea31f7c237ca1a553bf0cd1[5]);
            Ic3c59a5167cb83fd76ec6236572b1f3d = I29b4fdd4c13c96461c76660df767ea73(I6821e897aea31f7c237ca1a553bf0cd1[6]);
            I3e8e280553edaa5c8555ace81ecc10e0 = I29b4fdd4c13c96461c76660df767ea73(I6821e897aea31f7c237ca1a553bf0cd1[7]);
            I3e466d40a4447a23953d96d2e6d61d47 = I29b4fdd4c13c96461c76660df767ea73(I6821e897aea31f7c237ca1a553bf0cd1[8]);
            I76e4c55148effeba62a4837cd19c5e51 = I29b4fdd4c13c96461c76660df767ea73(I6821e897aea31f7c237ca1a553bf0cd1[9]);
            Ie335e68643fd2b0a53351f4bd45c3475 = I29b4fdd4c13c96461c76660df767ea73(I6821e897aea31f7c237ca1a553bf0cd1[10]);
            I89f75107ea95f207b9e664a1f4f0746a = I29b4fdd4c13c96461c76660df767ea73(I6821e897aea31f7c237ca1a553bf0cd1[11]);
            Ic8f0049e1298b14b4e039075dc0d5f74 = I29b4fdd4c13c96461c76660df767ea73(I6821e897aea31f7c237ca1a553bf0cd1[12]);
            I382153cec6f7d6258574e7c532186473 = I29b4fdd4c13c96461c76660df767ea73(I6821e897aea31f7c237ca1a553bf0cd1[13]);
            I351dc309e916f282cc1e19303eee4112 = I29b4fdd4c13c96461c76660df767ea73(I6821e897aea31f7c237ca1a553bf0cd1[14]);
            I9de5e90485b3f22e9003dc8a7b22a79b = I29b4fdd4c13c96461c76660df767ea73(I6821e897aea31f7c237ca1a553bf0cd1[15]);
            Idc4171a40dd2470e852af37a461013c7 = I29b4fdd4c13c96461c76660df767ea73(I290499340d94dd8e234f53f9962a182b[0]);
            Ifae488cb68d95ea517376319eb11f1bf = I29b4fdd4c13c96461c76660df767ea73(I290499340d94dd8e234f53f9962a182b[1]);
            I9cab38b69794ab661e12750cf69c822c = I29b4fdd4c13c96461c76660df767ea73(I290499340d94dd8e234f53f9962a182b[2]);
            I24180fba17c21bacefa8a4514e4b685c = I29b4fdd4c13c96461c76660df767ea73(I290499340d94dd8e234f53f9962a182b[3]);
            I83bbe6fa947f9f909e1a6785ab31901f = I29b4fdd4c13c96461c76660df767ea73(I290499340d94dd8e234f53f9962a182b[4]);
            I202c385beeccee309104b66f8f096b2c = I29b4fdd4c13c96461c76660df767ea73(I290499340d94dd8e234f53f9962a182b[5]);
            Idc549661d6694035874a3366704801c7 = I29b4fdd4c13c96461c76660df767ea73(I290499340d94dd8e234f53f9962a182b[6]);
            I778fbaea65beeb6de599490daf3b7e3c = I29b4fdd4c13c96461c76660df767ea73(I290499340d94dd8e234f53f9962a182b[7]);
            I4fd45670f88265e5d7aa6582f3ad3ff8 = I29b4fdd4c13c96461c76660df767ea73(I290499340d94dd8e234f53f9962a182b[8]);
            I2d636a246d815a4d12c478794860dd40 = I29b4fdd4c13c96461c76660df767ea73(I290499340d94dd8e234f53f9962a182b[9]);
            I3319313fe1d2b4ec2626711b187b4a5a = I29b4fdd4c13c96461c76660df767ea73(I290499340d94dd8e234f53f9962a182b[10]);
            I586aaa5c55efd37996b01febd3bc60a4 = I29b4fdd4c13c96461c76660df767ea73(I290499340d94dd8e234f53f9962a182b[11]);
            I95ccc219b5f5038641b38dff6db0b222 = I29b4fdd4c13c96461c76660df767ea73(I290499340d94dd8e234f53f9962a182b[12]);
            I5001118df37d08bd19d322aca8ff3996 = I29b4fdd4c13c96461c76660df767ea73(I290499340d94dd8e234f53f9962a182b[13]);
            I22c15857572603cc24d8a87cb47c33b0 = I29b4fdd4c13c96461c76660df767ea73(I290499340d94dd8e234f53f9962a182b[14]);
            Ifdcd91f925b63e0817798aa6e9200e50 = I29b4fdd4c13c96461c76660df767ea73(I290499340d94dd8e234f53f9962a182b[15]);
            I8435e69bc1ff06e7edfabbee7b9aa49e = I29b4fdd4c13c96461c76660df767ea73(I5ce387684404cf922955e4af33ed2367[0]);
            Ibeff607ba15fd8ef504224a9c1d102fc = I29b4fdd4c13c96461c76660df767ea73(I5ce387684404cf922955e4af33ed2367[1]);
            Id15c3bdce785df234c68432ccec8f959 = I29b4fdd4c13c96461c76660df767ea73(I5ce387684404cf922955e4af33ed2367[2]);
            I25888aa2135fc403ca9eac4df634549a = I29b4fdd4c13c96461c76660df767ea73(I5ce387684404cf922955e4af33ed2367[3]);
            I632ffd09a9091335b3aa91ab2a8f1cce = I29b4fdd4c13c96461c76660df767ea73(I5ce387684404cf922955e4af33ed2367[4]);
            I283331db80e6d0891b13dc55e6a7d76c = I29b4fdd4c13c96461c76660df767ea73(I5ce387684404cf922955e4af33ed2367[5]);
            I134a734d93e62f6ac6635015fe3a2096 = I29b4fdd4c13c96461c76660df767ea73(I5ce387684404cf922955e4af33ed2367[6]);
            Id66798f8ea67e74a67f264fe6b4503a3 = I29b4fdd4c13c96461c76660df767ea73(I5ce387684404cf922955e4af33ed2367[7]);
            If2ce7b8d2573494564393f7d426fa47f = I29b4fdd4c13c96461c76660df767ea73(I5ce387684404cf922955e4af33ed2367[8]);
            Id59cf860d9f4aff11b205b8970d93df3 = I29b4fdd4c13c96461c76660df767ea73(I5ce387684404cf922955e4af33ed2367[9]);
            I75aaeab4f372e28a8e51453540f9c6b2 = I29b4fdd4c13c96461c76660df767ea73(I5ce387684404cf922955e4af33ed2367[10]);
            I2266afbacf1ba750ce18f296aba1181d = I29b4fdd4c13c96461c76660df767ea73(I5ce387684404cf922955e4af33ed2367[11]);
            I69c2b063e61e14f5d49b907095ece00f = I29b4fdd4c13c96461c76660df767ea73(I5ce387684404cf922955e4af33ed2367[12]);
            If077c67a062095cfe69f2260cee82833 = I29b4fdd4c13c96461c76660df767ea73(I5ce387684404cf922955e4af33ed2367[13]);
            Ibc03a9b6115d0941ce9233df7ef2fa57 = I29b4fdd4c13c96461c76660df767ea73(I5ce387684404cf922955e4af33ed2367[14]);
            Ia18bdb8d2f02b50281f0acd4a45ac973 = I29b4fdd4c13c96461c76660df767ea73(I5ce387684404cf922955e4af33ed2367[15]);
            Ib88c884e54d6e6ecf5ac015bc304e4f3 = I29b4fdd4c13c96461c76660df767ea73(I1ae87f851f8bd64e6e1428a143e82151[0]);
            If6f5efee5e1f9709d86bf28cfb741955 = I29b4fdd4c13c96461c76660df767ea73(I1ae87f851f8bd64e6e1428a143e82151[1]);
            Ia0caf6693d441ac622f416a86b665166 = I29b4fdd4c13c96461c76660df767ea73(I1ae87f851f8bd64e6e1428a143e82151[2]);
            I85dd6a9634284c22027b4241551ea628 = I29b4fdd4c13c96461c76660df767ea73(I1ae87f851f8bd64e6e1428a143e82151[3]);
            Id5cedaa397ebfc2567efcc2f8a648db5 = I29b4fdd4c13c96461c76660df767ea73(I1ae87f851f8bd64e6e1428a143e82151[4]);
            Ica0a119af1728ae253c16cc3eb93f802 = I29b4fdd4c13c96461c76660df767ea73(I1ae87f851f8bd64e6e1428a143e82151[5]);
            Ie7274a7ffa053ced4f12a67986d3c81b = I29b4fdd4c13c96461c76660df767ea73(I1ae87f851f8bd64e6e1428a143e82151[6]);
            Ife7985db888089ea618413810611bfca = I29b4fdd4c13c96461c76660df767ea73(I1ae87f851f8bd64e6e1428a143e82151[7]);
            If49068db99aa9d09302eda27ab51fcb7 = I29b4fdd4c13c96461c76660df767ea73(I1ae87f851f8bd64e6e1428a143e82151[8]);
            I2959f2dc554e599d675eb6912757e413 = I29b4fdd4c13c96461c76660df767ea73(I646767a2d4b3029ed7acb73a15af1682[0]);
            I898d1b59aab3d5d4adce8ec3c0e14a0d = I29b4fdd4c13c96461c76660df767ea73(I646767a2d4b3029ed7acb73a15af1682[1]);
            Ibb6e54edb9d277242c06d386a9a75a26 = I29b4fdd4c13c96461c76660df767ea73(I646767a2d4b3029ed7acb73a15af1682[2]);
            I51b1cd475d0e389326b182cbe680a402 = I29b4fdd4c13c96461c76660df767ea73(I646767a2d4b3029ed7acb73a15af1682[3]);
            If12366160fdc899bd71cb0de5bcfd84d = I29b4fdd4c13c96461c76660df767ea73(I646767a2d4b3029ed7acb73a15af1682[4]);
            I44e5ce0cdf812c5b73e6e638da36e414 = I29b4fdd4c13c96461c76660df767ea73(I646767a2d4b3029ed7acb73a15af1682[5]);
            I4f38c3d620b72f21cf6d54c7df4ba816 = I29b4fdd4c13c96461c76660df767ea73(I646767a2d4b3029ed7acb73a15af1682[6]);
            Ib66b897398ea0702b74bdd03774f3ae4 = I29b4fdd4c13c96461c76660df767ea73(I646767a2d4b3029ed7acb73a15af1682[7]);
            I0b3a936c3f7e0391111e696b2445803b = I29b4fdd4c13c96461c76660df767ea73(I646767a2d4b3029ed7acb73a15af1682[8]);
            I10f045edf47784a91a5599494c2d3de2 = I29b4fdd4c13c96461c76660df767ea73(I48001f5c6554999a2178308ae271b70e[0]);
            I6a81b4485598387e4656c35e83866209 = I29b4fdd4c13c96461c76660df767ea73(I48001f5c6554999a2178308ae271b70e[1]);
            Icf7630b6002db2f9b59d5323d6cc8105 = I29b4fdd4c13c96461c76660df767ea73(I48001f5c6554999a2178308ae271b70e[2]);
            I3db0adb3457cb22c755f5d29a8fe7ed8 = I29b4fdd4c13c96461c76660df767ea73(I48001f5c6554999a2178308ae271b70e[3]);
            I887911fd9466f4d4fa7f50642d610d88 = I29b4fdd4c13c96461c76660df767ea73(I48001f5c6554999a2178308ae271b70e[4]);
            I9ae284c0089ae462a1bb9d168bde2fd0 = I29b4fdd4c13c96461c76660df767ea73(I48001f5c6554999a2178308ae271b70e[5]);
            I342a563de39175fe4a6eb7e3e1ccac9a = I29b4fdd4c13c96461c76660df767ea73(I48001f5c6554999a2178308ae271b70e[6]);
            Idc758f8e6fabb6b31b0a7d9c0c590310 = I29b4fdd4c13c96461c76660df767ea73(I48001f5c6554999a2178308ae271b70e[7]);
            I72b4ef48363856af7faacc85eafbaf2f = I29b4fdd4c13c96461c76660df767ea73(I48001f5c6554999a2178308ae271b70e[8]);
            I4ae2f2330a8ee7d5626499f2a030c7a5 = I29b4fdd4c13c96461c76660df767ea73(I7fe6d853fc1c11142b64ff8f40783246[0]);
            I4aa98503fc71292d42dba1cab6db952f = I29b4fdd4c13c96461c76660df767ea73(I7fe6d853fc1c11142b64ff8f40783246[1]);
            Ic35d5ac4dac46d47b2796bbac6452161 = I29b4fdd4c13c96461c76660df767ea73(I7fe6d853fc1c11142b64ff8f40783246[2]);
            I32679702c19eab37b46d13bb372967ea = I29b4fdd4c13c96461c76660df767ea73(I7fe6d853fc1c11142b64ff8f40783246[3]);
            I6a86b03402bd2e35208d3fc74601f9cf = I29b4fdd4c13c96461c76660df767ea73(I7fe6d853fc1c11142b64ff8f40783246[4]);
            If8a259e0c4f1839e852abec6e1b904ee = I29b4fdd4c13c96461c76660df767ea73(I7fe6d853fc1c11142b64ff8f40783246[5]);
            I938dd59e4cdf3434086f60d000113430 = I29b4fdd4c13c96461c76660df767ea73(I7fe6d853fc1c11142b64ff8f40783246[6]);
            Idc198bd5732ca5760d1a700a25273ce3 = I29b4fdd4c13c96461c76660df767ea73(I7fe6d853fc1c11142b64ff8f40783246[7]);
            I9dfdffbfdb83572cc3205f674e5db753 = I29b4fdd4c13c96461c76660df767ea73(I7fe6d853fc1c11142b64ff8f40783246[8]);
            I60520c850a95b893528569c4069bd677 = I29b4fdd4c13c96461c76660df767ea73(Iadc98deb917f599574e99a90e3230e88[0]);
            If525ac3dc97e3187e036d70e9984939d = I29b4fdd4c13c96461c76660df767ea73(Iadc98deb917f599574e99a90e3230e88[1]);
            I0c1e4d400520935c5c78b792a9d554ba = I29b4fdd4c13c96461c76660df767ea73(Iadc98deb917f599574e99a90e3230e88[2]);
            Ic7d5fe6c4b1dcb97d10ba3de2f95d1df = I29b4fdd4c13c96461c76660df767ea73(Iadc98deb917f599574e99a90e3230e88[3]);
            I8efad9622c05177563ab8a2747879044 = I29b4fdd4c13c96461c76660df767ea73(Iadc98deb917f599574e99a90e3230e88[4]);
            Ied4ddedaf801fbd7238d8a55c17c8090 = I29b4fdd4c13c96461c76660df767ea73(Iadc98deb917f599574e99a90e3230e88[5]);
            Ieb9720b6beb2363d651346ef0233cd49 = I29b4fdd4c13c96461c76660df767ea73(Iadc98deb917f599574e99a90e3230e88[6]);
            I202aa0814e7e28a6bd21db116b652b4d = I29b4fdd4c13c96461c76660df767ea73(Iadc98deb917f599574e99a90e3230e88[7]);
            Id201f81bbd80a70006a10866b8efeeff = I29b4fdd4c13c96461c76660df767ea73(Iadc98deb917f599574e99a90e3230e88[8]);
            Ic227f42a20219c6638ee3343ca445acf = I29b4fdd4c13c96461c76660df767ea73(Iadc98deb917f599574e99a90e3230e88[9]);
            I507e9bd0265d9ca6cd21a46fa21ba084 = I29b4fdd4c13c96461c76660df767ea73(Iadc98deb917f599574e99a90e3230e88[10]);
            Ie04e44d8e0756cdf34cf9ad53da76e47 = I29b4fdd4c13c96461c76660df767ea73(Iadc98deb917f599574e99a90e3230e88[11]);
            Ic92ab3dac1a151d6ff0b4e0c21003eb0 = I29b4fdd4c13c96461c76660df767ea73(I3d79461a85cd6a58bf9f96f6e0d704ac[0]);
            I3da241c7f221413abfbf1b4384bfca5a = I29b4fdd4c13c96461c76660df767ea73(I3d79461a85cd6a58bf9f96f6e0d704ac[1]);
            I0807a826e91f92ef279ccf0b6512a428 = I29b4fdd4c13c96461c76660df767ea73(I3d79461a85cd6a58bf9f96f6e0d704ac[2]);
            I05aabdf73200996b7bea8db700fa8930 = I29b4fdd4c13c96461c76660df767ea73(I3d79461a85cd6a58bf9f96f6e0d704ac[3]);
            I03038b940be8bd21bd26b150b28754a6 = I29b4fdd4c13c96461c76660df767ea73(I3d79461a85cd6a58bf9f96f6e0d704ac[4]);
            Ibf547f8a5e1059ffaabeb3f447904dcf = I29b4fdd4c13c96461c76660df767ea73(I3d79461a85cd6a58bf9f96f6e0d704ac[5]);
            I2ea27544ba4cc14d0f7ccf7158a27a2f = I29b4fdd4c13c96461c76660df767ea73(I3d79461a85cd6a58bf9f96f6e0d704ac[6]);
            Ib2f34922b0d5346500de093275bebc94 = I29b4fdd4c13c96461c76660df767ea73(I3d79461a85cd6a58bf9f96f6e0d704ac[7]);
            Id2e223005a932987b6f60663773187f8 = I29b4fdd4c13c96461c76660df767ea73(I3d79461a85cd6a58bf9f96f6e0d704ac[8]);
            I3188d354c2ba494ffe210dcd89c00620 = I29b4fdd4c13c96461c76660df767ea73(I3d79461a85cd6a58bf9f96f6e0d704ac[9]);
            I09faa07bf38acd96c4e29afd8a5167e8 = I29b4fdd4c13c96461c76660df767ea73(I3d79461a85cd6a58bf9f96f6e0d704ac[10]);
            I6d4867d03d9187e95e27e99f7aecddec = I29b4fdd4c13c96461c76660df767ea73(I3d79461a85cd6a58bf9f96f6e0d704ac[11]);
            Ifb09b84f9681c7bc28ffd562b633ffd9 = I29b4fdd4c13c96461c76660df767ea73(I2fcbccd884710be9c6a34f78d2ae6a18[0]);
            Ib55b0e4c45ebbdb605f0ba9d62bff21c = I29b4fdd4c13c96461c76660df767ea73(I2fcbccd884710be9c6a34f78d2ae6a18[1]);
            I4319fa23d59f4e690e31fb7e3a823d17 = I29b4fdd4c13c96461c76660df767ea73(I2fcbccd884710be9c6a34f78d2ae6a18[2]);
            I4ee3f608cc8f8df27345949f1a3713a7 = I29b4fdd4c13c96461c76660df767ea73(I2fcbccd884710be9c6a34f78d2ae6a18[3]);
            Iede5d56e52612e083407888da49470e5 = I29b4fdd4c13c96461c76660df767ea73(I2fcbccd884710be9c6a34f78d2ae6a18[4]);
            I3b2739319710681986b9d3f8cd04f619 = I29b4fdd4c13c96461c76660df767ea73(I2fcbccd884710be9c6a34f78d2ae6a18[5]);
            I850c257a0412bd9bd6001817bd9d0ee1 = I29b4fdd4c13c96461c76660df767ea73(I2fcbccd884710be9c6a34f78d2ae6a18[6]);
            Ib7875bf9d30d071e62a474c50d88ba06 = I29b4fdd4c13c96461c76660df767ea73(I2fcbccd884710be9c6a34f78d2ae6a18[7]);
            Ia92b76ee5b7d82a992a1b58147c0c0be = I29b4fdd4c13c96461c76660df767ea73(I2fcbccd884710be9c6a34f78d2ae6a18[8]);
            I2253b32e46200a23dba243819fce02f0 = I29b4fdd4c13c96461c76660df767ea73(I2fcbccd884710be9c6a34f78d2ae6a18[9]);
            I1b01cadaac7d3d15007f0afe5c0ab0f2 = I29b4fdd4c13c96461c76660df767ea73(I2fcbccd884710be9c6a34f78d2ae6a18[10]);
            Ie96877deef8b1676138f814c4a720800 = I29b4fdd4c13c96461c76660df767ea73(I2fcbccd884710be9c6a34f78d2ae6a18[11]);
            I8ce945d9f70bb317064a8d2d4eafd2d3 = I29b4fdd4c13c96461c76660df767ea73(I3d3df5d4d89adf508497bac8d75ef0c6[0]);
            Iaed105b99eae5b078521e3a94d8a79b7 = I29b4fdd4c13c96461c76660df767ea73(I3d3df5d4d89adf508497bac8d75ef0c6[1]);
            I05a812cd935867d1e417c64c26ea0952 = I29b4fdd4c13c96461c76660df767ea73(I3d3df5d4d89adf508497bac8d75ef0c6[2]);
            Ic0a580f94f3d03f72e3a487f84bf6612 = I29b4fdd4c13c96461c76660df767ea73(I3d3df5d4d89adf508497bac8d75ef0c6[3]);
            I39d9044227c161f0163e58dd82aadc90 = I29b4fdd4c13c96461c76660df767ea73(I3d3df5d4d89adf508497bac8d75ef0c6[4]);
            I5f607bdc9b276fdf07a17a11a20a6720 = I29b4fdd4c13c96461c76660df767ea73(I3d3df5d4d89adf508497bac8d75ef0c6[5]);
            I12e8b8cf609c2fbdc72efce9bb5dabee = I29b4fdd4c13c96461c76660df767ea73(I3d3df5d4d89adf508497bac8d75ef0c6[6]);
            I6fdccefd034e8b4b86cfa997502512ae = I29b4fdd4c13c96461c76660df767ea73(I3d3df5d4d89adf508497bac8d75ef0c6[7]);
            Idcd5283cf7b42d403ee0e4404b5b311b = I29b4fdd4c13c96461c76660df767ea73(I3d3df5d4d89adf508497bac8d75ef0c6[8]);
            Ia020344403aad35e050765a4b0cc42b7 = I29b4fdd4c13c96461c76660df767ea73(I3d3df5d4d89adf508497bac8d75ef0c6[9]);
            Id11fd3a31b70da0e64138e71840cfb83 = I29b4fdd4c13c96461c76660df767ea73(I3d3df5d4d89adf508497bac8d75ef0c6[10]);
            Ie9c5e7c98281cd1deb6acc51590c9d9a = I29b4fdd4c13c96461c76660df767ea73(I3d3df5d4d89adf508497bac8d75ef0c6[11]);
            Ia0e77e9544481aa0f56dfdb6eb253137 = I29b4fdd4c13c96461c76660df767ea73(Iadecdac113e45cd08e095317d07766e5[0]);
            Iec0d7ea31e0f1a75b15121090dcf1e11 = I29b4fdd4c13c96461c76660df767ea73(I2e4a339cb29f80caa8cbd630a0372ae8[0]);
            Ia98bb3648ce3719b1c31ce0f41121c63 = I29b4fdd4c13c96461c76660df767ea73(I423e8e9a9f19cf712372622e5c80c732[0]);
            Id9c8055ef530f2cb8096cb7bb2af55a4 = I29b4fdd4c13c96461c76660df767ea73(I5434db7480d96327d98156af57961745[0]);
            Ib9081d438413a627f5b16f68c2eabb80 = I29b4fdd4c13c96461c76660df767ea73(I20ebcbecf2c13a53be05ff26552b4e72[0]);
            I9c5bf5451736358f8c84e150004fa5a9 = I29b4fdd4c13c96461c76660df767ea73(I7ba72e4bac9bd64d046733ce50f43769[0]);
            I377933518c3807edb71f648c65ad5c85 = I29b4fdd4c13c96461c76660df767ea73(I6614526a756edaabd6a25e858b472d14[0]);
            Icec98d794a64752081fadfa74308fad3 = I29b4fdd4c13c96461c76660df767ea73(I47b2e8ee0c69e5301365a25d512b1ece[0]);
            I7bbe4d0a7d61d3f7da346de71b9a3a5f = I29b4fdd4c13c96461c76660df767ea73(Ibb72eb38996b41ce253875df0f620eb7[0]);
            I197c05f74bf7fb8d44124d40bd7c6563 = I29b4fdd4c13c96461c76660df767ea73(I66944cd8c5bc22cd92a5cfcd68cee426[0]);
            I92acc55d81ec6e02880337b0a451ae21 = I29b4fdd4c13c96461c76660df767ea73(I8f2ff78b78e43fe7f6780f19d92ff7b8[0]);
            I35c0ca76b28cd2f9355276b5d2f29ad4 = I29b4fdd4c13c96461c76660df767ea73(Ieea0e49da41cdf0d062217a6e6591728[0]);
            I29da0e5661f29bd8493c19885c998582 = I29b4fdd4c13c96461c76660df767ea73(I699c35d4b3c36c35ecaadb87c8b35d9a[0]);
            I9426c8c1b4d988d5cd7d89a7aed4f8fc = I29b4fdd4c13c96461c76660df767ea73(Ie6c95c6ddde379ca7437e78c42a8245e[0]);
            Ibd010f15e36194cbd2ce9f01c98a2b6f = I29b4fdd4c13c96461c76660df767ea73(I85e05de515eb28d7172a95ba55da82a2[0]);
            I7e86ab53e6d9647b230a94e076831ba2 = I29b4fdd4c13c96461c76660df767ea73(I7ed14b994ecbeae0536a721e16c88489[0]);
            Ia0ecfaedbc1d546d484978fd50096d10 = I29b4fdd4c13c96461c76660df767ea73(Iad29b892bf50a3e83e4eb9b7c271292a[0]);
            I27098cbe2d4fdd634385d771cc290c2b = I29b4fdd4c13c96461c76660df767ea73(I35d2bc3f0efd23ded421f195b62a6a33[0]);
            I5d7a0739e447775e00115799c52b11dd = I29b4fdd4c13c96461c76660df767ea73(I4aaa94237ac5b28ce1d0db0d4e15ff81[0]);
            Ie95793e09085b6de1383a37cc7fc41ac = I29b4fdd4c13c96461c76660df767ea73(I137145b608dfe5138d4bdbea237743bd[0]);
            Ib24b68cb35da39a743e1d90bba3f0836 = I29b4fdd4c13c96461c76660df767ea73(I68a784efb51b172af79e3dec88d529e1[0]);
            Id4cdd72193e90dddd211af73d7f3634a = I29b4fdd4c13c96461c76660df767ea73(Ic3036adab4495c6a59055dd34a28b2e5[0]);
            Iccab4c19a9190689f90a42160e2379de = I29b4fdd4c13c96461c76660df767ea73(I84a699063d2a7944f4a1b72b67ab5b4f[0]);
            I275ea08a3dc0600d8ccb6300eb7f2a6b = I29b4fdd4c13c96461c76660df767ea73(I63acf3ed504ad084a12a219790842b4a[0]);
            I1b53098a7240d2b5dc1f5c5c3b4bcc11 = I29b4fdd4c13c96461c76660df767ea73(I23a2a7fb24650eec8812d8671d92bf2b[0]);
            I278659ca1a0b093fc883d01987989dc0 = I29b4fdd4c13c96461c76660df767ea73(I6f9156b7b5e13529ec0c34da34cb2b04[0]);
            If92e66cba66732798dd19f968a5ef8ce = I29b4fdd4c13c96461c76660df767ea73(I09a4c92baceef72d764c6880fb62c1f7[0]);
            I784c4e9fb75c314f271477e0621aaf7c = I29b4fdd4c13c96461c76660df767ea73(I13a44a5dfbb198be64c99845122a6e97[0]);
            I3d3aafdd4d9d3e9fdab1f487c48a0ea9 = I29b4fdd4c13c96461c76660df767ea73(I2b57472e34677b9aafb852a3e421270d[0]);
            Idb4c722992139f39914af7085378c6cc = I29b4fdd4c13c96461c76660df767ea73(Ic96e056f2208c211122e5008d5fd8ced[0]);
            I63c9deb7e6a4b400e0aff6887a09e647 = I29b4fdd4c13c96461c76660df767ea73(Ie6b1ee6dfca427a82e4d1016585682d9[0]);
            Ie6f67c6e4c5e2b8357c0a902979e8722 = I29b4fdd4c13c96461c76660df767ea73(Ieb0276790e2d912809acc7f3a409ac37[0]);
            I1d7a4f99e3975fd01bfe5a9a1da84765 = I29b4fdd4c13c96461c76660df767ea73(I9883bdcc250c2eb1f8e691d0f18b3cbc[0]);
            I059d847e09f5aa3f6a8147062f4b13bf = I29b4fdd4c13c96461c76660df767ea73(I28f58fec52ea2df3fa3d8e4a2722468b[0]);
            I48e5256ade4d061a3b5ba08a53252bc3 = I29b4fdd4c13c96461c76660df767ea73(Ibf1bb88a30c8519cf22f684a9bc552e9[0]);
            I635fb29c55e0fb5cff0b6f443c2e3de5 = I29b4fdd4c13c96461c76660df767ea73(I9d2131bc965972708385d8d79c5b1687[0]);
            I088c5b971a2def57248769a33b7d2a2d = I29b4fdd4c13c96461c76660df767ea73(I65dc268c49445ceeef922f9c273df755[0]);
            Ide22394fce1658f9e7002bdb30d03c2f = I29b4fdd4c13c96461c76660df767ea73(I7c0af5fba885dca550df150029e9ee36[0]);
            I9ff276a14d3205b98174a8a736f79774 = I29b4fdd4c13c96461c76660df767ea73(If26299fbf3d11a469aa2bc573760fed0[0]);
            I123255637493b9c7924e3a72d1b86ee9 = I29b4fdd4c13c96461c76660df767ea73(I2ba80daf0c2b625370644ab47cef63e9[0]);
            I87e6ef84894cfc86b94e19c9d3065bc6 = I29b4fdd4c13c96461c76660df767ea73(I0911e01c831a9e46568122fa6dab2357[0]);
            I4c32900878260a261bc5403e8abd6258 = I29b4fdd4c13c96461c76660df767ea73(Ic8f0aa27dadc689b1bfb5b284fc13562[0]);
            Ifc100357ae3f754fb0e3863334bcc764 = I29b4fdd4c13c96461c76660df767ea73(I5ad4c6aba210a8b2d343ab17b49c38a3[0]);
            Iefe9e5376010997c0ee52eeb28e57a25 = I29b4fdd4c13c96461c76660df767ea73(I34947a54412d287f3ff730332211dc5a[0]);
            Ie6060acdcb16b6fa6aeeb649ed621053 = I29b4fdd4c13c96461c76660df767ea73(Ia6ac380b9be591fb53c0f36f4d417a7e[0]);
            I46c2b923860b0d1c01b9475f4467f280 = I29b4fdd4c13c96461c76660df767ea73(Ia5d5342af30d46f66f0e4f41e5170b87[0]);
            I38b4eceb159ecb0dda3920290a21a02a = I29b4fdd4c13c96461c76660df767ea73(Ica011579f46e949eda7f8eed2e4d3ada[0]);
            Ic45561ffe1837c3d5bb42c695a377f82 = I29b4fdd4c13c96461c76660df767ea73(I88b214aeebaffa768ccf7c70423fb0c3[0]);
            I3e76abc721bf7ed186f4d0f8f4bbf4e3 = I29b4fdd4c13c96461c76660df767ea73(If46340645f788fdde3bb8f4d176aae52[0]);
            I1afb4061458e9d2f5799afa1f2373bd2 = I29b4fdd4c13c96461c76660df767ea73(Ib59f285283d8c3013c20aad73ed9d148[0]);
            I18bb9a781a4c314fe6bd990e4c275f67 = I29b4fdd4c13c96461c76660df767ea73(I3229ea9a0c348b17fcaedf6565d6d7cc[0]);
            I49d7342f105c4502377abd23db973752 = I29b4fdd4c13c96461c76660df767ea73(I3ba17818aa7ea9bbfcebb2a5f405fec1[0]);
            Ieeb12d463444ca36af1ecf2e09504c06 = I29b4fdd4c13c96461c76660df767ea73(I2ad1769ceb4cf0013f7b032c6e583745[0]);
            I17525df1798fa2c1c4bbc4a1ddcdd0a5 = I29b4fdd4c13c96461c76660df767ea73(Ib35d4bfa08a9364f7f6c8be7feaf15ba[0]);
            I90c44c31fa7903a81826c1c568597362 = I29b4fdd4c13c96461c76660df767ea73(I216edc2024d31f612d05617f6696c6c5[0]);
            I3997cf122743b612f49cd5dd125a9201 = I29b4fdd4c13c96461c76660df767ea73(I2be51c29373fe2ddfe456265a54bcc08[0]);
            I1112c4267582ddb8148ee40d9529beee = I29b4fdd4c13c96461c76660df767ea73(Ib3561cb8090e7787ad8c324db3a5456a[0]);
            I21c207af859b94634d3750482b42a2ca = I29b4fdd4c13c96461c76660df767ea73(I5d701e34c6fea83dccbac286a36fcbbc[0]);
            I2ff2421bd86bf9ec110724460f1171e9 = I29b4fdd4c13c96461c76660df767ea73(Ie479179aee4de4208dda8af63ed9fb66[0]);
            I6ba5c453b17e4b33c61caf5d70041c4a = I29b4fdd4c13c96461c76660df767ea73(I0acbd9a7ed1409c7958d6c630a7f96d7[0]);
            I08318099725fbe033ab8d5427eb8b278 = I29b4fdd4c13c96461c76660df767ea73(I390dbe9907497b62162445c90f2f27fc[0]);
            If36cb462cdf20b0b1758cd6417e524fa = I29b4fdd4c13c96461c76660df767ea73(I01d386885d97d770ff2ab01da72631a0[0]);
            I40e8463645b1122b7cb224770fa00447 = I29b4fdd4c13c96461c76660df767ea73(Iedbfdad739e796202d764f909e6ac6b2[0]);
            Ide386e751e06dd5df0c042cd76f0f800 = I29b4fdd4c13c96461c76660df767ea73(I41ded014d071bd714d053a8aed21cf5a[0]);
            If63bb4681bf1116c0d1db3aa21bf52ac = I29b4fdd4c13c96461c76660df767ea73(I1f14df209c8c73fe390873ae05063afe[0]);
            I566c72342c69969892480fae41232c37 = I29b4fdd4c13c96461c76660df767ea73(I510a362375a9b9c75436ad01388de6db[0]);
            Ia0f7deea6b1ce1050dcf97fa99de9178 = I29b4fdd4c13c96461c76660df767ea73(Ic2f0b44a83961b8b49f4637ec6750f27[0]);
            I992b9876530d53c1b62d98511bf41942 = I29b4fdd4c13c96461c76660df767ea73(Id5cbccb1a2ccacf28b64ece8eec0099e[0]);
            Ib8861f627f6273c0a031bf43e7812a5d = I29b4fdd4c13c96461c76660df767ea73(I9686b2d0e5248bfb6d3ef9b7c687ed05[0]);
            Ieb5bac4ef0f5e4e0b826cdc43ae71471 = I29b4fdd4c13c96461c76660df767ea73(Ibe5129eb30f626925a3ab5ed5e239bb3[0]);
            I3cd0883d9f0ba7475f474f1e318ef023 = I29b4fdd4c13c96461c76660df767ea73(I2a656dad40cec86a53e732e78f00c269[0]);
            I5f8a41ab83a9257e534973e981e28e9b = I29b4fdd4c13c96461c76660df767ea73(If06132c6a0060efdbd695b31c338faf6[0]);
            I0e420136675d5f0d1aa027d589ee8741 = I29b4fdd4c13c96461c76660df767ea73(I02fd20ab9e4fa12009b63fbe41d647fb[0]);
            I4aab6ff52e3fba90bb7417cb50766125 = I29b4fdd4c13c96461c76660df767ea73(Ibb97d541a2ed2b0cbad273a09fef5594[0]);
            I1ba7f209cb735471073e8051026a148c = I29b4fdd4c13c96461c76660df767ea73(I0905c7e3678f66095194058bb72d22fe[0]);
            I711c5cf9fd8c5161bac36060b3443503 = I29b4fdd4c13c96461c76660df767ea73(I81433ae67b7cb4dee0b2091f3819ea88[0]);
            Ie3591b22e0e127f04658da68d4846be9 = I29b4fdd4c13c96461c76660df767ea73(Ia6249382442d1dd3062acc63f891465b[0]);
            I409129c0bf5d361e9916b6dc98e69a7d = I29b4fdd4c13c96461c76660df767ea73(Ie4bd4c14051455f00efdb023c3b58173[0]);
            Ie4f4faa470f572da2081b63b6df6e392 = I29b4fdd4c13c96461c76660df767ea73(Ie64e67a2316af18c5835c3a32ae9290f[0]);
            I5011dfbbb0eccfebcff255e4a2c5e64c = I29b4fdd4c13c96461c76660df767ea73(Icaf94b3fea3e29ff77d4793b389c9d14[0]);
            Ie32ca6b91d1c55883be8f63acca78764 = I29b4fdd4c13c96461c76660df767ea73(I334991f6bfe06389e35b7a580982de1f[0]);
            I6c7965d39dc839a9df56e628c77a5457 = I29b4fdd4c13c96461c76660df767ea73(I6390495458553670944cdbf57bd6ce7b[0]);
            Ieac9cea5f36bd82f87105b530e8fb614 = I29b4fdd4c13c96461c76660df767ea73(Ibafc73f0a3486943914e197a7af4505c[0]);
            I79657595561eac53237215fb4110f09d = I29b4fdd4c13c96461c76660df767ea73(I2ec83b82756dda6035ddff10dd41fed5[0]);
            I9b46463a6c54c3668e76190d942b7b38 = I29b4fdd4c13c96461c76660df767ea73(I5f6abb1000e5416dd4d43fcd052321fb[0]);
            I3ff883ad434cd5153b67186b6b21418d = I29b4fdd4c13c96461c76660df767ea73(Icc865d7264dd89944317be21610dcf9d[0]);
            I92abaae6fb89206885616877cca1e25a = I29b4fdd4c13c96461c76660df767ea73(I6a301412ef9235f3a609baf10a4200dd[0]);
            I33668b0ef7defef974b7a4c0f87689c0 = I29b4fdd4c13c96461c76660df767ea73(I9840f42586460341bb39256726d39ca1[0]);
            I338daeacf82ad288b14c6b5bd4099870 = I29b4fdd4c13c96461c76660df767ea73(I0837554bfb175a9ac8a4cb17e091fa9e[0]);
            Ibe085a39ecb07a8dca62002afa38df93 = I29b4fdd4c13c96461c76660df767ea73(Iacd698956b9ea6f1649063ee612c7e76[0]);
            I1f88dddf05f255942e2749891a7733da = I29b4fdd4c13c96461c76660df767ea73(I68928b2759202e358f75b08e162e6a68[0]);
            If1d0be4e9b995ec98c346e8392b9518a = I29b4fdd4c13c96461c76660df767ea73(I609f881624ec9034823c9f54f4fb9b6d[0]);
            I56a4443759b3d786bc9a34a0dc32abf0 = I29b4fdd4c13c96461c76660df767ea73(I075a0a1afc1463e92edb5f7658395424[0]);
            Ic826d371f2cfc503f5d9e43dc17481e1 = I29b4fdd4c13c96461c76660df767ea73(Idf1030f0e2aa5e2605bcea5fbe0428f8[0]);
            I5502f383dff392ef1be4cbbf9dbc3c2f = I29b4fdd4c13c96461c76660df767ea73(I1b82e98260c3bdeb5183a3af470e2d4a[0]);
            I96e6f1dc0cd451da6ac9170d5f83976d = I29b4fdd4c13c96461c76660df767ea73(I75338af3ebc7b7061a499e98a5be1674[0]);
            I10cd840a369d3e25556a41beede2be27 = I29b4fdd4c13c96461c76660df767ea73(I9f863d33f3c727e13eb52e7563ef9d1e[0]);
            Id85c2285fcc45211f0fa6963b74a663a = I29b4fdd4c13c96461c76660df767ea73(I56b8e0a7e6d2229baa9908843c0208ce[0]);
            Ie0bdfac78159144aa65090028931a3bf = I29b4fdd4c13c96461c76660df767ea73(I3d04bcd17aa2b98b69dcd671b9666c50[0]);
            I28fa30cd1f3b476fa6a354863108cbcf = I29b4fdd4c13c96461c76660df767ea73(Id254880ed38db79c53facbdc0c4a6d1a[0]);
            I7a927f4f266cc5253ec30f5c127bb17a = I29b4fdd4c13c96461c76660df767ea73(I988a7c2c284c38fcd6682236dc2d6151[0]);
            I7571c7c306861230de71a75fca79c5dc = I29b4fdd4c13c96461c76660df767ea73(Ida4c48caeba43eccdddd1748824ec551[0]);
            Ic79811a48840357d0b6303e7b19413dc = I29b4fdd4c13c96461c76660df767ea73(If9936b476bb351a9ecbb97e2088cdd6f[0]);
            I0f29300446f020dd23cf847d3e3d3530 = I29b4fdd4c13c96461c76660df767ea73(I6cbccfdeeb675a8a99d4c394bc8e71cd[0]);
            I802bd5b13c183c37e842f7e9278f35a9 = I29b4fdd4c13c96461c76660df767ea73(I79a4a9dfcecca4073c101bdd9b738c7c[0]);
            I0297905b35f06697625420b7fc2434f7 = I29b4fdd4c13c96461c76660df767ea73(Ice57a50f53d13e7eaf25af23547b5fb0[0]);
            I8487a819dcb61016798cde56f9662fcf = I29b4fdd4c13c96461c76660df767ea73(I8ff8106a70daac7c8932e88aeb6d198b[0]);
            Ia2904a5d5db43a209bd4b358ace68c6a = I29b4fdd4c13c96461c76660df767ea73(I8f9d1ec03357f7f045196050511341a2[0]);
            Ia8b29ca047a643f47bd3a0ffb50bf8cb = I29b4fdd4c13c96461c76660df767ea73(Ic423bfa7639075130324da59f2cca2fc[0]);
            Ic45d0537b94bc30713c0a0ee07b1ec40 = I29b4fdd4c13c96461c76660df767ea73(I4eed402353a7fa22fcb11f2adbf6be03[0]);
            I337231f0dc7eb85f7d950262e0adb724 = I29b4fdd4c13c96461c76660df767ea73(Ieb579bed6711928456b296873c5da9cd[0]);
            I530cf1f747d1df44b913f49eee90c079 = I29b4fdd4c13c96461c76660df767ea73(Ifdf316d14ef99080247091609b2c2a8f[0]);
            Ief52461e4a5ddb128be5e439edf34862 = I29b4fdd4c13c96461c76660df767ea73(I2a1afeffe5592e35349bfd4384de834e[0]);
            I46d86bfa6de26f3cfef9d802549ef2ad = I29b4fdd4c13c96461c76660df767ea73(I93f88eac6c04d26228b5d7a3b1d00a42[0]);
            If6a3bd6f002d91e0773c4ab9caaaa01e = I29b4fdd4c13c96461c76660df767ea73(I8c32ed7572af2a6a41a415ff6c580f3d[0]);
            Ib33e1c6d57e5e6fc465dc9c9a7cf29fa = I29b4fdd4c13c96461c76660df767ea73(I9cc4cd2860ebe1e5d43eb6024ea32dcf[0]);
            Id92a319da408be46970faf524513fdd8 = I29b4fdd4c13c96461c76660df767ea73(I35b73e275ce37c06d10c227595c7c3f6[0]);
            Iae182ffae6cea89363f0ccc8b5679561 = I29b4fdd4c13c96461c76660df767ea73(Iac4ee00e62d47494b2bfe3aff55506ea[0]);
            Idfe6aecb694385ce8c3c1544a4992a20 = I29b4fdd4c13c96461c76660df767ea73(I6023ec90efcd1ac53ea71eeee1c996e2[0]);
            Idfbc5726963cfa31bb4324143ffd08c7 = I29b4fdd4c13c96461c76660df767ea73(I6f2b0c5e254aeb7e967f86e914876171[0]);
            I205d5fdeae55fae7be2f06f11c949244 = I29b4fdd4c13c96461c76660df767ea73(Ie9353d9dd97f3536dfa6bcc2c662bf40[0]);
            Ie667e1755ae1561a2eefae9b63845dec = I29b4fdd4c13c96461c76660df767ea73(I09fd28ae4656b1282feb899a40b9b233[0]);
            If7348fdbe0400aab92e8fd6a7cf6c267 = I29b4fdd4c13c96461c76660df767ea73(Iabbb1734d7e19cd9c7329b30cb26cd3b[0]);
            I143b91852fddcdcc30bf1041332c4ed7 = I29b4fdd4c13c96461c76660df767ea73(Iacc03e49c3cd6749e4c49e13c8c8593e[0]);
            Iee5e74945ba15220f0f707c9c1927ba1 = I29b4fdd4c13c96461c76660df767ea73(I7913101e04088970adf3f1e7429cd06a[0]);
            I4d1c47569b0bc8c651c897ac8e88bd1f = I29b4fdd4c13c96461c76660df767ea73(Ibddcea3450984eb0b3cc3ca6961fa646[0]);
            Ib9d6c5be487a434fbafcda25ca9351dc = I29b4fdd4c13c96461c76660df767ea73(I0a863fcba425a8683ebbb35195ea70a4[0]);
            Ib0d033ba28e8c606ed92207049c76884 = I29b4fdd4c13c96461c76660df767ea73(I8138f45ab1b8a10869a2a6078b6c214c[0]);
            I300d9f403e33d860ff5dde9f91bae11b = I29b4fdd4c13c96461c76660df767ea73(Ie4c27f8574c8bad0b923796d2544f858[0]);
            Iebfe0fa45e4b34e142e82ddaa15243cf = I29b4fdd4c13c96461c76660df767ea73(Ibea29d15c71d594e4e9cbe6a58ebc550[0]);
            Ieb778442bc855e93e11c9b13f1a7ae06 = I29b4fdd4c13c96461c76660df767ea73(I0b249349485591abcc09c4587efca78d[0]);
            I57a393cc9cc9e1abc7962aa2cc840a7c = I29b4fdd4c13c96461c76660df767ea73(I6bbe05bfdabac8f312c7800eca53be62[0]);
            I0ffb8b65525af38861280645ac310e3d = I29b4fdd4c13c96461c76660df767ea73(Ie28e38c9881297e7ffae5c3aed4dfdd3[0]);
            I30fb41a57460a0b1f21065b4b97ddd42 = I29b4fdd4c13c96461c76660df767ea73(I1358b8ab0933bd596c33b622d2f9523f[0]);
            Ie8298c5c8ff538a3e37af46798f6d753 = I29b4fdd4c13c96461c76660df767ea73(I46ce01ea907e88cafb7d96d22b5fffd6[0]);
            Ie7dc322fee8ca0b6b9659e5183e0d6d6 = I29b4fdd4c13c96461c76660df767ea73(I64c0e39b2f3c34d724ecf0f511a413c9[0]);
            I91bbec0523f77fc52a88ebcc49267e9c = I29b4fdd4c13c96461c76660df767ea73(I6ffbd03867a92aea248506af197c2e86[0]);
            I38ae79956762380fadc94f8126dc1c90 = I29b4fdd4c13c96461c76660df767ea73(Ie0a0c3e63be2145dc838faf227a84044[0]);
            Id55a1ab9d158ea509e5f57286a3d1b67 = I29b4fdd4c13c96461c76660df767ea73(I58265e8a07eede7063d5a80db2412214[0]);
            Ice615e7e18356ae4c3f615dd997be943 = I29b4fdd4c13c96461c76660df767ea73(I6734d5f87b795f4a05510778c22b555c[0]);
            I57b40c72004f2c3072cbdefbeef72b7c = I29b4fdd4c13c96461c76660df767ea73(I314ced88cfc50d8b2edf129a6a3bf1a6[0]);
            Ie38351e19bdc4f2ce9caf75fc3937dd4 = I29b4fdd4c13c96461c76660df767ea73(I8cc6f1dc58a26262f18f334b751385ea[0]);
            Ibba6269b560db9d4913e1e515ed8270d = I29b4fdd4c13c96461c76660df767ea73(I18d34c481f17aae6b16b6d0a5aa85357[0]);
            Ie392719059587a201c0148138ba2a2d4 = I29b4fdd4c13c96461c76660df767ea73(Ib54b35abe1088393d275f4f45f7ed966[0]);
            I4852d6bacfd82fef6fab4502d61e9a37 = I29b4fdd4c13c96461c76660df767ea73(Ie339493197828e5bd69bc49ca91aeb1d[0]);
            I9200526d94c38e638370e9a2d7fed75c = I29b4fdd4c13c96461c76660df767ea73(Ic5084e34e9626f2e423283a87ea0d91d[0]);
            I15b8aa7d973edcf3b2365040f5570d82 = I29b4fdd4c13c96461c76660df767ea73(I3fee16f7ef907bcf1e2f5b2e7ec77866[0]);
            Ic3f8e77259ee3eb5be80e11b607818bd = I29b4fdd4c13c96461c76660df767ea73(Iee529a0d30e79cdc9b33dd3d876a0f23[0]);
            Iabf228f57ac154c417389f6711af1950 = I29b4fdd4c13c96461c76660df767ea73(I6c7373fafcfbb14c527e38e0f4440404[0]);
            If37de611ce4fa330c4fc9dcb87d4d95c = I29b4fdd4c13c96461c76660df767ea73(Ided1b79349f8806da8f5c6898cea94bc[0]);
            If3c44eb85217da3b6bddb5aed97a9bb7 = I29b4fdd4c13c96461c76660df767ea73(Id77e3ee5aded95fe141c26ad08639538[0]);
            I8c36318c45dabe6bf540381373f09fe5 = I29b4fdd4c13c96461c76660df767ea73(I3c286283659a38021c27b5e5346b59b0[0]);
end


   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
            Ib0973b6e90e7678addcb064fded7ce0f <=  1'b0;
            I5033323484d90d6bfbe03749019fc6dd <= {MAX_SUM_WDTH_LONG{1'b0}};
            Iee06707670e19a82d911c1750bcfc811 <=  1'b0;
            If5dad13ac41b3034bdb034bc86c9b348 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Id8d5df9e869aaeb107a41a6bca3b89bd <=  1'b0;
            Iac428f9f798618e1ef495c626c41892b <= {MAX_SUM_WDTH_LONG{1'b0}};
            I507f8602a99a1096e4c293ba3c235bbb <=  1'b0;
            I5a6427c8f18b36d2ea18fe60a0831ef1 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ibdf2178bd18783c4797c21e642388d16 <=  1'b0;
            Icc29441eac6ca7a138d45743d37505e3 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I2c690809d9b9e3482fe5a133b5c00afa <=  1'b0;
            I0e7754dcbc04a4850e052ae4a2fbe328 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I369ffa98995ba0834f8029ecce705c56 <=  1'b0;
            Ia30c019ed8ce395556494a92e7b42a92 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I9ccef4c47ae7cfab43584de0f2e193d3 <=  1'b0;
            I9799695ea8244992a6694eaf5c8ae64d <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ief31fe169c1b360d5933558208dbb602 <=  1'b0;
            I4524cd664b4cb41f642c675fa484c84b <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ib8c0317dafcfb91b3da5eb5afae1f2e2 <=  1'b0;
            I64e959d80af111ed2fcd54a5407d21bf <= {MAX_SUM_WDTH_LONG{1'b0}};
            I54e3f08f6f4cf784da57ac39f246b8fd <=  1'b0;
            I3e0da4bcbab4804b5397fb3aa2c94f51 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I16c7f1b874b0d05c6d120bbede254416 <=  1'b0;
            I3740b30d31f3c61d93a14a46e3199c4d <= {MAX_SUM_WDTH_LONG{1'b0}};
            I0c3cb2de514ecab0dd311e86a4dc3cdb <=  1'b0;
            Ibf0a30abfec9031737eada436ac1a0d4 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Icc5ba4554d7a44bc3b43377efbe3b5f8 <=  1'b0;
            Id36e8953a02400a5ab1f4dfdb0422e6d <= {MAX_SUM_WDTH_LONG{1'b0}};
            I5e51f49adb6dce65a9f19ff736526c4b <=  1'b0;
            Ica71108a53bfcfd1892b4d03ef68110c <= {MAX_SUM_WDTH_LONG{1'b0}};
            Id57092394c7cda397f42374df4aa3fec <=  1'b0;
            I7c97629ec6e594f9b2160815ddd133cc <= {MAX_SUM_WDTH_LONG{1'b0}};
            Idd6a4f8ae94c431f2fa3312b4fd287ba <=  1'b0;
            I4823c8239ace86dc399e906c1b5a0d74 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I9f1f8590dcf596097bc81001d51684b9 <=  1'b0;
            I10ad572ca72c2ea991487c39f7eabd7b <= {MAX_SUM_WDTH_LONG{1'b0}};
            Icecd765baa87877675b0f3972d78c02f <=  1'b0;
            Ie9f3fd3a6d16316e55addbe0e336519f <= {MAX_SUM_WDTH_LONG{1'b0}};
            I401a38ea1d71dcc71d17a4694ceb0988 <=  1'b0;
            I07965bca84276dd56da1af98e64b0adc <= {MAX_SUM_WDTH_LONG{1'b0}};
            I3db9b61e28a51e974e2d5e323ad53c1e <=  1'b0;
            Ic2ade31b8bcf68c4dcc1a371ff14074b <= {MAX_SUM_WDTH_LONG{1'b0}};
            I96d0a4387f9b959bc779ac13351182cc <=  1'b0;
            Ic0edcf240048fbfde4e938c3e4c5e281 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I64082bc75fdbeb69a52a4361ed2d5883 <=  1'b0;
            I8b42e89ff5f780d4ef8cd1cd5c99ef61 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I62929057b7c214bd38fd532e20ba5623 <=  1'b0;
            I70b1b8521b36920707e95fc9418eb8a9 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I641179f37fef63e7deec603b3291381c <=  1'b0;
            I4fb1c32a62cbbaeb585c6564a3c938f9 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Iff04b7ec87148f5bd408b4ec4b0590a5 <=  1'b0;
            Iefc37daeec14e14ef2fe0716f73109dc <= {MAX_SUM_WDTH_LONG{1'b0}};
            I198bfb18d6f91c8f62777e6f592a88fa <=  1'b0;
            Ibd15f164f6d2ac9e5721a21464bc2c5c <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ia1562c88b4f56d8935c3a5d6ead0f816 <=  1'b0;
            I951dfff9507bb70214d48e03a0ebb3a7 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Iaccba3030d9d9f8a56f86d6e34ed6325 <=  1'b0;
            Ie78e30b2a2eda75d0df7d10fd67b5e36 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I953dfeeacee8c44c08d0a425fa549e49 <=  1'b0;
            Ia0b83a372dd4115dc4d61eb8ff0811b9 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I214a50bf9f879fe747904f4679fdd1f6 <=  1'b0;
            If5c5bcbbea01aa22f242b913f0d01929 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ic88f2c344a8ad254fc7d7034cb594f6d <=  1'b0;
            Iccba58cd3519fb4cc75a61b50da1d562 <= {MAX_SUM_WDTH_LONG{1'b0}};
            If299d1a4e044acbc70bc3b7bce9f86e9 <=  1'b0;
            Ibc0999e4d0b3cc2650f9348b8c204b14 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Idb373d2cf788f6a93a0e5df7f9179292 <=  1'b0;
            I2aeff1fb4b839a581acaf26f90f9113c <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ic73b8c8f76a985330d4ac1fa0cc28e7f <=  1'b0;
            I7d60d53f883f8187700c4e78b4c22f1c <= {MAX_SUM_WDTH_LONG{1'b0}};
            I134dfb2c57d8cdffd2789e2f442c3247 <=  1'b0;
            Id6fcf4b7af4a37c854a12e2ae80851fa <= {MAX_SUM_WDTH_LONG{1'b0}};
            I0c735e43be8030078ec10bdb6882e79c <=  1'b0;
            Ifa5e5f7d753964f14f0f16dbe552fd85 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ie9951415c1d599570af1787767caa2dc <=  1'b0;
            I900d471b087cf5a436c2ad66a84d8280 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I2630f187d63ba9b0af52c77093e6b760 <=  1'b0;
            I6d1434907f0292ea2ee47cbc5b52bfb9 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I83db667ace2f04ef4950e2c186e0e6a4 <=  1'b0;
            I938bef7ba7ae1739d8e6a6a7c117a1b1 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ie818c5ea3f3b879fded32e6cb06ca546 <=  1'b0;
            I6384a9416b2d1da01df1b2d7b16c5390 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I3a67a175863091a52844aae6ad277da0 <=  1'b0;
            I5097a79e7cf7a30d38ba198d1407119c <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ia3aba80aead67feab12e4800fef82322 <=  1'b0;
            Ib113c26c8dcf49c972c41a938059a787 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I1181d42b560fca7bb5c924a81a5db1fc <=  1'b0;
            I970c4a25a8bce82a9d2846679029fcab <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ie4e5f3d7c5d2df30653f5666d14567bf <=  1'b0;
            Ibe2af096ad2db26e54d8b4b3bb05175c <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ifd9345cf219c58291c0b437aac093d78 <=  1'b0;
            Ie48569c467fba0c1291f71d6080ebedc <= {MAX_SUM_WDTH_LONG{1'b0}};
            I4f2d7bb48918ce51efe6b3b12f9f8e65 <=  1'b0;
            I90e7ded06617b49cdb8b5301fe9c6a20 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ifa612e6208151c616c3a0319182a96f1 <=  1'b0;
            I4920014f5d017f4e840dc3b88526955f <= {MAX_SUM_WDTH_LONG{1'b0}};
            I9cb28a0cc6358610854c8f8d1dd3c707 <=  1'b0;
            I03b70553f1c501609400574ae7cd73f5 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I40bcc924f5cf1f7d587aa35267022261 <=  1'b0;
            I63c9bf68b43ed66c51b0f4c0ed92e9ab <= {MAX_SUM_WDTH_LONG{1'b0}};
            I5238f7273b05b8b9f376314acdc6cc42 <=  1'b0;
            If408dfead07757878cc878131bc7d6a3 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I7137f56eeb4c4ae08bbc238db4cd3441 <=  1'b0;
            Ia0857d63d309807789b6ff4f6028f1b3 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I02335be013799e2560a98b6a82a0c528 <=  1'b0;
            I53921b825c5e434b63bee0e1ecb7a517 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Id327bb65156c8307901dfcb4184bb65f <=  1'b0;
            I5e68f84e123c37f19a03c13892c77e19 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I56331cb7b310613016958553732cdf40 <=  1'b0;
            Id5270b57c6fb4b18db3bbd0a523e467e <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ie3b00960f8af88a5aba7a2104dfca9a7 <=  1'b0;
            I3c18a84617eb21472d53e598700d7f4c <= {MAX_SUM_WDTH_LONG{1'b0}};
            I7d1ef47f35b7a4c3ea2e4383732de398 <=  1'b0;
            Id36663e7a01fff3170833ecfecac1321 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ibb013f036fc42687a04bdcbe2d0bbd8a <=  1'b0;
            I8d3be15109c7007a79fecaac0d891626 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I77eae49d321f1d1e39dd7c75829aaedc <=  1'b0;
            I92169cc57291f20d336a479e392ec271 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I420a4d69a077dc1996ddb4b715d63e15 <=  1'b0;
            I6178b220b469b40dac39168057023a1c <= {MAX_SUM_WDTH_LONG{1'b0}};
            I652202a4dc8f102d29334b4811f5628d <=  1'b0;
            I55342938216a0ea0889f96c2f6c05ce5 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I0e33e0cdf39fc4cc99f6696e9f2784de <=  1'b0;
            Idf28431c76a84a48dd895979d2b11a63 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ib9479328689dec62f900946e56ba0eb4 <=  1'b0;
            I1ef61124c8d62e8f6a82a729fb091694 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I2728682c0f749d1a9e8afeacdf44bfb7 <=  1'b0;
            Ib8bb96f0372323e6a8072ca56fb9396d <= {MAX_SUM_WDTH_LONG{1'b0}};
            I07da3bb5f943db6271fe1867a358df35 <=  1'b0;
            I432f74dda4f6b1cebdf5ad59c659080b <= {MAX_SUM_WDTH_LONG{1'b0}};
            I61fc44808c85a75909b9d9fd4035f147 <=  1'b0;
            Idc689442305acd00f0f32416d8fb3773 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ic5075ee0ad355c20dd45ed594f2a8c3f <=  1'b0;
            Ida03738adc101c03c2229756bed2469d <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ic0a651f45a502ead495cf14f97d65bfc <=  1'b0;
            I4d14c75f28f3e516c259ea288996131b <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ic1c05ea22f708f620f626cc8c5ca309c <=  1'b0;
            I6e6cbbf430d57f347a0d70558af143d8 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I61a18378aadae4556da501ce997321b4 <=  1'b0;
            Ib7487df45118e44acec6b9d07bbd5969 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ib1fc521709a1ce2198fd8df5b41d0177 <=  1'b0;
            I492f382fea500462b3d0866240fb91b2 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I1bb5511c9cda1a595c45ecde48e9ebc7 <=  1'b0;
            I3fb3ebddaf28efb56092d19a1b4695de <= {MAX_SUM_WDTH_LONG{1'b0}};
            I4a29c37ed36b6e12f1f8e263c92bdbc1 <=  1'b0;
            I22a26b7f0b1c8c16b00597732ce2ab23 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I4bf02a07719402890405fb2e7b679ed9 <=  1'b0;
            I2ac08a2d8c917ecb37fbaf5325cb0473 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I75bd82990cb60b6d7ccd7aa2982da7aa <=  1'b0;
            I50ff8f51e75fb9ce3db983c2a0f57196 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ia6d3e38249f8a1208540b68f54c46769 <=  1'b0;
            I444bc340ffb7ef7b72d4d2e761d58872 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Idf548b72357ab28fd956791e84e5d65c <=  1'b0;
            I039c6cac5830759529595a958b7f65c9 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I50b6f2e0ef2831535ac8c18cd7ca9379 <=  1'b0;
            I0584de7d919236ab138e288a27d08ff1 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I4003a2515229ca8eb6fefa2bef289ca6 <=  1'b0;
            I086402c82ec67ae09a9e6360c58904b4 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I48672f8b83eef8c406694676746469e7 <=  1'b0;
            I1cefdc831c146187c77f861b3e2d1af0 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ia14a60c9497c0faf3f1f448ff2abe553 <=  1'b0;
            Ida9c16ae57d17b6faee8a54838860447 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I0ef3962dd323e8ec64c4a881bd4b3044 <=  1'b0;
            Ia3b9fb112f39dd0ccbf7555659369efb <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ie9b64c34e31dab63c03b3de4528d53fe <=  1'b0;
            Ib1bfcdc0c972aafc99116ed8c0511445 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I5941476ded9f6dc25d7394f5d133955b <=  1'b0;
            I7adff505c50450a04f1717cac1adebe7 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ib46c78ff661ee6fb69c704d39235ffe1 <=  1'b0;
            I699feb4382974a02b21cb387c13f7f3f <= {MAX_SUM_WDTH_LONG{1'b0}};
            Iadabc5abc7dfbc1dd747179ad7e37850 <=  1'b0;
            Idc99c3b23e49aca3c98f0685ea34441c <= {MAX_SUM_WDTH_LONG{1'b0}};
            I97a6b5f0976feceee3a5b5890d4d76a0 <=  1'b0;
            Ib67318fa6954ec8f3247927d34e74f8c <= {MAX_SUM_WDTH_LONG{1'b0}};
            I7217d4790fec9797a1eb8cab1ebce71b <=  1'b0;
            I8774ce3f11362915c4331d1026e452dd <= {MAX_SUM_WDTH_LONG{1'b0}};
            I3dd024db4130c105a6817e8a4935de0d <=  1'b0;
            I2392b2d17ffed6073875fbe8e92534cf <= {MAX_SUM_WDTH_LONG{1'b0}};
            Iae502e5a5ae518fb7b817afff28b7932 <=  1'b0;
            I3a4f0d3e32596ef05477f494768d4266 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ib8b2b1d90204af5b100379ecad20fc0f <=  1'b0;
            Icd08ff59cf6be3ba97698dd55703339e <= {MAX_SUM_WDTH_LONG{1'b0}};
            Idf0e651d0b13e167df3c0cc40d149c29 <=  1'b0;
            I985fb7ed22a8476ea322c9e3c2b3851c <= {MAX_SUM_WDTH_LONG{1'b0}};
            I89daaca029498d05ca62c095db439eb5 <=  1'b0;
            Ib985709316b1b0a9d3fa3c1eaf6c641f <= {MAX_SUM_WDTH_LONG{1'b0}};
            I0fe5a34ceda936d0924efdd07fad11e5 <=  1'b0;
            I4be898887dff6e2cebe53f135ece131b <= {MAX_SUM_WDTH_LONG{1'b0}};
            I7876cbb2b5d8aba3652ec8b218080dff <=  1'b0;
            I004db04f61fb57aba81e15cc015442b3 <= {MAX_SUM_WDTH_LONG{1'b0}};
            If692ff56ce90d22d7af881599c54df75 <=  1'b0;
            I8f7e3dfb2f728d4cd1e79b82b62b0406 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I18a7a4fe8931c79df3a69223af46c440 <=  1'b0;
            I991054370345e61638ddaf81785505bd <= {MAX_SUM_WDTH_LONG{1'b0}};
            I8eec3538b8cc9c046954b6804cc656b0 <=  1'b0;
            Ifa1f503965270d10e7a5c9a15576069b <= {MAX_SUM_WDTH_LONG{1'b0}};
            I653767e659590c1676edf6c25fc0e253 <=  1'b0;
            I24f773842a4742fb58d09cae45717b2f <= {MAX_SUM_WDTH_LONG{1'b0}};
            I5ff863be142b92dff89f7916d0d088c1 <=  1'b0;
            I5bac7e0d778a547a0ae764fe259b6f7a <= {MAX_SUM_WDTH_LONG{1'b0}};
            I49f9fd0e0719be527f2a54814dab83ea <=  1'b0;
            I255577ebee6768871df0224fc1db2db3 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I945f2476eb599844cbee0cd89038e392 <=  1'b0;
            Ia7fb4af3d3529a32f902a52cf5598474 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ied0c5f8a9243cd9d93672ad6cc907d21 <=  1'b0;
            I2c98806141f064c9e92935b23a84ede1 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I9134c7f579723c7615af60b4344efe76 <=  1'b0;
            I5680847bc8d224fa4ed93b2fc0d841e1 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ie92388a9d1e71d73c07ed86e9bf6c887 <=  1'b0;
            I365254279ebb10dd7ba0b3482d5e34cd <= {MAX_SUM_WDTH_LONG{1'b0}};
            I6804fecdf59233c6cf14409bf2f1e430 <=  1'b0;
            I57bf4ad773cc058ae1bb7b1911dc3174 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I9e777a342bf53eaba0280737ae404bc1 <=  1'b0;
            I57072dfb29c4a3d2e2b40e46e62f0d95 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ied53820aab06b5c3423b1d878c71948f <=  1'b0;
            Id8cafb6f76321bdaba9711133be7be99 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I24cceded372d782c67b33f3a78b16045 <=  1'b0;
            I6344e71ca2b0fd39d36caedd889c3085 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I2e78d36bca5bfb016af674c343f9c041 <=  1'b0;
            I0c99a68e0bed90afce18807acf7d55bb <= {MAX_SUM_WDTH_LONG{1'b0}};
            I17a9a995de58643dbbfb78604f26198b <=  1'b0;
            I1c95650979c86310ae2a949961c9db11 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Iad642c4c62766e8f8bd5a1e9e73bdc80 <=  1'b0;
            I04eaefa5d133e53494fc270b07be7043 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I96f92481be1ac6cf985b8ab387d326bf <=  1'b0;
            I4a64fa2412eb8058c2dfd9351d7b297d <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ie03c09039ccafb427153d2347c1caea8 <=  1'b0;
            Ie8bb2fcb752c6a33254963d1ebb4130d <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ie7381a8294b4cdf669b9c57cfe4012b5 <=  1'b0;
            Iac05b7e3ae18f948b72c356ccfb8000f <= {MAX_SUM_WDTH_LONG{1'b0}};
            I61c9e3f8e42f869f4c9c1386325100b3 <=  1'b0;
            I27da3f75cca6c49e55db90306aa68e94 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I24c5b2de59eb1f43fe1efe687231c4b7 <=  1'b0;
            Idc7fed723190098341225fe01ba65ced <= {MAX_SUM_WDTH_LONG{1'b0}};
            I43d43acde5f831fc32b7bf5f10b9b3a9 <=  1'b0;
            Ife9065805598960919ee4f14c3cc6fd4 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ib06e93161fc8ca3be232f4261b04feb1 <=  1'b0;
            I717c5c2d6a2be61593492ae5f17a112f <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ia0dd00f83afc805036f2c6a0e38f725e <=  1'b0;
            I4c31fa8e6eb648439cdae1de1afe0d6f <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ib0a0f924fe3757a1e0aade7017ad9277 <=  1'b0;
            Iead549a9af27f1fced7d9c36e7b5c3f5 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I1ca949071d734d230cdb8adda46c9d79 <=  1'b0;
            I10422eb79364e7d0e21e1643d9060331 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I40170922c652fa7fa42abc6f580b5e3d <=  1'b0;
            I914cb87eba8baa40cd515334e59f26b2 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ib1ad0b531ac9028971d68f533e7ae566 <=  1'b0;
            I32ed679af4ab759901aee43c9d93eb67 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I0ab0170c7ceffbb58377b65d2ad92093 <=  1'b0;
            Id376dfa5141402f4d41a8858180ed87e <= {MAX_SUM_WDTH_LONG{1'b0}};
            I9ac68f228a93bbf4aa4a559b1364e42e <=  1'b0;
            I98a384bc62ee03f5ad7df20ef2d9af95 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I375c5f7eac92d853e85e0606011f3fb0 <=  1'b0;
            Icfed259ca2bb2732d8e0c26ef67cd4cf <= {MAX_SUM_WDTH_LONG{1'b0}};
            I94f9b1f2e63748c21ec7222c9641366a <=  1'b0;
            I20861535c450d6e6bf11c45dac120454 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I55500c1d85c4970932be67cc5cd2e023 <=  1'b0;
            I013929385ad819ddfcfcc59c22902ee3 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I36b487cd1a57a3a503e587fdefbb19e4 <=  1'b0;
            I34fffcb07fe82f11fe142f7c37f39155 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Icb5350e8c55a2adb370078a7575e28f8 <=  1'b0;
            I61ca60fde05ed88cce714dcd8c13b827 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I8a7a31327c9e4cbd88ce39fea8971caf <=  1'b0;
            I4907dd45c158dc7e0041c64f1fb388f6 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ied069655ed3775819d0bcb722d6d0488 <=  1'b0;
            I2c8f6a9b9f655b317bb0af4d60fdbc4b <= {MAX_SUM_WDTH_LONG{1'b0}};
            I78a5fc80d42e8db1b56cce5f4c97e325 <=  1'b0;
            Ic7dff631559304ec59f0696c66436d62 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I3ade7e345432319c1a9c91d4068b3ec9 <=  1'b0;
            I6a239d3e55b4a9a3be9989a85bbec545 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I88aed46f6dad7a81006562a720670654 <=  1'b0;
            I630f905e55f08e7d1569a08e937ad216 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I79e574dc9c7e18b695c9a2619b71b995 <=  1'b0;
            I8d13eb3669785c4279c685763d4f3fad <= {MAX_SUM_WDTH_LONG{1'b0}};
            I800ef583bec1d46d3d4ffdea6b312ef9 <=  1'b0;
            I25a6f3de9a9a01cbbdd32ed848561aa4 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I56cc5cd6d0a5a4e4601fd48e838fdaf3 <=  1'b0;
            Iba3dd4b2c2c85c4cfe770d9b52ef4634 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I21047a3955b8b89bdb9013d571b2bd0d <=  1'b0;
            Ie1b744387b5200a504e4874e14d2f282 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I56eb529a34b484cd20e29958cd6878eb <=  1'b0;
            Icf76cb69aedf4db01cd3444f4c4ba471 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I74588df6399af2c1112e3fa557e89e17 <=  1'b0;
            I4857b5b50556c8e7fff4b2d3e08e4b28 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ic8eae1a92f46db040eb22d726c3a0e6d <=  1'b0;
            I0a1e9cf99f1d4725327615f50fcc3ad0 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I854a15bc7e9728b01c9a1960f6248dc9 <=  1'b0;
            Ie844f4c446983ce381b0bc4c0e8ef7d7 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Iae332cfd000fd0529684ab787041b5dc <=  1'b0;
            I6067f47cccceea96ac46ff0d457b25f2 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I70148fe95244eebf7f0ec953703398de <=  1'b0;
            Ifd6fd1f3cbf8884ca7f64bc42278e4fa <= {MAX_SUM_WDTH_LONG{1'b0}};
            I24ee2d953e65fefdc73b3d3c4c0ddd05 <=  1'b0;
            Iaec9fd9e79371676bfa8ff14b4feae52 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ie3a5f8eec283fd4f682b5d0f909b051c <=  1'b0;
            I500757c4eda5d3d899aee47b87da585b <= {MAX_SUM_WDTH_LONG{1'b0}};
            I781d986d7fd6c2fec3a8cf3f29545174 <=  1'b0;
            I47bf091b0fa74ad511a760bad9d2506c <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ib4db8131350f8605e00907234aff901d <=  1'b0;
            Ia4c3d0cd9957f678880de5775de76e0d <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ie093f0750b60d3aed75705637933f34c <=  1'b0;
            If5f957fa2f055b1c2c28e8d7cfe3e9ad <= {MAX_SUM_WDTH_LONG{1'b0}};
            Id2fba7c1b3dc7a75a5e0d90494d56962 <=  1'b0;
            I3608378a5da8c66bef58528d56192530 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I9ecee74c445711a376133636ef414666 <=  1'b0;
            Ie6dead855e00ea0a8e6a9b7503aaebb8 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ifb3cf6b88835d27220df837682c4dc93 <=  1'b0;
            I3bae5e6862e003a8b9a476f72cc6858b <= {MAX_SUM_WDTH_LONG{1'b0}};
            I386fbb3bd550891d682e137044e8773a <=  1'b0;
            I4431adecba8be9e5f21bc6b3e1f8cb10 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I7ede7d2e1c2730b3b71340b11e880f5b <=  1'b0;
            I21c7a2885126d532d00484376588a469 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I64c65fad4a7d958d625c783626808175 <=  1'b0;
            I2c4d7339ff2fe68d060dd8d961dcab8c <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ib2e0cd0a2b51c3a265bdd20834c0ed2d <=  1'b0;
            Iee518b15b067eec58cccfa37f7432ea5 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I67be0b66c8d0680eb23290a4b3885af3 <=  1'b0;
            I42145be9c2a80288ba4a2edd91f661a3 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I01148401f7d058614dc1ae6ed3c8bd94 <=  1'b0;
            I9dc297ad41fafcda77f5347f331cfc25 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I3394319c370daf6102be00d938d55769 <=  1'b0;
            I846700c79f30ca954cc2933fc94d355b <= {MAX_SUM_WDTH_LONG{1'b0}};
            I24d6a334dd15ccdea558f32cd029e6d1 <=  1'b0;
            I8af96a91457316e49e3f7dd5e57c82da <= {MAX_SUM_WDTH_LONG{1'b0}};
            I3a41f68bca2d7edd1f5738c4fda8e73c <=  1'b0;
            I7d1c247500d7d32e406b2a5f7e2b745b <= {MAX_SUM_WDTH_LONG{1'b0}};
            I9ef1784d165492f3482d14f475732451 <=  1'b0;
            I66d85c030a8864505298919046056305 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I9d9378337a77515a4e8d04fb88938808 <=  1'b0;
            I4841257ae596d9d3e4eb1e6f886956b0 <= {MAX_SUM_WDTH_LONG{1'b0}};
            If0e20ef9aa69b77ae0e58ca3dfc9998f <=  1'b0;
            Icd6f7ec117f9ab4eda8c5eba41386ffa <= {MAX_SUM_WDTH_LONG{1'b0}};
            Iec2cb48bb1b58f268bf164d5e8a8120f <=  1'b0;
            Ibc0498839d1d9b6dc853b8e5d7a88fa3 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ia4ae7c98720d43a604f28dfc5dd67d50 <=  1'b0;
            I142ebca7f155e287e38ddf45423ab0fd <= {MAX_SUM_WDTH_LONG{1'b0}};
       end else begin
          Ib0973b6e90e7678addcb064fded7ce0f <=
            Ibc0871b3c992fd278815fdbefcd2bac0[0] ^
            Ibeb5edab51cd6aedad9c2ecedaded6f5[0] ^
            Ib0bf69cc797f330fb2546eb46d2d6f76[0] ^
            I5686b595177e07dd5bf231a35ee41659[0] ^
            I33a6ffad80ddf99a4d316a049078244d[0] ^
            I72a2f42b727a0503d43332c0f22d5ae3[0] ^
            Ic2580cbeec8c11a19bd1e2ebc29d255e[0] ^
            I6f5c991e5fdcf56d582c6f80eb6731df[0] ^
            exp_syn[0];
          Iee06707670e19a82d911c1750bcfc811 <=
            I8695e1e94cbfcbe4b9eae315b042529e[0] ^
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[0] ^
            Iec7404bc79c58d4d2538fcdf659e9134[0] ^
            I9c0b88a0be66d62f8ab061aeaee7e60f[0] ^
            I980165c1147ac5ff86619c841c6031dc[0] ^
            I8b8b9c4777e6df3eb2b9313e69ef2c8c[0] ^
            If79ed5ee2b8710da0608c1e245d07d55[0] ^
            Ia5cc3055ba3365e64cf59c4d4fd3f093[0] ^
            exp_syn[1];
          Id8d5df9e869aaeb107a41a6bca3b89bd <=
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[0] ^
            I5b7caaeb34c43e66e8d095a859e708fe[0] ^
            Ie1cd04c7668d3f450c387a6c1ad778c7[0] ^
            Id88b9265ff08e0730e6a41abe1f80a32[0] ^
            I19df055705f322292a3601fa63f0e5f9[0] ^
            I4a16e8e7946d9a8220304fc1be3fb362[0] ^
            I9497bbb4f746969a95cff948a3ee9ade[0] ^
            Iea7da1f43ba202d753b0edb0be8b3fcf[0] ^
            exp_syn[2];
          I507f8602a99a1096e4c293ba3c235bbb <=
            Ib58043c04b5c4c86c1c67e57cc66dcf7[0] ^
            I61f0c04673dfb262ef6912eb2df39120[0] ^
            If511a6ea6aa5cda5353658d8e192791f[0] ^
            I6330943c9295298c53e889d47c7904d9[0] ^
            I3d50cfeaa4b69c09bb648b8873a6bc24[0] ^
            I07930a807994815de45864af579902c4[0] ^
            I651d700a00d7004d8728bc7356f30926[0] ^
            I872f61d20baf011e867b44dc5539fc37[0] ^
            exp_syn[3];
          Ibdf2178bd18783c4797c21e642388d16 <=
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[1] ^
            I5686b595177e07dd5bf231a35ee41659[1] ^
            Ic2941d16ae6a5cbce70e8546a18ca4ff[0] ^
            I480a0f6d6c3eb936de10a72749f6cd3f[0] ^
            I980165c1147ac5ff86619c841c6031dc[1] ^
            I0e0b15868b02ca52b260f17f150d237e[0] ^
            I6ebab438dc55ccf6c1600313891d9c38[0] ^
            I07930a807994815de45864af579902c4[1] ^
            I6f5c991e5fdcf56d582c6f80eb6731df[1] ^
            Ieb244944e7ee8236a207924f56fbc689[0] ^
            exp_syn[4];
          I2c690809d9b9e3482fe5a133b5c00afa <=
            Ib58043c04b5c4c86c1c67e57cc66dcf7[1] ^
            I9c0b88a0be66d62f8ab061aeaee7e60f[1] ^
            I8e29ebe9ee25ea8ef3e52ff56fc29157[0] ^
            I50976b0051e84b6a42fc1dbabd7d20ae[0] ^
            I19df055705f322292a3601fa63f0e5f9[1] ^
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[0] ^
            I2fbf89398a148c47810456812dbee5a6[0] ^
            I72a2f42b727a0503d43332c0f22d5ae3[1] ^
            Ia5cc3055ba3365e64cf59c4d4fd3f093[1] ^
            Ie9b2be4c32334220e134e041ca8dfc06[0] ^
            exp_syn[5];
          I369ffa98995ba0834f8029ecce705c56 <=
            Ibc0871b3c992fd278815fdbefcd2bac0[1] ^
            Id88b9265ff08e0730e6a41abe1f80a32[1] ^
            Ic3742290179b27b9865f9d1f88d66266[0] ^
            I82e0e091fba6f79cef97eacac4b43ecb[0] ^
            I3d50cfeaa4b69c09bb648b8873a6bc24[1] ^
            I8e591d83170c8ba46d31c61935311b22[0] ^
            Icac5a9001ee113e612e3457b4b49ee68[0] ^
            I8b8b9c4777e6df3eb2b9313e69ef2c8c[1] ^
            Iea7da1f43ba202d753b0edb0be8b3fcf[1] ^
            Id6f07dee3e47f39e3b43329c26f690f7[0] ^
            exp_syn[6];
          I9ccef4c47ae7cfab43584de0f2e193d3 <=
            I8695e1e94cbfcbe4b9eae315b042529e[1] ^
            I6330943c9295298c53e889d47c7904d9[1] ^
            I9ef21ef20099af28d9a8c794f70d45a5[0] ^
            I04302edb2671c5bc0ca2673cd53935e1[0] ^
            I33a6ffad80ddf99a4d316a049078244d[1] ^
            I02b62fafd371de339f299f8aefec6c43[0] ^
            I9461e92a5880cb9e04fcece2ef4674f0[0] ^
            I4a16e8e7946d9a8220304fc1be3fb362[1] ^
            I872f61d20baf011e867b44dc5539fc37[1] ^
            Ic7f04c065f8ff82c2288f1de77d37189[0] ^
            exp_syn[7];
          Ief31fe169c1b360d5933558208dbb602 <=
            Ibc0871b3c992fd278815fdbefcd2bac0[2] ^
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[1] ^
            Id88b9265ff08e0730e6a41abe1f80a32[2] ^
            I9ef21ef20099af28d9a8c794f70d45a5[1] ^
            I6ebab438dc55ccf6c1600313891d9c38[1] ^
            Ic2580cbeec8c11a19bd1e2ebc29d255e[1] ^
            Ieb244944e7ee8236a207924f56fbc689[1] ^
            I4267622319ca65909a3b40484dc74d3a[0] ^
            exp_syn[8];
          Ib8c0317dafcfb91b3da5eb5afae1f2e2 <=
            I8695e1e94cbfcbe4b9eae315b042529e[2] ^
            I5b7caaeb34c43e66e8d095a859e708fe[1] ^
            I6330943c9295298c53e889d47c7904d9[2] ^
            Ic2941d16ae6a5cbce70e8546a18ca4ff[1] ^
            I2fbf89398a148c47810456812dbee5a6[1] ^
            If79ed5ee2b8710da0608c1e245d07d55[1] ^
            Ie9b2be4c32334220e134e041ca8dfc06[1] ^
            Iedd7d4ea8d082b40244c04946dfb14a0[0] ^
            exp_syn[9];
          I54e3f08f6f4cf784da57ac39f246b8fd <=
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[2] ^
            I61f0c04673dfb262ef6912eb2df39120[1] ^
            I5686b595177e07dd5bf231a35ee41659[2] ^
            I8e29ebe9ee25ea8ef3e52ff56fc29157[1] ^
            Icac5a9001ee113e612e3457b4b49ee68[1] ^
            I9497bbb4f746969a95cff948a3ee9ade[1] ^
            Id6f07dee3e47f39e3b43329c26f690f7[1] ^
            I56e1fe0c7a62589c123876f2b4e57a26[0] ^
            exp_syn[10];
          I16c7f1b874b0d05c6d120bbede254416 <=
            Ib58043c04b5c4c86c1c67e57cc66dcf7[2] ^
            Ibeb5edab51cd6aedad9c2ecedaded6f5[1] ^
            I9c0b88a0be66d62f8ab061aeaee7e60f[2] ^
            Ic3742290179b27b9865f9d1f88d66266[1] ^
            I9461e92a5880cb9e04fcece2ef4674f0[1] ^
            I651d700a00d7004d8728bc7356f30926[1] ^
            Ic7f04c065f8ff82c2288f1de77d37189[1] ^
            Ia8a468877c9f96713c8141df9205f92a[0] ^
            exp_syn[11];
          I0c3cb2de514ecab0dd311e86a4dc3cdb <=
            I61f0c04673dfb262ef6912eb2df39120[2] ^
            Ie1cd04c7668d3f450c387a6c1ad778c7[1] ^
            I8e29ebe9ee25ea8ef3e52ff56fc29157[2] ^
            I04302edb2671c5bc0ca2673cd53935e1[1] ^
            I33a6ffad80ddf99a4d316a049078244d[2] ^
            I8e591d83170c8ba46d31c61935311b22[1] ^
            Icac5a9001ee113e612e3457b4b49ee68[2] ^
            I07930a807994815de45864af579902c4[2] ^
            Ic2580cbeec8c11a19bd1e2ebc29d255e[2] ^
            I4267622319ca65909a3b40484dc74d3a[1] ^
            exp_syn[12];
          Icc5ba4554d7a44bc3b43377efbe3b5f8 <=
            Ibeb5edab51cd6aedad9c2ecedaded6f5[2] ^
            If511a6ea6aa5cda5353658d8e192791f[1] ^
            Ic3742290179b27b9865f9d1f88d66266[2] ^
            I480a0f6d6c3eb936de10a72749f6cd3f[1] ^
            I980165c1147ac5ff86619c841c6031dc[2] ^
            I02b62fafd371de339f299f8aefec6c43[1] ^
            I9461e92a5880cb9e04fcece2ef4674f0[2] ^
            I72a2f42b727a0503d43332c0f22d5ae3[2] ^
            If79ed5ee2b8710da0608c1e245d07d55[2] ^
            Iedd7d4ea8d082b40244c04946dfb14a0[1] ^
            exp_syn[13];
          I5e51f49adb6dce65a9f19ff736526c4b <=
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[2] ^
            Ib0bf69cc797f330fb2546eb46d2d6f76[1] ^
            I9ef21ef20099af28d9a8c794f70d45a5[2] ^
            I50976b0051e84b6a42fc1dbabd7d20ae[1] ^
            I19df055705f322292a3601fa63f0e5f9[2] ^
            I0e0b15868b02ca52b260f17f150d237e[1] ^
            I6ebab438dc55ccf6c1600313891d9c38[2] ^
            I8b8b9c4777e6df3eb2b9313e69ef2c8c[2] ^
            I9497bbb4f746969a95cff948a3ee9ade[2] ^
            I56e1fe0c7a62589c123876f2b4e57a26[1] ^
            exp_syn[14];
          Id57092394c7cda397f42374df4aa3fec <=
            I5b7caaeb34c43e66e8d095a859e708fe[2] ^
            Iec7404bc79c58d4d2538fcdf659e9134[1] ^
            Ic2941d16ae6a5cbce70e8546a18ca4ff[2] ^
            I82e0e091fba6f79cef97eacac4b43ecb[1] ^
            I3d50cfeaa4b69c09bb648b8873a6bc24[2] ^
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[1] ^
            I2fbf89398a148c47810456812dbee5a6[2] ^
            I4a16e8e7946d9a8220304fc1be3fb362[2] ^
            I651d700a00d7004d8728bc7356f30926[2] ^
            Ia8a468877c9f96713c8141df9205f92a[1] ^
            exp_syn[15];
          Idd6a4f8ae94c431f2fa3312b4fd287ba <=
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[3] ^
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[3] ^
            I872f61d20baf011e867b44dc5539fc37[2] ^
            Ida6059c6e0890f730536f97dfb83770b[0] ^
            exp_syn[16];
          I9f1f8590dcf596097bc81001d51684b9 <=
            Ib58043c04b5c4c86c1c67e57cc66dcf7[3] ^
            I5b7caaeb34c43e66e8d095a859e708fe[3] ^
            I6f5c991e5fdcf56d582c6f80eb6731df[2] ^
            I1993c1ed200d7cdf838d23c72a0c1c0b[0] ^
            exp_syn[17];
          Icecd765baa87877675b0f3972d78c02f <=
            Ibc0871b3c992fd278815fdbefcd2bac0[3] ^
            I61f0c04673dfb262ef6912eb2df39120[3] ^
            Ia5cc3055ba3365e64cf59c4d4fd3f093[2] ^
            I07e04e352df9aa1988ccf05d9cb2d1d7[0] ^
            exp_syn[18];
          I401a38ea1d71dcc71d17a4694ceb0988 <=
            I8695e1e94cbfcbe4b9eae315b042529e[3] ^
            Ibeb5edab51cd6aedad9c2ecedaded6f5[3] ^
            Iea7da1f43ba202d753b0edb0be8b3fcf[2] ^
            Ic4c0ebcc3711c9844a3aa3875483d2f7[0] ^
            exp_syn[19];
          I3db9b61e28a51e974e2d5e323ad53c1e <=
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[4] ^
            Ibeb5edab51cd6aedad9c2ecedaded6f5[4] ^
            I50976b0051e84b6a42fc1dbabd7d20ae[2] ^
            I02b62fafd371de339f299f8aefec6c43[2] ^
            I872f61d20baf011e867b44dc5539fc37[3] ^
            I28e344560ba76bb3b76d01d8c53693a9[0] ^
            exp_syn[20];
          I96d0a4387f9b959bc779ac13351182cc <=
            Ib58043c04b5c4c86c1c67e57cc66dcf7[4] ^
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[4] ^
            I82e0e091fba6f79cef97eacac4b43ecb[2] ^
            I0e0b15868b02ca52b260f17f150d237e[2] ^
            I6f5c991e5fdcf56d582c6f80eb6731df[3] ^
            I0600def6e6caada88ba6dedbb0d322ac[0] ^
            exp_syn[21];
          I64082bc75fdbeb69a52a4361ed2d5883 <=
            Ibc0871b3c992fd278815fdbefcd2bac0[4] ^
            I5b7caaeb34c43e66e8d095a859e708fe[4] ^
            I04302edb2671c5bc0ca2673cd53935e1[2] ^
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[2] ^
            Ia5cc3055ba3365e64cf59c4d4fd3f093[3] ^
            Iddbf50612c89b5b95a5c9efb5575cae3[0] ^
            exp_syn[22];
          I62929057b7c214bd38fd532e20ba5623 <=
            I8695e1e94cbfcbe4b9eae315b042529e[4] ^
            I61f0c04673dfb262ef6912eb2df39120[4] ^
            I480a0f6d6c3eb936de10a72749f6cd3f[2] ^
            I8e591d83170c8ba46d31c61935311b22[2] ^
            Iea7da1f43ba202d753b0edb0be8b3fcf[3] ^
            Iadc8f7f87b50bfff53d2d12d82489829[0] ^
            exp_syn[23];
          I641179f37fef63e7deec603b3291381c <=
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[5] ^
            I04302edb2671c5bc0ca2673cd53935e1[3] ^
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[3] ^
            I07930a807994815de45864af579902c4[3] ^
            Iea7da1f43ba202d753b0edb0be8b3fcf[4] ^
            I53a658b443200b9f11f1830547b5f42d[0] ^
            exp_syn[24];
          Iff04b7ec87148f5bd408b4ec4b0590a5 <=
            Ib58043c04b5c4c86c1c67e57cc66dcf7[5] ^
            I480a0f6d6c3eb936de10a72749f6cd3f[3] ^
            I8e591d83170c8ba46d31c61935311b22[3] ^
            I72a2f42b727a0503d43332c0f22d5ae3[3] ^
            I872f61d20baf011e867b44dc5539fc37[4] ^
            I170f424df45651abe215ec74d649a9eb[0] ^
            exp_syn[25];
          I198bfb18d6f91c8f62777e6f592a88fa <=
            Ibc0871b3c992fd278815fdbefcd2bac0[5] ^
            I50976b0051e84b6a42fc1dbabd7d20ae[3] ^
            I02b62fafd371de339f299f8aefec6c43[3] ^
            I8b8b9c4777e6df3eb2b9313e69ef2c8c[3] ^
            I6f5c991e5fdcf56d582c6f80eb6731df[4] ^
            I3c897bfed190017a876c44fd73a7ecea[0] ^
            exp_syn[26];
          Ia1562c88b4f56d8935c3a5d6ead0f816 <=
            I8695e1e94cbfcbe4b9eae315b042529e[5] ^
            I82e0e091fba6f79cef97eacac4b43ecb[3] ^
            I0e0b15868b02ca52b260f17f150d237e[3] ^
            I4a16e8e7946d9a8220304fc1be3fb362[3] ^
            Ia5cc3055ba3365e64cf59c4d4fd3f093[4] ^
            Iaecbbae967be2c62cacf2fa7f9801899[0] ^
            exp_syn[27];
          Iaccba3030d9d9f8a56f86d6e34ed6325 <=
            Ibeb5edab51cd6aedad9c2ecedaded6f5[5] ^
            I82e0e091fba6f79cef97eacac4b43ecb[4] ^
            I0e0b15868b02ca52b260f17f150d237e[4] ^
            I872f61d20baf011e867b44dc5539fc37[5] ^
            I4267622319ca65909a3b40484dc74d3a[2] ^
            I52f867f1009f2e8d18b50a777942bde3[0] ^
            exp_syn[28];
          I953dfeeacee8c44c08d0a425fa549e49 <=
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[5] ^
            I04302edb2671c5bc0ca2673cd53935e1[4] ^
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[4] ^
            I6f5c991e5fdcf56d582c6f80eb6731df[5] ^
            Iedd7d4ea8d082b40244c04946dfb14a0[2] ^
            I56a39a0c67b1de0a3cab6c61af3eebcf[0] ^
            exp_syn[29];
          I214a50bf9f879fe747904f4679fdd1f6 <=
            I5b7caaeb34c43e66e8d095a859e708fe[5] ^
            I480a0f6d6c3eb936de10a72749f6cd3f[4] ^
            I8e591d83170c8ba46d31c61935311b22[4] ^
            Ia5cc3055ba3365e64cf59c4d4fd3f093[5] ^
            I56e1fe0c7a62589c123876f2b4e57a26[2] ^
            I490a65b3f7b30540906262ec5e12717b[0] ^
            exp_syn[30];
          Ic88f2c344a8ad254fc7d7034cb594f6d <=
            I61f0c04673dfb262ef6912eb2df39120[5] ^
            I50976b0051e84b6a42fc1dbabd7d20ae[4] ^
            I02b62fafd371de339f299f8aefec6c43[4] ^
            Iea7da1f43ba202d753b0edb0be8b3fcf[5] ^
            Ia8a468877c9f96713c8141df9205f92a[2] ^
            Ib3c52fef8251d95e9abc8df0aad45d4e[0] ^
            exp_syn[31];
          If299d1a4e044acbc70bc3b7bce9f86e9 <=
            I8695e1e94cbfcbe4b9eae315b042529e[6] ^
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[6] ^
            Id6f07dee3e47f39e3b43329c26f690f7[2] ^
            If75725e534dcb00364d73a42769539fb[0] ^
            exp_syn[32];
          Idb373d2cf788f6a93a0e5df7f9179292 <=
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[6] ^
            I5b7caaeb34c43e66e8d095a859e708fe[6] ^
            Ic7f04c065f8ff82c2288f1de77d37189[2] ^
            I9ddc427eef437ecc3ac4a2cf52aad4c3[0] ^
            exp_syn[33];
          Ic73b8c8f76a985330d4ac1fa0cc28e7f <=
            Ib58043c04b5c4c86c1c67e57cc66dcf7[6] ^
            I61f0c04673dfb262ef6912eb2df39120[6] ^
            Ieb244944e7ee8236a207924f56fbc689[2] ^
            I8999ca1f2fe9d4a30bd38fcb0daad2a4[0] ^
            exp_syn[34];
          I134dfb2c57d8cdffd2789e2f442c3247 <=
            Ibc0871b3c992fd278815fdbefcd2bac0[6] ^
            Ibeb5edab51cd6aedad9c2ecedaded6f5[6] ^
            Ie9b2be4c32334220e134e041ca8dfc06[2] ^
            Ie11cf6677812bb739255b053a9c9cd56[0] ^
            exp_syn[35];
          I0c735e43be8030078ec10bdb6882e79c <=
            I5b7caaeb34c43e66e8d095a859e708fe[7] ^
            I2fbf89398a148c47810456812dbee5a6[3] ^
            If79ed5ee2b8710da0608c1e245d07d55[3] ^
            I872f61d20baf011e867b44dc5539fc37[6] ^
            Iacc1d5a5c7811f0c9326ef80d1154fbb[0] ^
            exp_syn[36];
          Ie9951415c1d599570af1787767caa2dc <=
            I61f0c04673dfb262ef6912eb2df39120[7] ^
            Icac5a9001ee113e612e3457b4b49ee68[3] ^
            I9497bbb4f746969a95cff948a3ee9ade[3] ^
            I6f5c991e5fdcf56d582c6f80eb6731df[6] ^
            I0efdadfd49c035a49d92243391395bca[0] ^
            exp_syn[37];
          I2630f187d63ba9b0af52c77093e6b760 <=
            Ibeb5edab51cd6aedad9c2ecedaded6f5[7] ^
            I9461e92a5880cb9e04fcece2ef4674f0[3] ^
            I651d700a00d7004d8728bc7356f30926[3] ^
            Ia5cc3055ba3365e64cf59c4d4fd3f093[6] ^
            Ie34d59bc77e06807937fe6f6860527e9[0] ^
            exp_syn[38];
          I83db667ace2f04ef4950e2c186e0e6a4 <=
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[7] ^
            I6ebab438dc55ccf6c1600313891d9c38[3] ^
            Ic2580cbeec8c11a19bd1e2ebc29d255e[3] ^
            Iea7da1f43ba202d753b0edb0be8b3fcf[6] ^
            I9661cb126908d8550b585e2bad383bd6[0] ^
            exp_syn[39];
          Ie818c5ea3f3b879fded32e6cb06ca546 <=
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[7] ^
            Ibeb5edab51cd6aedad9c2ecedaded6f5[8] ^
            I3d50cfeaa4b69c09bb648b8873a6bc24[3] ^
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[5] ^
            Ic0b832fbcbdb57745fefcc1ac1438808[0] ^
            exp_syn[40];
          I3a67a175863091a52844aae6ad277da0 <=
            Ib58043c04b5c4c86c1c67e57cc66dcf7[7] ^
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[8] ^
            I33a6ffad80ddf99a4d316a049078244d[3] ^
            I8e591d83170c8ba46d31c61935311b22[5] ^
            I2afd96714b26f30483c3935c2a68e64f[0] ^
            exp_syn[41];
          Ia3aba80aead67feab12e4800fef82322 <=
            Ibc0871b3c992fd278815fdbefcd2bac0[7] ^
            I5b7caaeb34c43e66e8d095a859e708fe[8] ^
            I980165c1147ac5ff86619c841c6031dc[3] ^
            I02b62fafd371de339f299f8aefec6c43[5] ^
            Id6d4165b752630a1ce7ceb77fdcee477[0] ^
            exp_syn[42];
          I1181d42b560fca7bb5c924a81a5db1fc <=
            I8695e1e94cbfcbe4b9eae315b042529e[7] ^
            I61f0c04673dfb262ef6912eb2df39120[8] ^
            I19df055705f322292a3601fa63f0e5f9[3] ^
            I0e0b15868b02ca52b260f17f150d237e[5] ^
            I59baaf1ad22721cde9064b8aad65ac76[0] ^
            exp_syn[43];
          Ie4e5f3d7c5d2df30653f5666d14567bf <=
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[8] ^
            I0e0b15868b02ca52b260f17f150d237e[6] ^
            I8b8b9c4777e6df3eb2b9313e69ef2c8c[4] ^
            I4267622319ca65909a3b40484dc74d3a[3] ^
            I9094f4e9c5b60add3acee212118a1dfa[0] ^
            exp_syn[44];
          Ifd9345cf219c58291c0b437aac093d78 <=
            Ib58043c04b5c4c86c1c67e57cc66dcf7[8] ^
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[6] ^
            I4a16e8e7946d9a8220304fc1be3fb362[4] ^
            Iedd7d4ea8d082b40244c04946dfb14a0[3] ^
            I13168bab2231ed22a3509142f990e408[0] ^
            exp_syn[45];
          I4f2d7bb48918ce51efe6b3b12f9f8e65 <=
            Ibc0871b3c992fd278815fdbefcd2bac0[8] ^
            I8e591d83170c8ba46d31c61935311b22[6] ^
            I07930a807994815de45864af579902c4[4] ^
            I56e1fe0c7a62589c123876f2b4e57a26[3] ^
            I280145f996e5e249788cacca7caf0095[0] ^
            exp_syn[46];
          Ifa612e6208151c616c3a0319182a96f1 <=
            I8695e1e94cbfcbe4b9eae315b042529e[8] ^
            I02b62fafd371de339f299f8aefec6c43[6] ^
            I72a2f42b727a0503d43332c0f22d5ae3[4] ^
            Ia8a468877c9f96713c8141df9205f92a[3] ^
            Ia9db6d176e9b9579a1aa5f257cd1a9f6[0] ^
            exp_syn[47];
          I9cb28a0cc6358610854c8f8d1dd3c707 <=
            I5b7caaeb34c43e66e8d095a859e708fe[9] ^
            I9c0b88a0be66d62f8ab061aeaee7e60f[3] ^
            Iea7da1f43ba202d753b0edb0be8b3fcf[7] ^
            I0ed43cf9eec83545457c57cfb6181d3c[0] ^
            exp_syn[48];
          I40bcc924f5cf1f7d587aa35267022261 <=
            I61f0c04673dfb262ef6912eb2df39120[9] ^
            Id88b9265ff08e0730e6a41abe1f80a32[3] ^
            I872f61d20baf011e867b44dc5539fc37[7] ^
            I5b74f5fc705a0406ff2376cb8ac11db4[0] ^
            exp_syn[49];
          I5238f7273b05b8b9f376314acdc6cc42 <=
            Ibeb5edab51cd6aedad9c2ecedaded6f5[9] ^
            I6330943c9295298c53e889d47c7904d9[3] ^
            I6f5c991e5fdcf56d582c6f80eb6731df[7] ^
            I14f0d3ad4fec9ca492d6b36eb29a5dea[0] ^
            exp_syn[50];
          I7137f56eeb4c4ae08bbc238db4cd3441 <=
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[9] ^
            I5686b595177e07dd5bf231a35ee41659[3] ^
            Ia5cc3055ba3365e64cf59c4d4fd3f093[7] ^
            I3a25c80d9bf7655f4ce70cf29843db43[0] ^
            exp_syn[51];
          I02335be013799e2560a98b6a82a0c528 <=
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[9] ^
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[10] ^
            Icac5a9001ee113e612e3457b4b49ee68[4] ^
            I56e1fe0c7a62589c123876f2b4e57a26[4] ^
            I260dc9154b3a9fe38b0948e807bdb42d[0] ^
            exp_syn[52];
          Id327bb65156c8307901dfcb4184bb65f <=
            Ib58043c04b5c4c86c1c67e57cc66dcf7[9] ^
            I5b7caaeb34c43e66e8d095a859e708fe[10] ^
            I9461e92a5880cb9e04fcece2ef4674f0[4] ^
            Ia8a468877c9f96713c8141df9205f92a[4] ^
            Ic49b2c150e2face8c362e33f2d87f9c4[0] ^
            exp_syn[53];
          I56331cb7b310613016958553732cdf40 <=
            Ibc0871b3c992fd278815fdbefcd2bac0[9] ^
            I61f0c04673dfb262ef6912eb2df39120[10] ^
            I6ebab438dc55ccf6c1600313891d9c38[4] ^
            I4267622319ca65909a3b40484dc74d3a[4] ^
            I714350b3b56a3249aad06d5f59fbb291[0] ^
            exp_syn[54];
          Ie3b00960f8af88a5aba7a2104dfca9a7 <=
            I8695e1e94cbfcbe4b9eae315b042529e[9] ^
            Ibeb5edab51cd6aedad9c2ecedaded6f5[10] ^
            I2fbf89398a148c47810456812dbee5a6[4] ^
            Iedd7d4ea8d082b40244c04946dfb14a0[4] ^
            Ia318eb500b8bd71048bde375c1db65a6[0] ^
            exp_syn[55];
          I7d1ef47f35b7a4c3ea2e4383732de398 <=
            I5b7caaeb34c43e66e8d095a859e708fe[11] ^
            I33a6ffad80ddf99a4d316a049078244d[4] ^
            I872f61d20baf011e867b44dc5539fc37[8] ^
            I4267622319ca65909a3b40484dc74d3a[5] ^
            Ia2c4192b1e4f180402550aebcf1dcd1f[0] ^
            exp_syn[56];
          Ibb013f036fc42687a04bdcbe2d0bbd8a <=
            I61f0c04673dfb262ef6912eb2df39120[11] ^
            I980165c1147ac5ff86619c841c6031dc[4] ^
            I6f5c991e5fdcf56d582c6f80eb6731df[8] ^
            Iedd7d4ea8d082b40244c04946dfb14a0[5] ^
            I1686a95674ecad0c4e234b8aa6e22dd9[0] ^
            exp_syn[57];
          I77eae49d321f1d1e39dd7c75829aaedc <=
            Ibeb5edab51cd6aedad9c2ecedaded6f5[11] ^
            I19df055705f322292a3601fa63f0e5f9[4] ^
            Ia5cc3055ba3365e64cf59c4d4fd3f093[8] ^
            I56e1fe0c7a62589c123876f2b4e57a26[5] ^
            I5ee21680396395f8338477fa2bb314ec[0] ^
            exp_syn[58];
          I420a4d69a077dc1996ddb4b715d63e15 <=
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[11] ^
            I3d50cfeaa4b69c09bb648b8873a6bc24[4] ^
            Iea7da1f43ba202d753b0edb0be8b3fcf[8] ^
            Ia8a468877c9f96713c8141df9205f92a[5] ^
            I005e89f0a9a9a52aec92752813a70f81[0] ^
            exp_syn[59];
          I652202a4dc8f102d29334b4811f5628d <=
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[10] ^
            I651d700a00d7004d8728bc7356f30926[4] ^
            Ia5cc3055ba3365e64cf59c4d4fd3f093[9] ^
            I0daca3ad02a67285295cd9fc330d8027[0] ^
            exp_syn[60];
          I0e33e0cdf39fc4cc99f6696e9f2784de <=
            Ib58043c04b5c4c86c1c67e57cc66dcf7[10] ^
            Ic2580cbeec8c11a19bd1e2ebc29d255e[4] ^
            Iea7da1f43ba202d753b0edb0be8b3fcf[9] ^
            I0d2ddde9edfef483482e6c177a084f6e[0] ^
            exp_syn[61];
          Ib9479328689dec62f900946e56ba0eb4 <=
            Ibc0871b3c992fd278815fdbefcd2bac0[10] ^
            If79ed5ee2b8710da0608c1e245d07d55[4] ^
            I872f61d20baf011e867b44dc5539fc37[9] ^
            I932ad562b582e2c9795f241c82901188[0] ^
            exp_syn[62];
          I2728682c0f749d1a9e8afeacdf44bfb7 <=
            I8695e1e94cbfcbe4b9eae315b042529e[10] ^
            I9497bbb4f746969a95cff948a3ee9ade[4] ^
            I6f5c991e5fdcf56d582c6f80eb6731df[9] ^
            Ifee4aa12e36833c935c54ef27b1917da[0] ^
            exp_syn[63];
          I07da3bb5f943db6271fe1867a358df35 <=
            I5b7caaeb34c43e66e8d095a859e708fe[12] ^
            I8b8b9c4777e6df3eb2b9313e69ef2c8c[5] ^
            I6f5c991e5fdcf56d582c6f80eb6731df[10] ^
            Id6f07dee3e47f39e3b43329c26f690f7[3] ^
            I51e5b79f738795719ac21c6a88711a01[0] ^
            exp_syn[64];
          I61fc44808c85a75909b9d9fd4035f147 <=
            I61f0c04673dfb262ef6912eb2df39120[12] ^
            I4a16e8e7946d9a8220304fc1be3fb362[5] ^
            Ia5cc3055ba3365e64cf59c4d4fd3f093[10] ^
            Ic7f04c065f8ff82c2288f1de77d37189[3] ^
            I4e41e628a8af629421544cb4c6f45265[0] ^
            exp_syn[65];
          Ic5075ee0ad355c20dd45ed594f2a8c3f <=
            Ibeb5edab51cd6aedad9c2ecedaded6f5[12] ^
            I07930a807994815de45864af579902c4[5] ^
            Iea7da1f43ba202d753b0edb0be8b3fcf[10] ^
            Ieb244944e7ee8236a207924f56fbc689[3] ^
            I9b2ec7db66661f7c9d85cfb1bc41893b[0] ^
            exp_syn[66];
          Ic0a651f45a502ead495cf14f97d65bfc <=
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[12] ^
            I72a2f42b727a0503d43332c0f22d5ae3[5] ^
            I872f61d20baf011e867b44dc5539fc37[10] ^
            Ie9b2be4c32334220e134e041ca8dfc06[3] ^
            I0a594a36728c7ac6244c504b8ea9c9af[0] ^
            exp_syn[67];
          Ic1c05ea22f708f620f626cc8c5ca309c <=
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[13] ^
            I04302edb2671c5bc0ca2673cd53935e1[5] ^
            Iea7da1f43ba202d753b0edb0be8b3fcf[11] ^
            Ieb244944e7ee8236a207924f56fbc689[4] ^
            Ibd943ebf64fe56a1818d2bb8b9f9f8bd[0] ^
            exp_syn[68];
          I61a18378aadae4556da501ce997321b4 <=
            I5b7caaeb34c43e66e8d095a859e708fe[13] ^
            I480a0f6d6c3eb936de10a72749f6cd3f[5] ^
            I872f61d20baf011e867b44dc5539fc37[11] ^
            Ie9b2be4c32334220e134e041ca8dfc06[4] ^
            I8c3ba90c84f9375001e727b711dead8d[0] ^
            exp_syn[69];
          Ib1fc521709a1ce2198fd8df5b41d0177 <=
            I61f0c04673dfb262ef6912eb2df39120[13] ^
            I50976b0051e84b6a42fc1dbabd7d20ae[5] ^
            I6f5c991e5fdcf56d582c6f80eb6731df[11] ^
            Id6f07dee3e47f39e3b43329c26f690f7[4] ^
            I387ca23d0e2183522ab041ec48bffef4[0] ^
            exp_syn[70];
          I1bb5511c9cda1a595c45ecde48e9ebc7 <=
            Ibeb5edab51cd6aedad9c2ecedaded6f5[13] ^
            I82e0e091fba6f79cef97eacac4b43ecb[5] ^
            Ia5cc3055ba3365e64cf59c4d4fd3f093[11] ^
            Ic7f04c065f8ff82c2288f1de77d37189[4] ^
            Ib933575f5224d414f87bc71fa7498534[0] ^
            exp_syn[71];
          I4a29c37ed36b6e12f1f8e263c92bdbc1 <=
            Ib58043c04b5c4c86c1c67e57cc66dcf7[11] ^
            I980165c1147ac5ff86619c841c6031dc[5] ^
            I8e591d83170c8ba46d31c61935311b22[7] ^
            Ibfe1bddf32fa63ea87c68de7a3af1815[0] ^
            exp_syn[72];
          I4bf02a07719402890405fb2e7b679ed9 <=
            Ibc0871b3c992fd278815fdbefcd2bac0[11] ^
            I19df055705f322292a3601fa63f0e5f9[5] ^
            I02b62fafd371de339f299f8aefec6c43[7] ^
            I719c50f9bbc66decebe794fe6ea017dd[0] ^
            exp_syn[73];
          I75bd82990cb60b6d7ccd7aa2982da7aa <=
            I8695e1e94cbfcbe4b9eae315b042529e[11] ^
            I3d50cfeaa4b69c09bb648b8873a6bc24[5] ^
            I0e0b15868b02ca52b260f17f150d237e[7] ^
            I833b0433a33dac70cb215bc8cc9f4863[0] ^
            exp_syn[74];
          Ia6d3e38249f8a1208540b68f54c46769 <=
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[11] ^
            I33a6ffad80ddf99a4d316a049078244d[5] ^
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[7] ^
            I9769761eb863e3273f9253ace4c69585[0] ^
            exp_syn[75];
          Idf548b72357ab28fd956791e84e5d65c <=
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[12] ^
            I61f0c04673dfb262ef6912eb2df39120[14] ^
            If79ed5ee2b8710da0608c1e245d07d55[5] ^
            I1fc63f388d047207a9375842c85e87f7[0] ^
            exp_syn[76];
          I50b6f2e0ef2831535ac8c18cd7ca9379 <=
            Ib58043c04b5c4c86c1c67e57cc66dcf7[12] ^
            Ibeb5edab51cd6aedad9c2ecedaded6f5[14] ^
            I9497bbb4f746969a95cff948a3ee9ade[5] ^
            I414c4d389ecc00197f2138eff0b6454e[0] ^
            exp_syn[77];
          I4003a2515229ca8eb6fefa2bef289ca6 <=
            Ibc0871b3c992fd278815fdbefcd2bac0[12] ^
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[14] ^
            I651d700a00d7004d8728bc7356f30926[5] ^
            Ibe387e8fe6f35588e028ba29cda5b912[0] ^
            exp_syn[78];
          I48672f8b83eef8c406694676746469e7 <=
            I8695e1e94cbfcbe4b9eae315b042529e[12] ^
            I5b7caaeb34c43e66e8d095a859e708fe[14] ^
            Ic2580cbeec8c11a19bd1e2ebc29d255e[5] ^
            I98191a7e6c56aae1b56e3d623004ed75[0] ^
            exp_syn[79];
          Ia14a60c9497c0faf3f1f448ff2abe553 <=
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[15] ^
            Ic2941d16ae6a5cbce70e8546a18ca4ff[3] ^
            Ia5cc3055ba3365e64cf59c4d4fd3f093[12] ^
            Icd0f5c370462670cd18d30dfc0c81c02[0] ^
            exp_syn[80];
          I0ef3962dd323e8ec64c4a881bd4b3044 <=
            I5b7caaeb34c43e66e8d095a859e708fe[15] ^
            I8e29ebe9ee25ea8ef3e52ff56fc29157[3] ^
            Iea7da1f43ba202d753b0edb0be8b3fcf[12] ^
            I15c59dc8eba10ff8eadfa6078678773b[0] ^
            exp_syn[81];
          Ie9b64c34e31dab63c03b3de4528d53fe <=
            I61f0c04673dfb262ef6912eb2df39120[15] ^
            Ic3742290179b27b9865f9d1f88d66266[3] ^
            I872f61d20baf011e867b44dc5539fc37[12] ^
            I3870d672343c002ad9c83c816fd40567[0] ^
            exp_syn[82];
          I5941476ded9f6dc25d7394f5d133955b <=
            Ibeb5edab51cd6aedad9c2ecedaded6f5[15] ^
            I9ef21ef20099af28d9a8c794f70d45a5[3] ^
            I6f5c991e5fdcf56d582c6f80eb6731df[12] ^
            Ic341b9d947f2d3ac57aa41f408214434[0] ^
            exp_syn[83];
          Ib46c78ff661ee6fb69c704d39235ffe1 <=
            Ib58043c04b5c4c86c1c67e57cc66dcf7[13] ^
            Icac5a9001ee113e612e3457b4b49ee68[5] ^
            I56e1fe0c7a62589c123876f2b4e57a26[6] ^
            Ied40f6b7847158bd08cbd932254dd6ba[0] ^
            exp_syn[84];
          Iadabc5abc7dfbc1dd747179ad7e37850 <=
            Ibc0871b3c992fd278815fdbefcd2bac0[13] ^
            I9461e92a5880cb9e04fcece2ef4674f0[5] ^
            Ia8a468877c9f96713c8141df9205f92a[6] ^
            I6ab04d323306b7290cc89ed66dbd93bf[0] ^
            exp_syn[85];
          I97a6b5f0976feceee3a5b5890d4d76a0 <=
            I8695e1e94cbfcbe4b9eae315b042529e[13] ^
            I6ebab438dc55ccf6c1600313891d9c38[5] ^
            I4267622319ca65909a3b40484dc74d3a[6] ^
            Iac4a5fdede87b021e6a8150d3bf34b66[0] ^
            exp_syn[86];
          I7217d4790fec9797a1eb8cab1ebce71b <=
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[13] ^
            I2fbf89398a148c47810456812dbee5a6[5] ^
            Iedd7d4ea8d082b40244c04946dfb14a0[6] ^
            Id92b1676e19c5818fa813d06dc9a01f3[0] ^
            exp_syn[87];
          I3dd024db4130c105a6817e8a4935de0d <=
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[16] ^
            If511a6ea6aa5cda5353658d8e192791f[2] ^
            I93da1192f27c33e21e03b9a2748774ea[0] ^
            exp_syn[88];
          Iae502e5a5ae518fb7b817afff28b7932 <=
            I5b7caaeb34c43e66e8d095a859e708fe[16] ^
            Ib0bf69cc797f330fb2546eb46d2d6f76[2] ^
            I69a0c79d41af6b6340430b8b337fb0ca[0] ^
            exp_syn[89];
          Ib8b2b1d90204af5b100379ecad20fc0f <=
            I61f0c04673dfb262ef6912eb2df39120[16] ^
            Iec7404bc79c58d4d2538fcdf659e9134[2] ^
            Ibd47f48d306ec44d94865a0a81e4f9dc[0] ^
            exp_syn[90];
          Idf0e651d0b13e167df3c0cc40d149c29 <=
            Ibeb5edab51cd6aedad9c2ecedaded6f5[16] ^
            Ie1cd04c7668d3f450c387a6c1ad778c7[2] ^
            Ia5707d1275138a5145b2a42190d95183[0] ^
            exp_syn[91];
          I89daaca029498d05ca62c095db439eb5 <=
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[14] ^
            I9c0b88a0be66d62f8ab061aeaee7e60f[4] ^
            I50976b0051e84b6a42fc1dbabd7d20ae[6] ^
            I33bc2f42d997a2963b063326eb210d1c[0] ^
            exp_syn[92];
          I0fe5a34ceda936d0924efdd07fad11e5 <=
            Ib58043c04b5c4c86c1c67e57cc66dcf7[14] ^
            Id88b9265ff08e0730e6a41abe1f80a32[4] ^
            I82e0e091fba6f79cef97eacac4b43ecb[6] ^
            Ib22e39b701614cd9986061c32adfbc66[0] ^
            exp_syn[93];
          I7876cbb2b5d8aba3652ec8b218080dff <=
            Ibc0871b3c992fd278815fdbefcd2bac0[14] ^
            I6330943c9295298c53e889d47c7904d9[4] ^
            I04302edb2671c5bc0ca2673cd53935e1[6] ^
            I9b08176fde1cd08c9d7686a659213580[0] ^
            exp_syn[94];
          If692ff56ce90d22d7af881599c54df75 <=
            I8695e1e94cbfcbe4b9eae315b042529e[14] ^
            I5686b595177e07dd5bf231a35ee41659[4] ^
            I480a0f6d6c3eb936de10a72749f6cd3f[6] ^
            I1b4e65357a818998d08b83d21584e18c[0] ^
            exp_syn[95];
          I18a7a4fe8931c79df3a69223af46c440 <=
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[17] ^
            If511a6ea6aa5cda5353658d8e192791f[3] ^
            I07930a807994815de45864af579902c4[6] ^
            Ibb865ea5891db706b7b54e5c6fa383d0[0] ^
            exp_syn[96];
          I8eec3538b8cc9c046954b6804cc656b0 <=
            I5b7caaeb34c43e66e8d095a859e708fe[17] ^
            Ib0bf69cc797f330fb2546eb46d2d6f76[3] ^
            I72a2f42b727a0503d43332c0f22d5ae3[6] ^
            I32d42cfd2d516af2e68fc2db4d5dce03[0] ^
            exp_syn[97];
          I653767e659590c1676edf6c25fc0e253 <=
            I61f0c04673dfb262ef6912eb2df39120[17] ^
            Iec7404bc79c58d4d2538fcdf659e9134[3] ^
            I8b8b9c4777e6df3eb2b9313e69ef2c8c[6] ^
            I4d0e8d475a5d2a7da24daca60f23f3d6[0] ^
            exp_syn[98];
          I5ff863be142b92dff89f7916d0d088c1 <=
            Ibeb5edab51cd6aedad9c2ecedaded6f5[17] ^
            Ie1cd04c7668d3f450c387a6c1ad778c7[3] ^
            I4a16e8e7946d9a8220304fc1be3fb362[6] ^
            Ie3850345b207e59aaaa5c944dab40b90[0] ^
            exp_syn[99];
          I49f9fd0e0719be527f2a54814dab83ea <=
            Ib58043c04b5c4c86c1c67e57cc66dcf7[15] ^
            I04302edb2671c5bc0ca2673cd53935e1[7] ^
            I4a9a1c932db30dcf04cb105a8d7384f9[0] ^
            exp_syn[100];
          I945f2476eb599844cbee0cd89038e392 <=
            Ibc0871b3c992fd278815fdbefcd2bac0[15] ^
            I480a0f6d6c3eb936de10a72749f6cd3f[7] ^
            I0ef689822226332f5feaf79fcf8f6674[0] ^
            exp_syn[101];
          Ied0c5f8a9243cd9d93672ad6cc907d21 <=
            I8695e1e94cbfcbe4b9eae315b042529e[15] ^
            I50976b0051e84b6a42fc1dbabd7d20ae[7] ^
            Ib5744c2130bb5a9d0ccdd975fdf2ff9c[0] ^
            exp_syn[102];
          I9134c7f579723c7615af60b4344efe76 <=
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[15] ^
            I82e0e091fba6f79cef97eacac4b43ecb[7] ^
            I039a7ddcb25972501d80c45c938cf683[0] ^
            exp_syn[103];
          Ie92388a9d1e71d73c07ed86e9bf6c887 <=
            Iec7404bc79c58d4d2538fcdf659e9134[4] ^
            I02b62fafd371de339f299f8aefec6c43[8] ^
            Ieb244944e7ee8236a207924f56fbc689[5] ^
            I56e1fe0c7a62589c123876f2b4e57a26[7] ^
            Ic5f36c15ebad061dfbd5301e02ce2ffe[0] ^
            exp_syn[104];
          I6804fecdf59233c6cf14409bf2f1e430 <=
            Ie1cd04c7668d3f450c387a6c1ad778c7[4] ^
            I0e0b15868b02ca52b260f17f150d237e[8] ^
            Ie9b2be4c32334220e134e041ca8dfc06[5] ^
            Ia8a468877c9f96713c8141df9205f92a[7] ^
            Idf0d9dac06522293f8d7e00a93b6bbb5[0] ^
            exp_syn[105];
          I9e777a342bf53eaba0280737ae404bc1 <=
            If511a6ea6aa5cda5353658d8e192791f[4] ^
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[8] ^
            Id6f07dee3e47f39e3b43329c26f690f7[5] ^
            I4267622319ca65909a3b40484dc74d3a[7] ^
            Id557db735a70dbb14504bc3088e8798e[0] ^
            exp_syn[106];
          Ied53820aab06b5c3423b1d878c71948f <=
            Ib0bf69cc797f330fb2546eb46d2d6f76[4] ^
            I8e591d83170c8ba46d31c61935311b22[8] ^
            Ic7f04c065f8ff82c2288f1de77d37189[5] ^
            Iedd7d4ea8d082b40244c04946dfb14a0[7] ^
            I150d31ef31093fdfc5f145d84bb35156[0] ^
            exp_syn[107];
          I24cceded372d782c67b33f3a78b16045 <=
            Ib58043c04b5c4c86c1c67e57cc66dcf7[16] ^
            I19df055705f322292a3601fa63f0e5f9[6] ^
            I7e40e6f9d82d9b9fc546672e8e8621bb[0] ^
            exp_syn[108];
          I2e78d36bca5bfb016af674c343f9c041 <=
            Ibc0871b3c992fd278815fdbefcd2bac0[16] ^
            I3d50cfeaa4b69c09bb648b8873a6bc24[6] ^
            I14133cbbfa6521c5b81477fa1c229cbf[0] ^
            exp_syn[109];
          I17a9a995de58643dbbfb78604f26198b <=
            I8695e1e94cbfcbe4b9eae315b042529e[16] ^
            I33a6ffad80ddf99a4d316a049078244d[6] ^
            I3728e31a7cf48639ce873d9135dc87fb[0] ^
            exp_syn[110];
          Iad642c4c62766e8f8bd5a1e9e73bdc80 <=
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[16] ^
            I980165c1147ac5ff86619c841c6031dc[6] ^
            Ic6be12e390bd3c25c66d9b9e7c0532b8[0] ^
            exp_syn[111];
          I96f92481be1ac6cf985b8ab387d326bf <=
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[18] ^
            Iec7404bc79c58d4d2538fcdf659e9134[5] ^
            I82e0e091fba6f79cef97eacac4b43ecb[8] ^
            Icc50e1923274729fe472ca578b68c0f5[0] ^
            exp_syn[112];
          Ie03c09039ccafb427153d2347c1caea8 <=
            I5b7caaeb34c43e66e8d095a859e708fe[18] ^
            Ie1cd04c7668d3f450c387a6c1ad778c7[5] ^
            I04302edb2671c5bc0ca2673cd53935e1[8] ^
            I4d98064f544a41b977ba945d2eecdf21[0] ^
            exp_syn[113];
          Ie7381a8294b4cdf669b9c57cfe4012b5 <=
            I61f0c04673dfb262ef6912eb2df39120[18] ^
            If511a6ea6aa5cda5353658d8e192791f[5] ^
            I480a0f6d6c3eb936de10a72749f6cd3f[8] ^
            I12f2a9f1e3e715d7e684ff39dd7942f0[0] ^
            exp_syn[114];
          I61c9e3f8e42f869f4c9c1386325100b3 <=
            Ibeb5edab51cd6aedad9c2ecedaded6f5[18] ^
            Ib0bf69cc797f330fb2546eb46d2d6f76[5] ^
            I50976b0051e84b6a42fc1dbabd7d20ae[8] ^
            Iaa4e3c53a0d55e8f42f60ff40893427e[0] ^
            exp_syn[115];
          I24c5b2de59eb1f43fe1efe687231c4b7 <=
            I8695e1e94cbfcbe4b9eae315b042529e[17] ^
            I9ef21ef20099af28d9a8c794f70d45a5[4] ^
            I26aae317b0b320df86ca4004f64aab88[0] ^
            exp_syn[116];
          I43d43acde5f831fc32b7bf5f10b9b3a9 <=
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[17] ^
            Ic2941d16ae6a5cbce70e8546a18ca4ff[4] ^
            I9344825cc2e5864f691043a1f94f86a4[0] ^
            exp_syn[117];
          Ib06e93161fc8ca3be232f4261b04feb1 <=
            Ib58043c04b5c4c86c1c67e57cc66dcf7[17] ^
            I8e29ebe9ee25ea8ef3e52ff56fc29157[4] ^
            I82988c3879c1de76fe2140c469f6a4c1[0] ^
            exp_syn[118];
          Ia0dd00f83afc805036f2c6a0e38f725e <=
            Ibc0871b3c992fd278815fdbefcd2bac0[17] ^
            Ic3742290179b27b9865f9d1f88d66266[4] ^
            I6bdd8334512c7c6a3226ebb4e928a270[0] ^
            exp_syn[119];
          Ib0a0f924fe3757a1e0aade7017ad9277 <=
            If511a6ea6aa5cda5353658d8e192791f[6] ^
            I04302edb2671c5bc0ca2673cd53935e1[9] ^
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[9] ^
            I07930a807994815de45864af579902c4[7] ^
            I0debec6ace7160558cce7f111dd1bea6[0] ^
            exp_syn[120];
          I1ca949071d734d230cdb8adda46c9d79 <=
            Ib0bf69cc797f330fb2546eb46d2d6f76[6] ^
            I480a0f6d6c3eb936de10a72749f6cd3f[9] ^
            I8e591d83170c8ba46d31c61935311b22[9] ^
            I72a2f42b727a0503d43332c0f22d5ae3[7] ^
            I8ee02e65ce9183683f0f3168bfd755c5[0] ^
            exp_syn[121];
          I40170922c652fa7fa42abc6f580b5e3d <=
            Iec7404bc79c58d4d2538fcdf659e9134[6] ^
            I50976b0051e84b6a42fc1dbabd7d20ae[9] ^
            I02b62fafd371de339f299f8aefec6c43[9] ^
            I8b8b9c4777e6df3eb2b9313e69ef2c8c[7] ^
            I80e6d2c9c5f7b6bc6bffa063c4959115[0] ^
            exp_syn[122];
          Ib1ad0b531ac9028971d68f533e7ae566 <=
            Ie1cd04c7668d3f450c387a6c1ad778c7[6] ^
            I82e0e091fba6f79cef97eacac4b43ecb[9] ^
            I0e0b15868b02ca52b260f17f150d237e[9] ^
            I4a16e8e7946d9a8220304fc1be3fb362[7] ^
            I0f21fb041239a7a8895c9506f2754595[0] ^
            exp_syn[123];
          I0ab0170c7ceffbb58377b65d2ad92093 <=
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[19] ^
            Iedd7d4ea8d082b40244c04946dfb14a0[8] ^
            I8ce37a8e81b54043276835c11e394df5[0] ^
            exp_syn[124];
          I9ac68f228a93bbf4aa4a559b1364e42e <=
            I5b7caaeb34c43e66e8d095a859e708fe[19] ^
            I56e1fe0c7a62589c123876f2b4e57a26[8] ^
            Idf7d1f78735ce1e9695d99a532a7726e[0] ^
            exp_syn[125];
          I375c5f7eac92d853e85e0606011f3fb0 <=
            I61f0c04673dfb262ef6912eb2df39120[19] ^
            Ia8a468877c9f96713c8141df9205f92a[8] ^
            I96a552ed2d18c0ba3fc6cb6d6b6a0f44[0] ^
            exp_syn[126];
          I94f9b1f2e63748c21ec7222c9641366a <=
            Ibeb5edab51cd6aedad9c2ecedaded6f5[19] ^
            I4267622319ca65909a3b40484dc74d3a[8] ^
            I3c76936e8e3467378210a13645a401d4[0] ^
            exp_syn[127];
          I55500c1d85c4970932be67cc5cd2e023 <=
            I8695e1e94cbfcbe4b9eae315b042529e[18] ^
            I04302edb2671c5bc0ca2673cd53935e1[10] ^
            Id6f07dee3e47f39e3b43329c26f690f7[6] ^
            Ic9a1d599fcfd5dd51265e5d0989719b6[0] ^
            exp_syn[128];
          I36b487cd1a57a3a503e587fdefbb19e4 <=
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[18] ^
            I480a0f6d6c3eb936de10a72749f6cd3f[10] ^
            Ic7f04c065f8ff82c2288f1de77d37189[6] ^
            I60156470e631268c392040d3c5582eca[0] ^
            exp_syn[129];
          Icb5350e8c55a2adb370078a7575e28f8 <=
            Ib58043c04b5c4c86c1c67e57cc66dcf7[18] ^
            I50976b0051e84b6a42fc1dbabd7d20ae[10] ^
            Ieb244944e7ee8236a207924f56fbc689[6] ^
            I821126d1516ad7e8191a7b2a3b5e4b47[0] ^
            exp_syn[130];
          I8a7a31327c9e4cbd88ce39fea8971caf <=
            Ibc0871b3c992fd278815fdbefcd2bac0[18] ^
            I82e0e091fba6f79cef97eacac4b43ecb[10] ^
            Ie9b2be4c32334220e134e041ca8dfc06[6] ^
            Ibe72e9f6d2c3cbbcf98f6b5aa6a4f93b[0] ^
            exp_syn[131];
          Ied069655ed3775819d0bcb722d6d0488 <=
            Ib0bf69cc797f330fb2546eb46d2d6f76[7] ^
            I0e0b15868b02ca52b260f17f150d237e[10] ^
            I651d700a00d7004d8728bc7356f30926[6] ^
            I1e8b6306d2dfde4a36ee9b9c2caf1c85[0] ^
            exp_syn[132];
          I78a5fc80d42e8db1b56cce5f4c97e325 <=
            Iec7404bc79c58d4d2538fcdf659e9134[7] ^
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[10] ^
            Ic2580cbeec8c11a19bd1e2ebc29d255e[6] ^
            I48ed92480f457fc3cc2ff0dd7d177a10[0] ^
            exp_syn[133];
          I3ade7e345432319c1a9c91d4068b3ec9 <=
            Ie1cd04c7668d3f450c387a6c1ad778c7[7] ^
            I8e591d83170c8ba46d31c61935311b22[10] ^
            If79ed5ee2b8710da0608c1e245d07d55[6] ^
            Iaed28d88a651f0151501ec4ea6ee3346[0] ^
            exp_syn[134];
          I88aed46f6dad7a81006562a720670654 <=
            If511a6ea6aa5cda5353658d8e192791f[7] ^
            I02b62fafd371de339f299f8aefec6c43[10] ^
            I9497bbb4f746969a95cff948a3ee9ade[6] ^
            I9d94d9b5414662de841443d7866e66b1[0] ^
            exp_syn[135];
          I79e574dc9c7e18b695c9a2619b71b995 <=
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[19] ^
            Ie9b2be4c32334220e134e041ca8dfc06[7] ^
            I4267622319ca65909a3b40484dc74d3a[9] ^
            I870b8a3b11be215a8704ba05568f05e2[0] ^
            exp_syn[136];
          I800ef583bec1d46d3d4ffdea6b312ef9 <=
            Ib58043c04b5c4c86c1c67e57cc66dcf7[19] ^
            Id6f07dee3e47f39e3b43329c26f690f7[7] ^
            Iedd7d4ea8d082b40244c04946dfb14a0[9] ^
            Ia8bbf21e040b326058a9acb7d198a835[0] ^
            exp_syn[137];
          I56cc5cd6d0a5a4e4601fd48e838fdaf3 <=
            Ibc0871b3c992fd278815fdbefcd2bac0[19] ^
            Ic7f04c065f8ff82c2288f1de77d37189[7] ^
            I56e1fe0c7a62589c123876f2b4e57a26[9] ^
            Ie852f207c8f537621b080ffa0a89bfdc[0] ^
            exp_syn[138];
          I21047a3955b8b89bdb9013d571b2bd0d <=
            I8695e1e94cbfcbe4b9eae315b042529e[19] ^
            Ieb244944e7ee8236a207924f56fbc689[7] ^
            Ia8a468877c9f96713c8141df9205f92a[9] ^
            If53029b05bea46d656a6ef72fb6d6642[0] ^
            exp_syn[139];
          I56eb529a34b484cd20e29958cd6878eb <=
            Ibeb5edab51cd6aedad9c2ecedaded6f5[20] ^
            I04302edb2671c5bc0ca2673cd53935e1[11] ^
            I872f61d20baf011e867b44dc5539fc37[13] ^
            I8e8a740d09e000444ba1f4931b5cccf4[0] ^
            exp_syn[140];
          I74588df6399af2c1112e3fa557e89e17 <=
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[20] ^
            I480a0f6d6c3eb936de10a72749f6cd3f[11] ^
            I6f5c991e5fdcf56d582c6f80eb6731df[13] ^
            I46605d823e06af5485e50b256b5c3f22[0] ^
            exp_syn[141];
          Ic8eae1a92f46db040eb22d726c3a0e6d <=
            I5b7caaeb34c43e66e8d095a859e708fe[20] ^
            I50976b0051e84b6a42fc1dbabd7d20ae[11] ^
            Ia5cc3055ba3365e64cf59c4d4fd3f093[13] ^
            I38344d68127f5c035193bb9030ce4d4d[0] ^
            exp_syn[142];
          I854a15bc7e9728b01c9a1960f6248dc9 <=
            I61f0c04673dfb262ef6912eb2df39120[20] ^
            I82e0e091fba6f79cef97eacac4b43ecb[11] ^
            Iea7da1f43ba202d753b0edb0be8b3fcf[13] ^
            Iba9f33c08db89a7f120cc1e3eaf05dec[0] ^
            exp_syn[143];
          Iae332cfd000fd0529684ab787041b5dc <=
            Ib58043c04b5c4c86c1c67e57cc66dcf7[20] ^
            Ie1cd04c7668d3f450c387a6c1ad778c7[8] ^
            I8e591d83170c8ba46d31c61935311b22[11] ^
            Ibde51eb91b3ca50a8a0513c94bd7be15[0] ^
            exp_syn[144];
          I70148fe95244eebf7f0ec953703398de <=
            Ibc0871b3c992fd278815fdbefcd2bac0[20] ^
            If511a6ea6aa5cda5353658d8e192791f[8] ^
            I02b62fafd371de339f299f8aefec6c43[11] ^
            Ifb94196d1653a0166567e170f06ec0db[0] ^
            exp_syn[145];
          I24ee2d953e65fefdc73b3d3c4c0ddd05 <=
            I8695e1e94cbfcbe4b9eae315b042529e[20] ^
            Ib0bf69cc797f330fb2546eb46d2d6f76[8] ^
            I0e0b15868b02ca52b260f17f150d237e[11] ^
            I9cf7557e2cac4532a77fcb212712db0f[0] ^
            exp_syn[146];
          Ie3a5f8eec283fd4f682b5d0f909b051c <=
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[20] ^
            Iec7404bc79c58d4d2538fcdf659e9134[8] ^
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[11] ^
            I3159d7faeee1a904c409bde1967d2c21[0] ^
            exp_syn[147];
          I781d986d7fd6c2fec3a8cf3f29545174 <=
            I651d700a00d7004d8728bc7356f30926[7] ^
            Ia8a468877c9f96713c8141df9205f92a[10] ^
            I35dfb5ece5e04504d6e74739ae99c9cc[0] ^
            exp_syn[148];
          Ib4db8131350f8605e00907234aff901d <=
            Ic2580cbeec8c11a19bd1e2ebc29d255e[7] ^
            I4267622319ca65909a3b40484dc74d3a[10] ^
            Iabff939ae4acf7d7b038e028c29b6166[0] ^
            exp_syn[149];
          Ie093f0750b60d3aed75705637933f34c <=
            If79ed5ee2b8710da0608c1e245d07d55[7] ^
            Iedd7d4ea8d082b40244c04946dfb14a0[10] ^
            Ia14159444578c6dc88f2d5ea0317774b[0] ^
            exp_syn[150];
          Id2fba7c1b3dc7a75a5e0d90494d56962 <=
            I9497bbb4f746969a95cff948a3ee9ade[7] ^
            I56e1fe0c7a62589c123876f2b4e57a26[10] ^
            Ie2306a5c441d621388b73195027fc118[0] ^
            exp_syn[151];
          I9ecee74c445711a376133636ef414666 <=
            I5b7caaeb34c43e66e8d095a859e708fe[21] ^
            I50976b0051e84b6a42fc1dbabd7d20ae[12] ^
            Iea7da1f43ba202d753b0edb0be8b3fcf[14] ^
            I700a0fbf81e57d4970ce07090ec4f2e2[0] ^
            exp_syn[152];
          Ifb3cf6b88835d27220df837682c4dc93 <=
            I61f0c04673dfb262ef6912eb2df39120[21] ^
            I82e0e091fba6f79cef97eacac4b43ecb[12] ^
            I872f61d20baf011e867b44dc5539fc37[14] ^
            I6007914b3fb3011c3ab2f9a9d7794ab2[0] ^
            exp_syn[153];
          I386fbb3bd550891d682e137044e8773a <=
            Ibeb5edab51cd6aedad9c2ecedaded6f5[21] ^
            I04302edb2671c5bc0ca2673cd53935e1[12] ^
            I6f5c991e5fdcf56d582c6f80eb6731df[14] ^
            I2096f40fe62e9d6f1ff96f258ffdbe33[0] ^
            exp_syn[154];
          I7ede7d2e1c2730b3b71340b11e880f5b <=
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[21] ^
            I480a0f6d6c3eb936de10a72749f6cd3f[12] ^
            Ia5cc3055ba3365e64cf59c4d4fd3f093[14] ^
            I93d8b7a24702bacbfc528242991516a9[0] ^
            exp_syn[155];
          I64c65fad4a7d958d625c783626808175 <=
            Ifeb6f8e9d7d86fb01ee8faed3bad6d6e[21] ^
            I0e0b15868b02ca52b260f17f150d237e[12] ^
            Id6f07dee3e47f39e3b43329c26f690f7[8] ^
            If0863fae91b2ec980ebdb26cfc90ae2e[0] ^
            exp_syn[156];
          Ib2e0cd0a2b51c3a265bdd20834c0ed2d <=
            Ib58043c04b5c4c86c1c67e57cc66dcf7[21] ^
            I3c0b6f53f0a5cda5b6758b2ee2c83b92[12] ^
            Ic7f04c065f8ff82c2288f1de77d37189[8] ^
            I9ec29a319384efd562c2337e1857cb4e[0] ^
            exp_syn[157];
          I67be0b66c8d0680eb23290a4b3885af3 <=
            Ibc0871b3c992fd278815fdbefcd2bac0[21] ^
            I8e591d83170c8ba46d31c61935311b22[12] ^
            Ieb244944e7ee8236a207924f56fbc689[8] ^
            Ia56ecc024eae608d7de1509d75139dc2[0] ^
            exp_syn[158];
          I01148401f7d058614dc1ae6ed3c8bd94 <=
            I8695e1e94cbfcbe4b9eae315b042529e[21] ^
            I02b62fafd371de339f299f8aefec6c43[12] ^
            Ie9b2be4c32334220e134e041ca8dfc06[8] ^
            Iebcd65ea41cd38bfe3c8577277809acd[0] ^
            exp_syn[159];
          I3394319c370daf6102be00d938d55769 <=
            Ib0bf69cc797f330fb2546eb46d2d6f76[9] ^
            I651d700a00d7004d8728bc7356f30926[8] ^
            I4267622319ca65909a3b40484dc74d3a[11] ^
            I75be12b14694ebcb5aff6e5d3e576315[0] ^
            exp_syn[160];
          I24d6a334dd15ccdea558f32cd029e6d1 <=
            Iec7404bc79c58d4d2538fcdf659e9134[9] ^
            Ic2580cbeec8c11a19bd1e2ebc29d255e[8] ^
            Iedd7d4ea8d082b40244c04946dfb14a0[11] ^
            I8e06fe414cd04103baf3882771a63e2c[0] ^
            exp_syn[161];
          I3a41f68bca2d7edd1f5738c4fda8e73c <=
            Ie1cd04c7668d3f450c387a6c1ad778c7[9] ^
            If79ed5ee2b8710da0608c1e245d07d55[8] ^
            I56e1fe0c7a62589c123876f2b4e57a26[11] ^
            I0fe8574049166c363c7cc816b1435009[0] ^
            exp_syn[162];
          I9ef1784d165492f3482d14f475732451 <=
            If511a6ea6aa5cda5353658d8e192791f[9] ^
            I9497bbb4f746969a95cff948a3ee9ade[8] ^
            Ia8a468877c9f96713c8141df9205f92a[11] ^
            Id5f435c07240d5fe4a0e48c8f25ad0b7[0] ^
            exp_syn[163];
          I9d9378337a77515a4e8d04fb88938808 <=
            Ibeb5edab51cd6aedad9c2ecedaded6f5[22] ^
            I480a0f6d6c3eb936de10a72749f6cd3f[13] ^
            Iea7da1f43ba202d753b0edb0be8b3fcf[15] ^
            I1ae21e0db88f955c4f08f6d52f58974d[0] ^
            exp_syn[164];
          If0e20ef9aa69b77ae0e58ca3dfc9998f <=
            Iceb64ab2ff8a2e0dfdb74803811d4cfe[22] ^
            I50976b0051e84b6a42fc1dbabd7d20ae[13] ^
            I872f61d20baf011e867b44dc5539fc37[15] ^
            I92efddd59e1ea92902a295c0b8385c68[0] ^
            exp_syn[165];
          Iec2cb48bb1b58f268bf164d5e8a8120f <=
            I5b7caaeb34c43e66e8d095a859e708fe[22] ^
            I82e0e091fba6f79cef97eacac4b43ecb[13] ^
            I6f5c991e5fdcf56d582c6f80eb6731df[15] ^
            I56948ad2b2cc245bb1003fd71ae5f899[0] ^
            exp_syn[166];
          Ia4ae7c98720d43a604f28dfc5dd67d50 <=
            I61f0c04673dfb262ef6912eb2df39120[22] ^
            I04302edb2671c5bc0ca2673cd53935e1[13] ^
            Ia5cc3055ba3365e64cf59c4d4fd3f093[15] ^
            I5fb5081b7a2da89115c0080b0967974d[0] ^
            exp_syn[167];



          I5033323484d90d6bfbe03749019fc6dd <=
            I1a632a3e06ad738d5865acc77e204f48 +
            I71b93abe4b20e6a17ff17e0f33ac2ca5 +
            I9184110e3e9b8614460fc0abe5fff2d9 +
            I535cad8c919a4330257eb5b4bed61b3a +
            I7ea8fe50c45e213f3257060e2813240b +
            Ifec9abca21cf476b70e0befa3926b46a +
            I7c191c2c2be09886d0f31e4368797afd +
            Idd01d014f0469f893305057ae3f4cb2e +
            {MAX_SUM_WDTH_LONG{1'h0}};
          If5dad13ac41b3034bdb034bc86c9b348 <=
            I3f59174b3764a0b0741462024be9fb92 +
            I0e112f1d4e9c934a118f79f3856744a9 +
            I65708fb59e90bb79b8107da619fe63eb +
            I0fc42ce9cc31d781ea3013318c25a571 +
            I8bc3210e86a523accdbeefe7e72ee4fc +
            I597c3f5c14e235f90dc8c796bc3e931d +
            I07d68462362d8453e83570cc793c55db +
            Ife6be241bc50560a14f97650e5cc2959 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Iac428f9f798618e1ef495c626c41892b <=
            Ie04ce30f26a4ef1ee5b34474368dbac7 +
            I546657528d591e8bb44c32fed7707af5 +
            I0ace1d51fdee91f8f3826a945c4e66a4 +
            I8dbe6497a8deabcc60783bfe7548d0fb +
            I9a57f2f03cf8a154c3a7d48ec089306d +
            Icda9a86a25dbe516a93b46fe487029e3 +
            I64ae3cd6f36b8bde29cd3e1fcba7bade +
            Idc4171a40dd2470e852af37a461013c7 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I5a6427c8f18b36d2ea18fe60a0831ef1 <=
            I43864225be03ea8e9379eb28dfa6c599 +
            I70e68beb262fbdeba621b3794adf9f84 +
            I656852be6f5b3542862e0f68d48be518 +
            I041f9455435bfa375395eb330a34993d +
            Iac48d2ccf6c6e0c555e874ae77123f2e +
            Ib76e892d1a1271844338042381b5690b +
            I45b64b2b963963d2d0a8318133941f1d +
            I8435e69bc1ff06e7edfabbee7b9aa49e +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Icc29441eac6ca7a138d45743d37505e3 <=
            Ibfee0b4ad5cdf16e88fcf469c5e031e9 +
            Ib2afdf9534deaae465d99b7e377788bb +
            Ib6cdbbb765694d822639b7c8fbfc50c4 +
            I8dddcade21ad3bb330c1c25970c32b73 +
            Ib63574478126e6ee30a388d9648cb548 +
            Ia1aedd38250e76763aaee3de2f832b3c +
            Id5ddf5331aba567aaf5b7eb88b31a52e +
            Icb158c031d434cb419c15e0510511231 +
            I79444eef1875b6ad1a0675b66392ff9d +
            Ib88c884e54d6e6ecf5ac015bc304e4f3 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I0e7754dcbc04a4850e052ae4a2fbe328 <=
            I31cb0c699cffcd2fedfbed0e1b86490e +
            I4363ca6b3d9ca9863f70958aa7c23777 +
            I25eb943ea517a4827efb1e797bfdc4f5 +
            I490996026af34eba5bcd8d553af818eb +
            I9d8f8c1792427975a9e7024041f59be9 +
            I452ba61d5fb5c7ead1824dade4bd7801 +
            I7e36dcae438a712fca2320117b7e3356 +
            Ifc527b6af9486df7f52d7eb9637c671f +
            I1062442edb2bff727ca6283c8270bf28 +
            I2959f2dc554e599d675eb6912757e413 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ia30c019ed8ce395556494a92e7b42a92 <=
            I4d4ec5540257040d10182ed478a71918 +
            Ifef870b405335975988b58b2273d4e1a +
            I9e0a36d0be66b4c02b03e5b75b686226 +
            If404a00ab81d6ebbc0dbdf4aecdce389 +
            Ic6f40833f5f6284c9015304fd3fc00f0 +
            Ib8664a2abe9d6326d6e45bb2a7ad59d0 +
            I36ed1a0d0d618f90443fbea17b7c97ec +
            I397a69dab323c7148b620dd6fe0b0c51 +
            Ifae488cb68d95ea517376319eb11f1bf +
            I10f045edf47784a91a5599494c2d3de2 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I9799695ea8244992a6694eaf5c8ae64d <=
            If0c2d002c315b21e11ae776bb48c9338 +
            Ifbe29365e7035c78af9f42902b0d303e +
            I6922b510e432e06d209095bcc6297e7e +
            I31bf4597a3b776962f5c820378254065 +
            Ic3e6e38a2986c7f14fd0db2246367a1c +
            Ia1d9dee7a9821283498d17de0cfacb32 +
            Ibac0851ce1a3c23f18b072d263afff36 +
            I53971b75cbd7ebc74b579776a6ea4778 +
            Ibeff607ba15fd8ef504224a9c1d102fc +
            I4ae2f2330a8ee7d5626499f2a030c7a5 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I4524cd664b4cb41f642c675fa484c84b <=
            I8da7e01f56dc9a70eb6b3f110dc005c2 +
            I005e8b590924f9486cb23191d35c9797 +
            Ic1f6842b4f246d624d91daa6ada10ca9 +
            Ief90f8a8efca2b06eff0d4cba1cbb342 +
            I0f46a17f14ab18e6338aa3d06678b0a5 +
            Ia3bfd86e26efbef2cf6bb72be7ac1453 +
            If6f5efee5e1f9709d86bf28cfb741955 +
            I60520c850a95b893528569c4069bd677 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I64e959d80af111ed2fcd54a5407d21bf <=
            I18e548b082364c75686f2b7ad2ef46ab +
            I6e4ae763dc4e8aa8afc4599de96c75d3 +
            Ic8759e2f58848b33082bd1b02acc9c0b +
            Ibdaa6d215d34aa0cc27d5234da6fd991 +
            I0f9bc36c9d40290f83489aac3d674924 +
            I9a2bba3f62de5f750dc8161a488dc331 +
            I898d1b59aab3d5d4adce8ec3c0e14a0d +
            Ic92ab3dac1a151d6ff0b4e0c21003eb0 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I3e0da4bcbab4804b5397fb3aa2c94f51 <=
            I3a4a965f22487553dec2a3e8e7836264 +
            Ie7bf11bab3d601fd0a6e3eb415e263c8 +
            I6eaffd980e4d77fdbda5e63bad9489d7 +
            Iac4b8906947fc90bfe76cee2f1d4c4ab +
            I612a41511db375f10f3c2b10d13edb24 +
            Ia6a78664c080829664158f53ba330312 +
            I6a81b4485598387e4656c35e83866209 +
            Ifb09b84f9681c7bc28ffd562b633ffd9 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I3740b30d31f3c61d93a14a46e3199c4d <=
            Ibed5004d869a01005768ba694c2234d6 +
            I91c2f3cdd7cc98a60090ec6e46d52ae7 +
            Ic902e09b33db1b919c102f7971cdef7b +
            I1eef40a71c8d1e2da9802929a5347e90 +
            Id58474582f209a3859f65a447fe99191 +
            I1939152ddbede923cde577984e0aa743 +
            I4aa98503fc71292d42dba1cab6db952f +
            I8ce945d9f70bb317064a8d2d4eafd2d3 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ibf0a30abfec9031737eada436ac1a0d4 <=
            Ica3d4ebff001fb6ee69a66eb898eb5bd +
            I99ff3922e018c409dc8ce5f3503e3c56 +
            I58a490344f87b4d5bb319e3e85ba9278 +
            I58361fb97f1b5aff0a2751d35c8da672 +
            I581eb136fdd08302e02c1fafb5d5c90b +
            I91893028c4409cfeceeb7976815b2d31 +
            I19032091a26dfdfffff60818041ec79e +
            I563802213afb6abe2f6e8c6f4d1e5b08 +
            I4ae59dd2f57bda295e11b077e8668f1a +
            If525ac3dc97e3187e036d70e9984939d +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Id36e8953a02400a5ab1f4dfdb0422e6d <=
            I4254f2987cd014ed703ae18e9963e585 +
            Id6551b6b053952162b90792ab73a1a49 +
            Ied41909cd443432dafadba42672151c1 +
            I74a7b85ddacad06ab1c6b0db9b084bd3 +
            Ic4501a8a1fb34c30a97e18a0ab189e3a +
            Idd8643af2515f65fd9a1dfe66494ccf2 +
            Ic9e06a355beabfacc053ec48f17f49de +
            I31d94aae2e3721045fe850d84dd2225a +
            I71da7e172b2b967040b6e6d02ef9949e +
            I3da241c7f221413abfbf1b4384bfca5a +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ica71108a53bfcfd1892b4d03ef68110c <=
            I8c5f98353b5b082dc3cf056469945a08 +
            If8865fee7dbf593b34ea54692d947f10 +
            Ib5334df42ee8f1574e41cb30b903fae9 +
            Icbc12ab47f586b12402ae5d4361c967d +
            Ie8644d7edbadf19937c399cf275946e5 +
            I2087576fbc15119bf5d9e8afa2603b69 +
            If1ec4241fd12255369f72b3f3310b6e7 +
            I401ab1ad994f5018061a3f57d3a51ad1 +
            I2ba16a10a82c20d54c776a9804ee50e4 +
            Ib55b0e4c45ebbdb605f0ba9d62bff21c +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I7c97629ec6e594f9b2160815ddd133cc <=
            Id8c36004ae8e550569a491f6b514945a +
            I840a1a7c0bf49f4f42499b33f32fa02d +
            Id769d4a92f5f6da262ce0521e5509368 +
            I19875f52f79482b477f1febaa7e97090 +
            I3f2507530dd648814af0964f7da11d35 +
            I8b5d10c412daccdcb07645bf239d61bd +
            I3a09554ca009781e28ef1b3ea70d39ad +
            I37e5c3118e8536e37bd797aeaa92476c +
            Ifbcebda2bb0ce58a0e1764c392a816df +
            Iaed105b99eae5b078521e3a94d8a79b7 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I4823c8239ace86dc399e906c1b5a0d74 <=
            I2a2d014f94d7a3b9fb3024a3e9107a73 +
            I9aa11f30712f1779339b985212a7979c +
            Id15c3bdce785df234c68432ccec8f959 +
            Ia0e77e9544481aa0f56dfdb6eb253137 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I10ad572ca72c2ea991487c39f7eabd7b <=
            Ia4b2db3d48f946b0bfd0be0e32d7518d +
            I111ac0aadbdd3e4479ca0786491a7b08 +
            I7caf8c7496dd96c1ed08e98b415f5775 +
            Iec0d7ea31e0f1a75b15121090dcf1e11 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ie9f3fd3a6d16316e55addbe0e336519f <=
            Icc5d7bcbd7fcdb5092e6d8e18f6de6ec +
            I27951ef3d612004abdc639662807426b +
            I6c9ae8b8191507f908c27bbde53bf2d5 +
            Ia98bb3648ce3719b1c31ce0f41121c63 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I07965bca84276dd56da1af98e64b0adc <=
            I5e0d6b44474a226ab2ce916a6d46072a +
            I9068cca0de6ecff56ca542d0998fcab2 +
            I9cab38b69794ab661e12750cf69c822c +
            Id9c8055ef530f2cb8096cb7bb2af55a4 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ic2ade31b8bcf68c4dcc1a371ff14074b <=
            I5bab5ae46114c487f67b8e779d7461df +
            Ib3ec015a3d43d46e0b7142b21a81cfee +
            Iee0e45914c52a357e1e32922299d6937 +
            I1684820afb9d9cec38cfdfcd6ca8b36a +
            I25888aa2135fc403ca9eac4df634549a +
            Ib9081d438413a627f5b16f68c2eabb80 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ic0edcf240048fbfde4e938c3e4c5e281 <=
            I4d908bbe633c193cd9fc93dd33c60bd2 +
            I65928407b1d5447dbc815cd2d2e7b37d +
            Ic7855ca956651bd368cbdde7ec93ba6d +
            I7a6ab9e700bd94208ab6528af413f3a9 +
            I7fc6e2aecff5bd691872d1e10a39103b +
            I9c5bf5451736358f8c84e150004fa5a9 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I8b42e89ff5f780d4ef8cd1cd5c99ef61 <=
            I83cec264bd378f1dc23f87e439e7310e +
            Ib83242b57ab050b0e5f9bdf91fa118fb +
            I8ab7efc436a0f2cc3efbc299a0ddf914 +
            I9b1390839ee2b9ba591e3873e967c8e2 +
            Iec936eeebd1f8c95307bd8705e6def81 +
            I377933518c3807edb71f648c65ad5c85 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I70b1b8521b36920707e95fc9418eb8a9 <=
            I0c53d8d6a5b92960e29fc31cf456c23b +
            Ice4f4ba8bb3381c8846941d5d5fe4534 +
            I2b0b168ce4fe8aa4a2e7cb69fe532aa3 +
            I2e14fb1e667e967ab4c116e0c7438aec +
            I24180fba17c21bacefa8a4514e4b685c +
            Icec98d794a64752081fadfa74308fad3 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I4fb1c32a62cbbaeb585c6564a3c938f9 <=
            I45373bff54eccf8137da2931d841934e +
            I3934ed7170967ff3852944cc39ba1de9 +
            I17e818b67440efaba9a5d19e7467bf85 +
            Ia5b779ef95333736b08f63770900e275 +
            I83bbe6fa947f9f909e1a6785ab31901f +
            I7bbe4d0a7d61d3f7da346de71b9a3a5f +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Iefc37daeec14e14ef2fe0716f73109dc <=
            Ib14733d3585dbf7f196cfc068e9508f0 +
            I3e8d26ea83937cae01aadf1092c59bdf +
            I0fb60c4f56f6d7b4007cf0dae39f4573 +
            If3bdbb4c20efca0c5af78614b4271ed1 +
            I632ffd09a9091335b3aa91ab2a8f1cce +
            I197c05f74bf7fb8d44124d40bd7c6563 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ibd15f164f6d2ac9e5721a21464bc2c5c <=
            Ied7e494fb288f78d110ed06662f1926a +
            Iefe423653d454e21324a6857b52f98ac +
            Ice8a82bdd966719098a8d5f2a826f73d +
            I3a47540f34ce47bcfa1da66cc4e6e088 +
            I49321308413cb4dbe5e6c01ba5b9023c +
            I92acc55d81ec6e02880337b0a451ae21 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I951dfff9507bb70214d48e03a0ebb3a7 <=
            Ib16c6096ce80e2f15a5ccea145e28510 +
            Ic57a2627a194099105a2908a41feddfb +
            I4481555c402ba99bee05658ba6017984 +
            I9c68bfa3b888b6a6d41e38e674578284 +
            I6332af145d560e3f22a4a88106749f98 +
            I35c0ca76b28cd2f9355276b5d2f29ad4 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ie78e30b2a2eda75d0df7d10fd67b5e36 <=
            I8cb171677016e4309034dc5d83981a48 +
            I4d1ba6ee8fb9505ba3b58b2b7553245b +
            Ib849494e5087777f646ee0947b4f634a +
            I283331db80e6d0891b13dc55e6a7d76c +
            I0c1e4d400520935c5c78b792a9d554ba +
            I29da0e5661f29bd8493c19885c998582 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ia0b83a372dd4115dc4d61eb8ff0811b9 <=
            If5b3850da967f6f3d7a71d680341ad1c +
            Ic690477b1672dea4905a5e1c92b47366 +
            Ifa67d343acc6f3ec50c2b01fc26b4374 +
            Id27560fb44b4f2fda98d47e9f20d6898 +
            I0807a826e91f92ef279ccf0b6512a428 +
            I9426c8c1b4d988d5cd7d89a7aed4f8fc +
            {MAX_SUM_WDTH_LONG{1'h0}};
          If5c5bcbbea01aa22f242b913f0d01929 <=
            I7be8b2f8a9fe8e13001c2a1fce4a8a3f +
            I90a4190941651d885d04deb86a163365 +
            I24b4c998d19ae97f7178e37f75c77d06 +
            I0c121fa3e9e6e0e2e8291a594d6b4ceb +
            I4319fa23d59f4e690e31fb7e3a823d17 +
            Ibd010f15e36194cbd2ce9f01c98a2b6f +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Iccba58cd3519fb4cc75a61b50da1d562 <=
            I223151b6414d9979d71023053dd3f5e2 +
            I6d6a242cdfadfc97fe656510bef73adc +
            I338400586daa58006c0a3dcd82ea8f4a +
            I202c385beeccee309104b66f8f096b2c +
            I05a812cd935867d1e417c64c26ea0952 +
            I7e86ab53e6d9647b230a94e076831ba2 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ibc0999e4d0b3cc2650f9348b8c204b14 <=
            I0e7ca2d6470b9bfc6a1ca6143b468507 +
            I0aa5522190c741b7df4c4d7d34e46987 +
            Icf7630b6002db2f9b59d5323d6cc8105 +
            Ia0ecfaedbc1d546d484978fd50096d10 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I2aeff1fb4b839a581acaf26f90f9113c <=
            Ib9322ec1d3866ba3cb42e96b5ff5cfb2 +
            If4d030e5858f325debc6f37abf4a7d6c +
            Ic35d5ac4dac46d47b2796bbac6452161 +
            I27098cbe2d4fdd634385d771cc290c2b +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I7d60d53f883f8187700c4e78b4c22f1c <=
            Idfcf7f3240d92bfc87d44833bc00ff9d +
            I73d2731c1b1ae5ef73ce0eb9c8995912 +
            Ia0caf6693d441ac622f416a86b665166 +
            I5d7a0739e447775e00115799c52b11dd +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Id6fcf4b7af4a37c854a12e2ae80851fa <=
            Idd5b362dab4f93bba0c39af78c4c5981 +
            I2a4b3573ae7c3b38ec34591f20c1d076 +
            Ibb6e54edb9d277242c06d386a9a75a26 +
            Ie95793e09085b6de1383a37cc7fc41ac +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ifa5e5f7d753964f14f0f16dbe552fd85 <=
            I627e4bdc8061c69e3fcac17535b9f1e0 +
            I28ea268c5b51ac1d9249e96599bb6b0d +
            Ib97b2670a6cd88b2327f07f62d887900 +
            I134a734d93e62f6ac6635015fe3a2096 +
            Ib24b68cb35da39a743e1d90bba3f0836 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I900d471b087cf5a436c2ad66a84d8280 <=
            I5ca15c7da1f49580ddedd9ff8ba822c0 +
            I6aba8ca0e4b20a6355b43a70f19d9d8c +
            Ie9a316de516ec4fb828a614c67e38b2a +
            I745187336b8a5ae4eac66e90539752cf +
            Id4cdd72193e90dddd211af73d7f3634a +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I6d1434907f0292ea2ee47cbc5b52bfb9 <=
            I276c2ce5d3a1b7551c2790971071b094 +
            I77fd8001d879fc9e9117464fba27902d +
            I6d0d098e6d47dea04d6d7be67b648a0d +
            Ic3c59a5167cb83fd76ec6236572b1f3d +
            Iccab4c19a9190689f90a42160e2379de +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I938bef7ba7ae1739d8e6a6a7c117a1b1 <=
            Iff777b2c4a3939e330c4cbb36cbe1ac5 +
            Iedf37dac8b3a5331277ae4f0176968aa +
            I3f6fad8bb0fba790fcdb1612b6fa7712 +
            Idc549661d6694035874a3366704801c7 +
            I275ea08a3dc0600d8ccb6300eb7f2a6b +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I6384a9416b2d1da01df1b2d7b16c5390 <=
            I0a9cb91319cc0d0c1c4d0020cce321d7 +
            I9dff504e40aaddefedbb7b0f822c844a +
            Id9edc6ac95a260bf5af3de25f00e9e9c +
            If0676ef300628c4097565b13ef2d8854 +
            I1b53098a7240d2b5dc1f5c5c3b4bcc11 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I5097a79e7cf7a30d38ba198d1407119c <=
            I1cff7306aaf303bb3342ea3d72048908 +
            I2d839c10960739097d449efab58b9fd4 +
            I080832c25509f7003ed50d71210bc7f7 +
            Idb73eba1bd4ce25a6109e296f51e7dc4 +
            I278659ca1a0b093fc883d01987989dc0 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ib113c26c8dcf49c972c41a938059a787 <=
            Id033e7adfcfb0420cc592a1fb6c297b6 +
            Ia443284a35e0873de59b3ae55b7f809d +
            I2b807c16cfc6d65cb2a7f28ffa837974 +
            Ie467c5fde1d123da4e9587b5a56748a0 +
            If92e66cba66732798dd19f968a5ef8ce +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I970c4a25a8bce82a9d2846679029fcab <=
            I4ba05e74c2f63e2f4c59268775d549aa +
            I8289bfc08a5d8979ec26825bcb6e3d18 +
            I2b32537c9178028493af165398a60875 +
            I18d0dd7a10d6533f721a2392d4ad2d02 +
            I784c4e9fb75c314f271477e0621aaf7c +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ibe2af096ad2db26e54d8b4b3bb05175c <=
            I299b37fd45c6ee2031fb2c74caac73be +
            Ib8603cb82ceb97c2f35bf8209306a457 +
            I18916d0023ca275d84c52af07dcc5ca2 +
            Ic7d5fe6c4b1dcb97d10ba3de2f95d1df +
            I3d3aafdd4d9d3e9fdab1f487c48a0ea9 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ie48569c467fba0c1291f71d6080ebedc <=
            I26bdcc44692db066911c8d5b0a1aae0c +
            I8d26e73fafa909f1e26e329828cf4888 +
            I2c72d6c5fa6968dffa6517cf81219875 +
            I05aabdf73200996b7bea8db700fa8930 +
            Idb4c722992139f39914af7085378c6cc +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I90e7ded06617b49cdb8b5301fe9c6a20 <=
            Iaee91a5e94c3f174682f72a1ebfd0021 +
            Ibc1a16427d8dfa5ee20dac15327a53ea +
            Ic1120eb027841908cd64fe5c7274da14 +
            I4ee3f608cc8f8df27345949f1a3713a7 +
            I63c9deb7e6a4b400e0aff6887a09e647 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I4920014f5d017f4e840dc3b88526955f <=
            Iaed26e1c4a2578d16b111d15d31339d2 +
            Ifc52604a4f9f9de392a35f2f9fe885b8 +
            I4037f1b207aa101f354e59eddd7c9eb4 +
            Ic0a580f94f3d03f72e3a487f84bf6612 +
            Ie6f67c6e4c5e2b8357c0a902979e8722 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I03b70553f1c501609400574ae7cd73f5 <=
            Ibafedcf9f2990ed9c1efa973a0b1d81d +
            Icf4405d4a4063448a2be8ad0354ab1a8 +
            I778fbaea65beeb6de599490daf3b7e3c +
            I1d7a4f99e3975fd01bfe5a9a1da84765 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I63c9bf68b43ed66c51b0f4c0ed92e9ab <=
            Ie3c88bc240576aa220f0f110b13bfdd3 +
            Ibc8679379ddc43ee4bc508a1f577eb2c +
            Id66798f8ea67e74a67f264fe6b4503a3 +
            I059d847e09f5aa3f6a8147062f4b13bf +
            {MAX_SUM_WDTH_LONG{1'h0}};
          If408dfead07757878cc878131bc7d6a3 <=
            I4ed5da534afbfe9ecbc10ef4cc649a55 +
            Ie2e3d64640c339dc51512979dbd6a173 +
            I772e844c41387e7079259875e0ba3fa0 +
            I48e5256ade4d061a3b5ba08a53252bc3 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ia0857d63d309807789b6ff4f6028f1b3 <=
            Ice8765807beffd3acf59fa137ee0baac +
            I6e4786234b286b12c83e06e93c628534 +
            I3e8e280553edaa5c8555ace81ecc10e0 +
            I635fb29c55e0fb5cff0b6f443c2e3de5 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I53921b825c5e434b63bee0e1ecb7a517 <=
            Ic2f450f7ab60ba57dfc1406c92c0f077 +
            I529eaa7e5eeb6d0a1aba78df5d5a2fa0 +
            I839895c8614ff28df83314c44824900b +
            Iede5d56e52612e083407888da49470e5 +
            I088c5b971a2def57248769a33b7d2a2d +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I5e68f84e123c37f19a03c13892c77e19 <=
            Id144785da9b171f1e2d0e9182d693e31 +
            I439c7c302b535bfd7db655c3c607d71f +
            I2a0dc4ed573a544cb13544e049514903 +
            I39d9044227c161f0163e58dd82aadc90 +
            Ide22394fce1658f9e7002bdb30d03c2f +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Id5270b57c6fb4b18db3bbd0a523e467e <=
            I0cd8a6e719305ee3fbe8228081993957 +
            I583c6d23506c7d7b84403bfe977ec1ec +
            Ia422fbdf8f318ff3ddc049d1374e7939 +
            I8efad9622c05177563ab8a2747879044 +
            I9ff276a14d3205b98174a8a736f79774 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I3c18a84617eb21472d53e598700d7f4c <=
            Ic566fe27ccaf2220101cbc49fc187a6b +
            I618363a8ac413dd0ee52eb658940eaed +
            I1d648ed8f07f0743a6d616584270c513 +
            I03038b940be8bd21bd26b150b28754a6 +
            I123255637493b9c7924e3a72d1b86ee9 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Id36663e7a01fff3170833ecfecac1321 <=
            I2133d362ba45ceb3dceaa84e95ace1e6 +
            Ib43383830037df764b48c637a28ab6b5 +
            If2ce7b8d2573494564393f7d426fa47f +
            Ied4ddedaf801fbd7238d8a55c17c8090 +
            I87e6ef84894cfc86b94e19c9d3065bc6 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I8d3be15109c7007a79fecaac0d891626 <=
            I768afe193d9d79b136736abc6846d945 +
            I0aa93075086164fdbab3814d60633141 +
            I32c35da92922c5b477f8aba837fa6d92 +
            Ibf547f8a5e1059ffaabeb3f447904dcf +
            I4c32900878260a261bc5403e8abd6258 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I92169cc57291f20d336a479e392ec271 <=
            I54166b387c02e12374d6febc425bfb7a +
            If06a1563b9d7348de03a98d31bd85b06 +
            I3e466d40a4447a23953d96d2e6d61d47 +
            I3b2739319710681986b9d3f8cd04f619 +
            Ifc100357ae3f754fb0e3863334bcc764 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I6178b220b469b40dac39168057023a1c <=
            Icb2805685607d5fedd0300c9d800f863 +
            I28fa295ebd90c2b7255d48ca9ffcfcf3 +
            I4fd45670f88265e5d7aa6582f3ad3ff8 +
            I5f607bdc9b276fdf07a17a11a20a6720 +
            Iefe9e5376010997c0ee52eeb28e57a25 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I55342938216a0ea0889f96c2f6c05ce5 <=
            Ieca5b21b91e150c9d509964bdcea500d +
            Icaeb9a2ec8ec5822658fa85b88cca04b +
            I76e4c55148effeba62a4837cd19c5e51 +
            Ie6060acdcb16b6fa6aeeb649ed621053 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Idf28431c76a84a48dd895979d2b11a63 <=
            I6b7a8ba12de5b44817ec99faebe54617 +
            I58416287b268462d28f55c6c2705e613 +
            I2d636a246d815a4d12c478794860dd40 +
            I46c2b923860b0d1c01b9475f4467f280 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I1ef61124c8d62e8f6a82a729fb091694 <=
            I9b8cfdb69b76453a3ac687a1e098417f +
            Ib2963b82260024e1853d297798d88d3c +
            Id59cf860d9f4aff11b205b8970d93df3 +
            I38b4eceb159ecb0dda3920290a21a02a +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ib8bb96f0372323e6a8072ca56fb9396d <=
            Ibf9f6d7baed9e761b69fb41442761ac6 +
            Ie945349d77442536992d9ad52ce84218 +
            I3bc01b072987a0c980615abbc2251e5f +
            Ic45561ffe1837c3d5bb42c695a377f82 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I432f74dda4f6b1cebdf5ad59c659080b <=
            I67534b68fee8f76ac0c5e64cd02aba42 +
            Ic79072d9e42dbc9974231f1d642b3f12 +
            If08adda7d796da7c7849e472a73282a3 +
            I3db0adb3457cb22c755f5d29a8fe7ed8 +
            I3e76abc721bf7ed186f4d0f8f4bbf4e3 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Idc689442305acd00f0f32416d8fb3773 <=
            I277d7065150714e33d8ba64875d18190 +
            I9bb4d58b1fe80549451b00c4ed2b3885 +
            Ie335e68643fd2b0a53351f4bd45c3475 +
            I32679702c19eab37b46d13bb372967ea +
            I1afb4061458e9d2f5799afa1f2373bd2 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ida03738adc101c03c2229756bed2469d <=
            I0b6cdfa1dbfa774fc9a12d856e61cddb +
            I5160de2c5ce4782d8f8be10dc740694b +
            I3319313fe1d2b4ec2626711b187b4a5a +
            I85dd6a9634284c22027b4241551ea628 +
            I18bb9a781a4c314fe6bd990e4c275f67 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I4d14c75f28f3e516c259ea288996131b <=
            Idadf072247b351cf51d718f797c3b375 +
            If4d63635a5f99c4dc9e5b57712830c20 +
            I75aaeab4f372e28a8e51453540f9c6b2 +
            I51b1cd475d0e389326b182cbe680a402 +
            I49d7342f105c4502377abd23db973752 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I6e6cbbf430d57f347a0d70558af143d8 <=
            I6fcb3b133a6a654b69f41468a713d922 +
            I5eaa11e26f19b94dcb7eaee7f09d24b4 +
            I586aaa5c55efd37996b01febd3bc60a4 +
            Id5cedaa397ebfc2567efcc2f8a648db5 +
            Ieeb12d463444ca36af1ecf2e09504c06 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ib7487df45118e44acec6b9d07bbd5969 <=
            I8613cac4ccd4f956e8a0ae7b627f5be2 +
            I7d85b73e85379bf3a480e954c05516f3 +
            I2266afbacf1ba750ce18f296aba1181d +
            If12366160fdc899bd71cb0de5bcfd84d +
            I17525df1798fa2c1c4bbc4a1ddcdd0a5 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I492f382fea500462b3d0866240fb91b2 <=
            Ia5c77c9be26d62b026f24ee5a5e25fb8 +
            Ib5c8d91204a2d313c9c23110a53cd0cf +
            Ife3bb8945e14d8746c82b66886293997 +
            I887911fd9466f4d4fa7f50642d610d88 +
            I90c44c31fa7903a81826c1c568597362 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I3fb3ebddaf28efb56092d19a1b4695de <=
            Ic4af6c9097257c9b22a57ce4b79b40fe +
            Ieb7b388ff89e352dd239e0ccbe7b9ecc +
            I89f75107ea95f207b9e664a1f4f0746a +
            I6a86b03402bd2e35208d3fc74601f9cf +
            I3997cf122743b612f49cd5dd125a9201 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I22a26b7f0b1c8c16b00597732ce2ab23 <=
            I4a403449a9ba75243369032e1cca1a0d +
            I886750aaf8d2040c3f12ff113294f658 +
            I0e52c25aa840402d944cbd81f73c1ffe +
            I1112c4267582ddb8148ee40d9529beee +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I2ac08a2d8c917ecb37fbaf5325cb0473 <=
            Ic2159627df2efa5e677fa6f4498bdd31 +
            I58a7c7b05b84d292cd06d68e96ecb9f8 +
            I20c4e393929b875521e5316f4d8e2d42 +
            I21c207af859b94634d3750482b42a2ca +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I50ff8f51e75fb9ce3db983c2a0f57196 <=
            Id5b4ee69444e5b499476c05a7f1d6e60 +
            Ia308e09137af1cb50167562efb5da628 +
            I2418ae211f327ed45cc70c42078180dc +
            I2ff2421bd86bf9ec110724460f1171e9 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I444bc340ffb7ef7b72d4d2e761d58872 <=
            I48b39ee498563e23c3a4be079b6100d8 +
            Iddf65ccb4396288264a400ba37cbb655 +
            If29fcea810adbdb1c4d8a4ace1d8081b +
            I6ba5c453b17e4b33c61caf5d70041c4a +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I039c6cac5830759529595a958b7f65c9 <=
            Iac8cb32c2d86b975f51a2ed605002e51 +
            I88a325547ccfe4eabf90792abd60e356 +
            I0722ec4e9d400f8eaeacd060e42de79c +
            I08318099725fbe033ab8d5427eb8b278 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I0584de7d919236ab138e288a27d08ff1 <=
            If85d9a95c1c02ce2da1dc3486b53eb81 +
            Iae21bdea20a6266d3f69aa680b6b2817 +
            Ic6a7a82d16e6106071934ba79d3698cd +
            If36cb462cdf20b0b1758cd6417e524fa +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I086402c82ec67ae09a9e6360c58904b4 <=
            I59fba74472ded0a985cb237104ac127f +
            I77e1f5f504a794edbb89c66cf1ffcf66 +
            I3cc30aaba3dcd3eda262a19e85e53117 +
            I40e8463645b1122b7cb224770fa00447 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I1cefdc831c146187c77f861b3e2d1af0 <=
            Id6105518ade80c89d4f20222a2382efb +
            I8493e2dac01f009db1d2d5504b49d135 +
            I106d0e71b7378d110b0a624e5cbf0d6e +
            Ide386e751e06dd5df0c042cd76f0f800 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ida9c16ae57d17b6faee8a54838860447 <=
            I185085cbf8da6df921ba32442b28bcca +
            Iaf3a0b5ea5d9eda47fcced9260922bc6 +
            Ic8f0049e1298b14b4e039075dc0d5f74 +
            If63bb4681bf1116c0d1db3aa21bf52ac +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ia3b9fb112f39dd0ccbf7555659369efb <=
            I5c278aad08b7c4b0237d68f88fcb3f3a +
            I9222c4c0eb2b110fd80547d46ba17036 +
            I95ccc219b5f5038641b38dff6db0b222 +
            I566c72342c69969892480fae41232c37 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ib1bfcdc0c972aafc99116ed8c0511445 <=
            I21842d06e25948ef461d1fd03485f86c +
            Ib2c1636a66f6479d6123a038cbc668d5 +
            I69c2b063e61e14f5d49b907095ece00f +
            Ia0f7deea6b1ce1050dcf97fa99de9178 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I7adff505c50450a04f1717cac1adebe7 <=
            I37e360420c7dd061de93a6647513676d +
            I535b29f7177b4fc009ee998f1f4f7d7f +
            I45ef0ac486fe043f57e8a46aa91461a3 +
            I992b9876530d53c1b62d98511bf41942 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I699feb4382974a02b21cb387c13f7f3f <=
            I8e470b68bf35c647af42b6e46201e570 +
            I8cbafa797ef136d7e50c909dc160deb1 +
            I850c257a0412bd9bd6001817bd9d0ee1 +
            Ib8861f627f6273c0a031bf43e7812a5d +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Idc99c3b23e49aca3c98f0685ea34441c <=
            Ia526539cc0f844b802d412b7a17cb6a6 +
            I71bc7271cc432bb3c5d0b7a416cdfc60 +
            I12e8b8cf609c2fbdc72efce9bb5dabee +
            Ieb5bac4ef0f5e4e0b826cdc43ae71471 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ib67318fa6954ec8f3247927d34e74f8c <=
            I26cf25e680483bf4e556d74efec35ee7 +
            I9cbe73d708c561d43d05945552d32dde +
            Ieb9720b6beb2363d651346ef0233cd49 +
            I3cd0883d9f0ba7475f474f1e318ef023 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I8774ce3f11362915c4331d1026e452dd <=
            Ic989dc794ce4356856b3916ab1889589 +
            I82a225237aeb1ceb31e8cd18b1e45c6f +
            I2ea27544ba4cc14d0f7ccf7158a27a2f +
            I5f8a41ab83a9257e534973e981e28e9b +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I2392b2d17ffed6073875fbe8e92534cf <=
            Ibcb80df5bed66f8498561e3f3ffa4ec4 +
            Ib7fde6a2ec1ff0a3af10bccf3012e63f +
            I0e420136675d5f0d1aa027d589ee8741 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I3a4f0d3e32596ef05477f494768d4266 <=
            Iba75ff0f3b67c7e28cf627706733d528 +
            I4854ff71aa885da3d07acaaa24740d7c +
            I4aab6ff52e3fba90bb7417cb50766125 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Icd08ff59cf6be3ba97698dd55703339e <=
            Id65f22fa8fc9c47bfd00c796b63c9fa4 +
            If7543e2f5a158b1f3f3a4078ec54cab5 +
            I1ba7f209cb735471073e8051026a148c +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I985fb7ed22a8476ea322c9e3c2b3851c <=
            Ia81c31ea4f4786136b539c9766987596 +
            I6a3824a6598bbaa138e1e763ad85f5f7 +
            I711c5cf9fd8c5161bac36060b3443503 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ib985709316b1b0a9d3fa3c1eaf6c641f <=
            Ie380b37a78242e6d45b659d568887457 +
            I72108531a608f6d5e51a481c68d7b271 +
            Ic9740baafb1c92e3a25f0a1e7bc46486 +
            Ie3591b22e0e127f04658da68d4846be9 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I4be898887dff6e2cebe53f135ece131b <=
            I484ec87270fcc959a486ebce40a9a03c +
            Ibdd9957b7f1a319b797c021933ff75d7 +
            Ib1461f456ebc14f449eee77e386a4c69 +
            I409129c0bf5d361e9916b6dc98e69a7d +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I004db04f61fb57aba81e15cc015442b3 <=
            I5d80b7c7d102d2c2bfa73a68c73376be +
            Ib2c327648cce481482eaf0467e9227d4 +
            Iaf1d3be13e6441a7a9ab3f286a7dc21b +
            Ie4f4faa470f572da2081b63b6df6e392 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I8f7e3dfb2f728d4cd1e79b82b62b0406 <=
            I8636f5c91b567780d3324e4b8a320fc2 +
            Idcc745602c4b7b34df9c3d68f9a9d76d +
            Id5c9a9b9c34c8f9d56df0aa8d780c9d3 +
            I5011dfbbb0eccfebcff255e4a2c5e64c +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I991054370345e61638ddaf81785505bd <=
            I2cf5304a672431888916e08b3c15f0c7 +
            I989091b3586964ab598f166a89279d16 +
            I5f7b6e6a30348ae86057f7e56f625846 +
            Ie32ca6b91d1c55883be8f63acca78764 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ifa1f503965270d10e7a5c9a15576069b <=
            I9164fa2a9a33da6612ea692cf3fa7d2f +
            Ie8befb003fe83e774e8d1d01d4e2f4ad +
            I1f1f2fefd3381ee48ab0ec9c9301754b +
            I6c7965d39dc839a9df56e628c77a5457 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I24f773842a4742fb58d09cae45717b2f <=
            I288ff69a7395e74f7de8da5a6a7f9062 +
            I98a2aa729628adde0b6047869bd12743 +
            I1140fa91b5e22ba0c094c03295781e5a +
            Ieac9cea5f36bd82f87105b530e8fb614 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I5bac7e0d778a547a0ae764fe259b6f7a <=
            I5a4f0749acdc34fd0786e4b3d062f88b +
            I283107989a436e2c720123b8d9e335c2 +
            Ic488e78b5c73251b673301e84c4b5b0b +
            I79657595561eac53237215fb4110f09d +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I255577ebee6768871df0224fc1db2db3 <=
            I079932780612fbce79cbe9b58bb6c2b5 +
            I61f5ebea2bbe443b644c95ee559c2234 +
            I9b46463a6c54c3668e76190d942b7b38 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ia7fb4af3d3529a32f902a52cf5598474 <=
            Ia92defa0ca87c7c30fbe901da40a575e +
            I21255a0ad20a9668c958faf68d53b2bc +
            I3ff883ad434cd5153b67186b6b21418d +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I2c98806141f064c9e92935b23a84ede1 <=
            I914bef0326cf82d350344317eb1359be +
            I6f69796a6fe6da57066319ec8210c1a3 +
            I92abaae6fb89206885616877cca1e25a +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I5680847bc8d224fa4ed93b2fc0d841e1 <=
            Ie43a7f8082f91c2955076a6373028b55 +
            I8786eb767f02164cdc32f14f41b5d0e1 +
            I33668b0ef7defef974b7a4c0f87689c0 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I365254279ebb10dd7ba0b3482d5e34cd <=
            Ibfb57f2b507c27759a3556759f23977b +
            I064499f0315fbeec7b6cb50583388a07 +
            Ica0a119af1728ae253c16cc3eb93f802 +
            Ib7875bf9d30d071e62a474c50d88ba06 +
            I338daeacf82ad288b14c6b5bd4099870 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I57bf4ad773cc058ae1bb7b1911dc3174 <=
            I7b12345fe53174cadef6811fb8869b42 +
            I6521c9167261db6eb37f50b66159ddb7 +
            I44e5ce0cdf812c5b73e6e638da36e414 +
            I6fdccefd034e8b4b86cfa997502512ae +
            Ibe085a39ecb07a8dca62002afa38df93 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I57072dfb29c4a3d2e2b40e46e62f0d95 <=
            I9785922874bba479ce4a9bf1759e2933 +
            I0e3286fca6cd040758950259ab663df7 +
            I9ae284c0089ae462a1bb9d168bde2fd0 +
            I202aa0814e7e28a6bd21db116b652b4d +
            I1f88dddf05f255942e2749891a7733da +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Id8cafb6f76321bdaba9711133be7be99 <=
            Ie7e196fbb66ba6bee51ef0064ca519c2 +
            Id7619819e1297844d92c8bf3a1d61926 +
            If8a259e0c4f1839e852abec6e1b904ee +
            Ib2f34922b0d5346500de093275bebc94 +
            If1d0be4e9b995ec98c346e8392b9518a +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I6344e71ca2b0fd39d36caedd889c3085 <=
            Ibb157b97546cb19fa7c1c0a7c79b1d38 +
            I3fdec80112b3fc543b217d1c253406da +
            I56a4443759b3d786bc9a34a0dc32abf0 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I0c99a68e0bed90afce18807acf7d55bb <=
            I8fb1602dcdcd2912ea8aec42e2b7848f +
            I5aa85d9503b0e4ff46bbd63e873053ca +
            Ic826d371f2cfc503f5d9e43dc17481e1 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I1c95650979c86310ae2a949961c9db11 <=
            I7de222bc26e38b8b6543819701740302 +
            Ia7673d73f0535906a99d6cb467892104 +
            I5502f383dff392ef1be4cbbf9dbc3c2f +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I04eaefa5d133e53494fc270b07be7043 <=
            Iea765ae5e9c65b3186445b15c56f69e5 +
            I103ec7cf279f527fc6e3648a19a12a8a +
            I96e6f1dc0cd451da6ac9170d5f83976d +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I4a64fa2412eb8058c2dfd9351d7b297d <=
            Icf266f710358631b7119ef526acb301c +
            Ib20dec1346f227042c749ec1abfa4d39 +
            Id6fa8ec5d1062fc3e09bdac65ff79f45 +
            I10cd840a369d3e25556a41beede2be27 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ie8bb2fcb752c6a33254963d1ebb4130d <=
            I0f3c4fb63ef1e88168b4d28175a0b68c +
            Iac6fcccf3a0cfe04edc0d998b60c2681 +
            I1fbcaf2f6be01b129ebc24dee8a65396 +
            Id85c2285fcc45211f0fa6963b74a663a +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Iac05b7e3ae18f948b72c356ccfb8000f <=
            I2ba94ef71f97b9ba731b306d4a5fd02c +
            Ifbaae8b3da03911a4c96d4efdb9283c5 +
            Ifba1584d599da13b98a3b76b4db10974 +
            Ie0bdfac78159144aa65090028931a3bf +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I27da3f75cca6c49e55db90306aa68e94 <=
            I5529d6db17b6184c45cc4487e5a2c24a +
            I685699f60c76b00df87c9c53e9a8e448 +
            Idb862697f62a6c678072de760e176096 +
            I28fa30cd1f3b476fa6a354863108cbcf +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Idc7fed723190098341225fe01ba65ced <=
            Ie3361a270ebc41698ef4651bb3548a49 +
            Id0842da8068ee88d99af7acea50e7b77 +
            I7a927f4f266cc5253ec30f5c127bb17a +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ife9065805598960919ee4f14c3cc6fd4 <=
            I74b55d2f94073ba8f948e4b02386867c +
            I03a8a458ee0942c35001cbfe8e589222 +
            I7571c7c306861230de71a75fca79c5dc +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I717c5c2d6a2be61593492ae5f17a112f <=
            I45cb51c25c426c296f97a5d23a08c063 +
            Ic1af7410a9d11c5324f3ee5b2e0e9dac +
            Ic79811a48840357d0b6303e7b19413dc +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I4c31fa8e6eb648439cdae1de1afe0d6f <=
            I0cedca0e2c589104d6f3318505910594 +
            Ica02d19b129c8b1d491ea4747a55113e +
            I0f29300446f020dd23cf847d3e3d3530 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Iead549a9af27f1fced7d9c36e7b5c3f5 <=
            I77a54091bc2c3d9006ecb3471b94d8c8 +
            I1c0df8c2c64b688ae417a238263f33db +
            I696db0b98e27dcc4657dc7feb23a881b +
            I9de41d0b279b84366640880dbd18c502 +
            I802bd5b13c183c37e842f7e9278f35a9 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I10422eb79364e7d0e21e1643d9060331 <=
            Ib6c0e635e659f54724737f0cffd1b0fc +
            Iad0f4602ec545dc6ef12aa34add00ed3 +
            Idfa432a87877e1ce103e56891745b62a +
            Iba52b84e6e215842e0ca8e72c42ebce7 +
            I0297905b35f06697625420b7fc2434f7 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I914cb87eba8baa40cd515334e59f26b2 <=
            Ifba318d4faf308168c5eac8fe92395b4 +
            I06e05a1ed002175a75d02b8b76f52c50 +
            I894ef04bfa1b7b39ef51b7c82f7686eb +
            Id2989aaee3930698cd374e6c9feedf82 +
            I8487a819dcb61016798cde56f9662fcf +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I32ed679af4ab759901aee43c9d93eb67 <=
            Ic9678deca4bf44a7b99f853334f6a05c +
            I83b77ad1a40dc102f28153f692516eb4 +
            I920f95bb52cdc9b07f93afc3a6b5c009 +
            I8d07beccef519ab4ce4024d911ac2346 +
            Ia2904a5d5db43a209bd4b358ace68c6a +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Id376dfa5141402f4d41a8858180ed87e <=
            Ia209e5b03deaf4fcb8ae12b731a49e0a +
            Id2e223005a932987b6f60663773187f8 +
            Ia8b29ca047a643f47bd3a0ffb50bf8cb +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I98a384bc62ee03f5ad7df20ef2d9af95 <=
            I99d236d41be79090ca7ba1fb6faaec4c +
            Ia92b76ee5b7d82a992a1b58147c0c0be +
            Ic45d0537b94bc30713c0a0ee07b1ec40 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Icfed259ca2bb2732d8e0c26ef67cd4cf <=
            I26ae9e570a101c6f8237d7941285b924 +
            Idcd5283cf7b42d403ee0e4404b5b311b +
            I337231f0dc7eb85f7d950262e0adb724 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I20861535c450d6e6bf11c45dac120454 <=
            Iabe5aea929c668c9b9728d073ffb00c8 +
            Id201f81bbd80a70006a10866b8efeeff +
            I530cf1f747d1df44b913f49eee90c079 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I013929385ad819ddfcfcc59c22902ee3 <=
            I1240c9410b897a4d0504affca5ba139e +
            I4f169c2c8c0768f2725ed655a03acfc2 +
            I342a563de39175fe4a6eb7e3e1ccac9a +
            Ief52461e4a5ddb128be5e439edf34862 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I34fffcb07fe82f11fe142f7c37f39155 <=
            I015630502f5cb4eb27b2a673e810f1dc +
            I8bb46c3eb9f54c5d1b28dc6aa0154358 +
            I938dd59e4cdf3434086f60d000113430 +
            I46d86bfa6de26f3cfef9d802549ef2ad +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I61ca60fde05ed88cce714dcd8c13b827 <=
            Iff1d4b06901796098f91e87a3c30f7a5 +
            I1e110e27162231650875dd1152d96e64 +
            Ie7274a7ffa053ced4f12a67986d3c81b +
            If6a3bd6f002d91e0773c4ab9caaaa01e +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I4907dd45c158dc7e0041c64f1fb388f6 <=
            I54c260db5c1b2c76527c8fc1cee229fe +
            I55e54359961ef6e5a63f1c2eb0ad4aa1 +
            I4f38c3d620b72f21cf6d54c7df4ba816 +
            Ib33e1c6d57e5e6fc465dc9c9a7cf29fa +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I2c8f6a9b9f655b317bb0af4d60fdbc4b <=
            I3a8bcfdab631a268d21c87b98e9d1c49 +
            Iad0ecc5208263d239e4a62c5563f52ab +
            Ic0b2f9717b8aacb34325fd5aaf03a366 +
            Id92a319da408be46970faf524513fdd8 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ic7dff631559304ec59f0696c66436d62 <=
            I95b923444062b4a98918c685c65996d0 +
            I06c0921675f464807a63c7965796f0d0 +
            I59adad4fd84c1fc233dc58f70a12779d +
            Iae182ffae6cea89363f0ccc8b5679561 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I6a239d3e55b4a9a3be9989a85bbec545 <=
            Ie40c90fdb38b3e4046ba89295ed77d7c +
            I13b9e098622d90a1074f636d8f351aca +
            I1972375d51767f0cffa5395a354b3493 +
            Idfe6aecb694385ce8c3c1544a4992a20 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I630f905e55f08e7d1569a08e937ad216 <=
            I9859b94cda465ceaaa5674eb19e94824 +
            I8d6927b0bcbbb318cf52987c121a07b5 +
            Ide40b1bf9c0b642c49a5685a62af1c93 +
            Idfbc5726963cfa31bb4324143ffd08c7 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I8d13eb3669785c4279c685763d4f3fad <=
            I5085f161323433d8d38be2e4511b0c46 +
            Ib66b897398ea0702b74bdd03774f3ae4 +
            Ic227f42a20219c6638ee3343ca445acf +
            I205d5fdeae55fae7be2f06f11c949244 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I25a6f3de9a9a01cbbdd32ed848561aa4 <=
            I16db9cab1981451a02dab21e2ca221b4 +
            Idc758f8e6fabb6b31b0a7d9c0c590310 +
            I3188d354c2ba494ffe210dcd89c00620 +
            Ie667e1755ae1561a2eefae9b63845dec +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Iba3dd4b2c2c85c4cfe770d9b52ef4634 <=
            I3d700e050cb7f22b0e381f3c72a20124 +
            Idc198bd5732ca5760d1a700a25273ce3 +
            I2253b32e46200a23dba243819fce02f0 +
            If7348fdbe0400aab92e8fd6a7cf6c267 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ie1b744387b5200a504e4874e14d2f282 <=
            If17b4f86674bc5fb212a1f7751fb043a +
            Ife7985db888089ea618413810611bfca +
            Ia020344403aad35e050765a4b0cc42b7 +
            I143b91852fddcdcc30bf1041332c4ed7 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Icf76cb69aedf4db01cd3444f4c4ba471 <=
            I4fb3fe065daa2708e55c812e57c19fb6 +
            I96f65790e2cacf7b529ce5b88598da00 +
            If077c67a062095cfe69f2260cee82833 +
            Iee5e74945ba15220f0f707c9c1927ba1 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I4857b5b50556c8e7fff4b2d3e08e4b28 <=
            Iffb7fe9c74dfc01a43e99a099c4e7e04 +
            Ic09b4671e867144fe9f54a09e74c5519 +
            Ic0ae1191869e636f9e4391efe93309ae +
            I4d1c47569b0bc8c651c897ac8e88bd1f +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I0a1e9cf99f1d4725327615f50fcc3ad0 <=
            I487b9b236d118786e475ccc5e4e56a6d +
            Ic46357bb77f6183329946f7e28294365 +
            I382153cec6f7d6258574e7c532186473 +
            Ib9d6c5be487a434fbafcda25ca9351dc +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ie844f4c446983ce381b0bc4c0e8ef7d7 <=
            Icb92c7c10f0bfc5d287228f98d8a235c +
            I90001da8c360ccff128f637cd672ad42 +
            I5001118df37d08bd19d322aca8ff3996 +
            Ib0d033ba28e8c606ed92207049c76884 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I6067f47cccceea96ac46ff0d457b25f2 <=
            I72756ea6a4997bc4afd4bfde1dfb2d26 +
            Iea4a7766d3b9d5d030ade1739859ef0d +
            I78e1205de9119fac3ae8f43c72ac71f4 +
            I300d9f403e33d860ff5dde9f91bae11b +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ifd6fd1f3cbf8884ca7f64bc42278e4fa <=
            I63c0c8bef1dea4e499a16ce01e781951 +
            I5a7746e9fbb8c009f83ae57423296cdf +
            Ie0ce2826fd13b0e0b23c91e97787691f +
            Iebfe0fa45e4b34e142e82ddaa15243cf +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Iaec9fd9e79371676bfa8ff14b4feae52 <=
            I275f6334127640b2de3f0f87f54fd74c +
            I3faeba79f7af7a006ab5cd256352e2db +
            I0c0be3347a7df9cc39997208b013f17b +
            Ieb778442bc855e93e11c9b13f1a7ae06 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I500757c4eda5d3d899aee47b87da585b <=
            Ie9fd8f7dc0c3849c0437a2a3d8607b4c +
            I45a6ef43e6e42594444adcbda26700ab +
            If36016df78d833c80e1355151c038225 +
            I57a393cc9cc9e1abc7962aa2cc840a7c +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I47bf091b0fa74ad511a760bad9d2506c <=
            I002869e450d79649d27441ce00bfb575 +
            Id11fd3a31b70da0e64138e71840cfb83 +
            I0ffb8b65525af38861280645ac310e3d +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ia4c3d0cd9957f678880de5775de76e0d <=
            I8e01532a1ab9534b8de0474549d41a2e +
            I507e9bd0265d9ca6cd21a46fa21ba084 +
            I30fb41a57460a0b1f21065b4b97ddd42 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          If5f957fa2f055b1c2c28e8d7cfe3e9ad <=
            Ifb19d75cfa0051107b5fba57bfc002b5 +
            I09faa07bf38acd96c4e29afd8a5167e8 +
            Ie8298c5c8ff538a3e37af46798f6d753 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I3608378a5da8c66bef58528d56192530 <=
            I79280400a4c9bed015106e5d006de757 +
            I1b01cadaac7d3d15007f0afe5c0ab0f2 +
            Ie7dc322fee8ca0b6b9659e5183e0d6d6 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ie6dead855e00ea0a8e6a9b7503aaebb8 <=
            I6cb09ac924c3b3b44443263e08c3315c +
            I8741c5cc763512d16cb1186fa3323f45 +
            I22c15857572603cc24d8a87cb47c33b0 +
            I91bbec0523f77fc52a88ebcc49267e9c +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I3bae5e6862e003a8b9a476f72cc6858b <=
            Iba4972a3b71a3101ab23190ed905dc17 +
            Ib38a46dc131d635b81fb7c196110fc4b +
            Ibc03a9b6115d0941ce9233df7ef2fa57 +
            I38ae79956762380fadc94f8126dc1c90 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I4431adecba8be9e5f21bc6b3e1f8cb10 <=
            I4bd98e902e805426fdd4606fcb5a5214 +
            I6b5720d71a0b4cd10ea34affa6631a25 +
            Id92d779518ae724b5fef5221372f8f26 +
            Id55a1ab9d158ea509e5f57286a3d1b67 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I21c7a2885126d532d00484376588a469 <=
            I43f52bcba1bd2e8ee5fac03320e4f19f +
            I391a2f354262558ff17d7d80b8c39e8c +
            I351dc309e916f282cc1e19303eee4112 +
            Ice615e7e18356ae4c3f615dd997be943 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I2c4d7339ff2fe68d060dd8d961dcab8c <=
            I9306d9ef7934ffe5902306b9783c351e +
            I70dc03a46e1ac0da826388abd3bdc503 +
            I72b4ef48363856af7faacc85eafbaf2f +
            I57b40c72004f2c3072cbdefbeef72b7c +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Iee518b15b067eec58cccfa37f7432ea5 <=
            I2882ae2eb6d79a5b96d1ed937dcfd8bf +
            I0dbf900b4f430b4c1106aa86b640bb37 +
            I9dfdffbfdb83572cc3205f674e5db753 +
            Ie38351e19bdc4f2ce9caf75fc3937dd4 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I42145be9c2a80288ba4a2edd91f661a3 <=
            Ia8abcb8cf8d9ecc17c27ff015aa0b71f +
            I5bbbc4eedb7c61516769f429a8498ea7 +
            If49068db99aa9d09302eda27ab51fcb7 +
            Ibba6269b560db9d4913e1e515ed8270d +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I9dc297ad41fafcda77f5347f331cfc25 <=
            Iec844d10736440b96f9d6c651e604efd +
            I7dbd1aeba00bb8b257990b7bb294211f +
            I0b3a936c3f7e0391111e696b2445803b +
            Ie392719059587a201c0148138ba2a2d4 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I846700c79f30ca954cc2933fc94d355b <=
            I02e672436ade3ee620c72c0d9ceee664 +
            Ie4d20df6b1e7a42f0df9a3cc26b12ac1 +
            Ie04e44d8e0756cdf34cf9ad53da76e47 +
            I4852d6bacfd82fef6fab4502d61e9a37 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I8af96a91457316e49e3f7dd5e57c82da <=
            I508cea40d87bec2672f980d145c89b55 +
            I80af3dcb716f3474a7257700aef89b81 +
            I6d4867d03d9187e95e27e99f7aecddec +
            I9200526d94c38e638370e9a2d7fed75c +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I7d1c247500d7d32e406b2a5f7e2b745b <=
            I844b9a89ffb7a5e48979fdea546e244a +
            I9d05dc0e39e85c23b62f343a8de12e64 +
            Ie96877deef8b1676138f814c4a720800 +
            I15b8aa7d973edcf3b2365040f5570d82 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I66d85c030a8864505298919046056305 <=
            Ibddcc2e26fba20dfe2a2d399be2bc45b +
            Ic6e3847f035738243f4c5f71f296da57 +
            Ie9c5e7c98281cd1deb6acc51590c9d9a +
            Ic3f8e77259ee3eb5be80e11b607818bd +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I4841257ae596d9d3e4eb1e6f886956b0 <=
            Ia5e26c2417aba1005971749f4ab2f367 +
            If6b40a030cb120fe017bf9d39e1a35d1 +
            Ifdcd91f925b63e0817798aa6e9200e50 +
            Iabf228f57ac154c417389f6711af1950 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Icd6f7ec117f9ab4eda8c5eba41386ffa <=
            I9fdfe73e77c384d33196c0f2d2a2fde2 +
            I30b5c7aadb5312ce96e833704bb3a320 +
            Ia18bdb8d2f02b50281f0acd4a45ac973 +
            If37de611ce4fa330c4fc9dcb87d4d95c +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ibc0498839d1d9b6dc853b8e5d7a88fa3 <=
            Id924dafd31fd0af0b28c7e6b7e95ec37 +
            I926c049036f53f0a0a6ad369de116c57 +
            Id0762ac7710c93249bc11c6ce4ae51a0 +
            If3c44eb85217da3b6bddb5aed97a9bb7 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I142ebca7f155e287e38ddf45423ab0fd <=
            I33703f538ec70268e6c00ad6eef6c4e0 +
            Ifc7eec6765af08463751db128f8818b3 +
            I9de5e90485b3f22e9003dc8a7b22a79b +
            I8c36318c45dabe6bf540381373f09fe5 +
            {MAX_SUM_WDTH_LONG{1'h0}};
       end
   end







always_comb begin

            I97afe24956b7f87cd431f048202bab67 = I5033323484d90d6bfbe03749019fc6dd + ~I1a632a3e06ad738d5865acc77e204f48 + 1;
            Ic188ebb37ff178022c61400613f4f3dc = I2bcab411f9bec1541259751bcb9e0823(I97afe24956b7f87cd431f048202bab67);
            Ifeb14203f4daf31c7701a6a742be57cc    = Ic188ebb37ff178022c61400613f4f3dc;

            I117235e3ac8e68e4c1ab34db1612aba0 = I5033323484d90d6bfbe03749019fc6dd + ~I71b93abe4b20e6a17ff17e0f33ac2ca5 + 1;
            I3f80921fd94cff373648fa34fcadd4d2 = I2bcab411f9bec1541259751bcb9e0823(I117235e3ac8e68e4c1ab34db1612aba0);
            Ib581c19864deecf01268595049268b19    = I3f80921fd94cff373648fa34fcadd4d2;

            Ifd700cc9d18f99b63f1947f3ae631976 = I5033323484d90d6bfbe03749019fc6dd + ~I9184110e3e9b8614460fc0abe5fff2d9 + 1;
            I229f7430f590d86a323b48806beec48c = I2bcab411f9bec1541259751bcb9e0823(Ifd700cc9d18f99b63f1947f3ae631976);
            I661d84af541e30828bcbd962d72baba3    = I229f7430f590d86a323b48806beec48c;

            Ifffbe3d1007fb07a20d3b37902b3ec95 = I5033323484d90d6bfbe03749019fc6dd + ~I535cad8c919a4330257eb5b4bed61b3a + 1;
            I26fa0a5f87600d9535e8f83fa1a11136 = I2bcab411f9bec1541259751bcb9e0823(Ifffbe3d1007fb07a20d3b37902b3ec95);
            I1c6928cccb4bf7ea7dfd74e425b9624d    = I26fa0a5f87600d9535e8f83fa1a11136;

            If5443777169422ea6e1e3f709b970e05 = I5033323484d90d6bfbe03749019fc6dd + ~I7ea8fe50c45e213f3257060e2813240b + 1;
            Id87360986474c9bfa5266a90b59a9a8b = I2bcab411f9bec1541259751bcb9e0823(If5443777169422ea6e1e3f709b970e05);
            I6eabc5c074fb1e2183a5f1ecee87a518    = Id87360986474c9bfa5266a90b59a9a8b;

            Ifaf9fc93e4609d818aa46751754c17f1 = I5033323484d90d6bfbe03749019fc6dd + ~Ifec9abca21cf476b70e0befa3926b46a + 1;
            Id63daaeb52208682533b5f136480a29c = I2bcab411f9bec1541259751bcb9e0823(Ifaf9fc93e4609d818aa46751754c17f1);
            I0107769bbd7c239685b4818731334437    = Id63daaeb52208682533b5f136480a29c;

            I419caf964986c655df84d043badc37c9 = I5033323484d90d6bfbe03749019fc6dd + ~I7c191c2c2be09886d0f31e4368797afd + 1;
            I1e9d5c2338b6f89e43c30c0ad71f675c = I2bcab411f9bec1541259751bcb9e0823(I419caf964986c655df84d043badc37c9);
            If723180430080198d18a08d6775ab208    = I1e9d5c2338b6f89e43c30c0ad71f675c;

            I3095214ac0e6c1323e75ee4ec85e6821 = I5033323484d90d6bfbe03749019fc6dd + ~Idd01d014f0469f893305057ae3f4cb2e + 1;
            I11cce7dd119eb0e3acafc12dbc6d3536 = I2bcab411f9bec1541259751bcb9e0823(I3095214ac0e6c1323e75ee4ec85e6821);
            I44abc734d6acf92a8e8209186d7a1676    = I11cce7dd119eb0e3acafc12dbc6d3536;

            Ided9739bf63937933250a6d0c37535f9 = If5dad13ac41b3034bdb034bc86c9b348 + ~I3f59174b3764a0b0741462024be9fb92 + 1;
            I934b111c08439d3797cb8928c7238f23 = I2bcab411f9bec1541259751bcb9e0823(Ided9739bf63937933250a6d0c37535f9);
            I72aa55988d58c664f3291b5786fc8ceb    = I934b111c08439d3797cb8928c7238f23;

            Id0f139b9f3848b45554ac8429230eea2 = If5dad13ac41b3034bdb034bc86c9b348 + ~I0e112f1d4e9c934a118f79f3856744a9 + 1;
            I508cb12fa71441b216fd7c1899d00e24 = I2bcab411f9bec1541259751bcb9e0823(Id0f139b9f3848b45554ac8429230eea2);
            Ie69528583db8155917ab3d32a446de04    = I508cb12fa71441b216fd7c1899d00e24;

            Id9feed58cf9565255abfd0bf7e3ec068 = If5dad13ac41b3034bdb034bc86c9b348 + ~I65708fb59e90bb79b8107da619fe63eb + 1;
            Ic69c6ea6b4f360efae87611c00b00fdb = I2bcab411f9bec1541259751bcb9e0823(Id9feed58cf9565255abfd0bf7e3ec068);
            Ib22b47d95b72871e74069fe80a191680    = Ic69c6ea6b4f360efae87611c00b00fdb;

            I30a3be3b5f6ad1880a917eb35659a1bf = If5dad13ac41b3034bdb034bc86c9b348 + ~I0fc42ce9cc31d781ea3013318c25a571 + 1;
            Ifccbe59b7ebe3f692f5b7e7564ca50ba = I2bcab411f9bec1541259751bcb9e0823(I30a3be3b5f6ad1880a917eb35659a1bf);
            Id9451e945bd26b8dcb4cb83ab4ade73b    = Ifccbe59b7ebe3f692f5b7e7564ca50ba;

            Ie8148d9aa962a733eb65877b902a187d = If5dad13ac41b3034bdb034bc86c9b348 + ~I8bc3210e86a523accdbeefe7e72ee4fc + 1;
            Ifd7275bc534fe9da81b12b25ed218e91 = I2bcab411f9bec1541259751bcb9e0823(Ie8148d9aa962a733eb65877b902a187d);
            Iba4627d3d3ef91f168068ed128c04113    = Ifd7275bc534fe9da81b12b25ed218e91;

            I69e98cf3e679183aef6005bb582b18dc = If5dad13ac41b3034bdb034bc86c9b348 + ~I597c3f5c14e235f90dc8c796bc3e931d + 1;
            I01a99ac2a3f919f4fc1680edb11c576b = I2bcab411f9bec1541259751bcb9e0823(I69e98cf3e679183aef6005bb582b18dc);
            I39bef4d462b0a3f88ce1485a58d66da0    = I01a99ac2a3f919f4fc1680edb11c576b;

            I7f42a504fc61c9548acebdd8b1858eaa = If5dad13ac41b3034bdb034bc86c9b348 + ~I07d68462362d8453e83570cc793c55db + 1;
            I322b3879383d75c43c55535f01fdfdd6 = I2bcab411f9bec1541259751bcb9e0823(I7f42a504fc61c9548acebdd8b1858eaa);
            Ib95e457d5ae9fc89e197c249414abbcd    = I322b3879383d75c43c55535f01fdfdd6;

            I08b1b4639b5a9ca509b943b977f6d4bb = If5dad13ac41b3034bdb034bc86c9b348 + ~Ife6be241bc50560a14f97650e5cc2959 + 1;
            I1adc689464e0b81fa165eb17e71310fa = I2bcab411f9bec1541259751bcb9e0823(I08b1b4639b5a9ca509b943b977f6d4bb);
            I2be28be47a38e9ca9d3b9167327d3d59    = I1adc689464e0b81fa165eb17e71310fa;

            I8d7296627d886566783e79c01b9fa423 = Iac428f9f798618e1ef495c626c41892b + ~Ie04ce30f26a4ef1ee5b34474368dbac7 + 1;
            I2bdc0908c3d365d25f8026263dc4a258 = I2bcab411f9bec1541259751bcb9e0823(I8d7296627d886566783e79c01b9fa423);
            I2ee6154b613d0d86c2354604e93a9a57    = I2bdc0908c3d365d25f8026263dc4a258;

            I4fc4c97229a8b1f631a3b505941159e4 = Iac428f9f798618e1ef495c626c41892b + ~I546657528d591e8bb44c32fed7707af5 + 1;
            Icf6c6fcfa42c48f16a1b30cd325c139f = I2bcab411f9bec1541259751bcb9e0823(I4fc4c97229a8b1f631a3b505941159e4);
            Ia7479d4940b575cf918cb8421f041e44    = Icf6c6fcfa42c48f16a1b30cd325c139f;

            Ib9b16bf51891c328dba2699eb9bcef95 = Iac428f9f798618e1ef495c626c41892b + ~I0ace1d51fdee91f8f3826a945c4e66a4 + 1;
            Ife8337f33629521c096d4dcfde96e879 = I2bcab411f9bec1541259751bcb9e0823(Ib9b16bf51891c328dba2699eb9bcef95);
            I3c5b1cddd608ad869e0182ad68bd0494    = Ife8337f33629521c096d4dcfde96e879;

            I6c30501ec81fce286817788d614a7824 = Iac428f9f798618e1ef495c626c41892b + ~I8dbe6497a8deabcc60783bfe7548d0fb + 1;
            I8afa93d48ae589bb90cc74897defe4de = I2bcab411f9bec1541259751bcb9e0823(I6c30501ec81fce286817788d614a7824);
            Ic4425ae997c479e05e12347a803213dd    = I8afa93d48ae589bb90cc74897defe4de;

            Ia4d4f37baec48121a88808075dd655ef = Iac428f9f798618e1ef495c626c41892b + ~I9a57f2f03cf8a154c3a7d48ec089306d + 1;
            I56d0b4df55f7f4181a51f58187d399e4 = I2bcab411f9bec1541259751bcb9e0823(Ia4d4f37baec48121a88808075dd655ef);
            I3a0518d0d382758ae579acd7e6cd634a    = I56d0b4df55f7f4181a51f58187d399e4;

            I385495ea2bf6442a95ab7561456254ac = Iac428f9f798618e1ef495c626c41892b + ~Icda9a86a25dbe516a93b46fe487029e3 + 1;
            I8ae9260d2a5dd6c2ed4b6157946e38d4 = I2bcab411f9bec1541259751bcb9e0823(I385495ea2bf6442a95ab7561456254ac);
            Ifd28c1cd286b7a483891bdd094b70db1    = I8ae9260d2a5dd6c2ed4b6157946e38d4;

            I5128e03d383c226befa6f7422f3a6f04 = Iac428f9f798618e1ef495c626c41892b + ~I64ae3cd6f36b8bde29cd3e1fcba7bade + 1;
            Ie405c3459c9caf16c0a257a059a9fa96 = I2bcab411f9bec1541259751bcb9e0823(I5128e03d383c226befa6f7422f3a6f04);
            Iadf7734be049c645819d9d023b58c4dc    = Ie405c3459c9caf16c0a257a059a9fa96;

            Ib208908bab4c20713cd17e20139c8db3 = Iac428f9f798618e1ef495c626c41892b + ~Idc4171a40dd2470e852af37a461013c7 + 1;
            Ie76a46f18cbb52a93a4fad65462da3e8 = I2bcab411f9bec1541259751bcb9e0823(Ib208908bab4c20713cd17e20139c8db3);
            I5f23af0d0853ea6de084ccf77702b78d    = Ie76a46f18cbb52a93a4fad65462da3e8;

            Id939992b99a11c09f4688c10ca1a34d1 = I5a6427c8f18b36d2ea18fe60a0831ef1 + ~I43864225be03ea8e9379eb28dfa6c599 + 1;
            I0445dbe40692ef21353aacc7b4f7a4c9 = I2bcab411f9bec1541259751bcb9e0823(Id939992b99a11c09f4688c10ca1a34d1);
            Ic5c99c42e9ebe5dded369ac78a1bedb5    = I0445dbe40692ef21353aacc7b4f7a4c9;

            I823453ccb90d5b2b2d9dfc6e8358224d = I5a6427c8f18b36d2ea18fe60a0831ef1 + ~I70e68beb262fbdeba621b3794adf9f84 + 1;
            Ie3be0f770c8ddbdf301ae23881499e9d = I2bcab411f9bec1541259751bcb9e0823(I823453ccb90d5b2b2d9dfc6e8358224d);
            I4f2498bec0e96802b82f0419d97c527f    = Ie3be0f770c8ddbdf301ae23881499e9d;

            I279c5c00b92eb1b872b5afa168b0306e = I5a6427c8f18b36d2ea18fe60a0831ef1 + ~I656852be6f5b3542862e0f68d48be518 + 1;
            I3a4d175e3b015a17f7a49cc6bacbd12f = I2bcab411f9bec1541259751bcb9e0823(I279c5c00b92eb1b872b5afa168b0306e);
            Icaf86e0abee612aa972388c0b6f90763    = I3a4d175e3b015a17f7a49cc6bacbd12f;

            I66f25b1c3c0eb226295179adcca2c3d2 = I5a6427c8f18b36d2ea18fe60a0831ef1 + ~I041f9455435bfa375395eb330a34993d + 1;
            Id85473220f4909f9182711939cf6a978 = I2bcab411f9bec1541259751bcb9e0823(I66f25b1c3c0eb226295179adcca2c3d2);
            I478c4f13c05651605a2045bb5fd6b60d    = Id85473220f4909f9182711939cf6a978;

            I3068627e91b667d14cd3e55a9371931a = I5a6427c8f18b36d2ea18fe60a0831ef1 + ~Iac48d2ccf6c6e0c555e874ae77123f2e + 1;
            If77ecdb29d692c01752be0908c4f4392 = I2bcab411f9bec1541259751bcb9e0823(I3068627e91b667d14cd3e55a9371931a);
            Ide67911b52687d67ef0c25f2aadf14c5    = If77ecdb29d692c01752be0908c4f4392;

            I44c4e0a2d8a7289f8660b81a9ecfa19b = I5a6427c8f18b36d2ea18fe60a0831ef1 + ~Ib76e892d1a1271844338042381b5690b + 1;
            Ia188482ea4a2696f188f637912aa6f3b = I2bcab411f9bec1541259751bcb9e0823(I44c4e0a2d8a7289f8660b81a9ecfa19b);
            Ie9e7630af25f39a0e820181918edd029    = Ia188482ea4a2696f188f637912aa6f3b;

            Ibe868e258dc87f0dd1460ba6b8354671 = I5a6427c8f18b36d2ea18fe60a0831ef1 + ~I45b64b2b963963d2d0a8318133941f1d + 1;
            Ibd0c9231ee029200ca39013c839bc4ae = I2bcab411f9bec1541259751bcb9e0823(Ibe868e258dc87f0dd1460ba6b8354671);
            I0e1f07f30cfe36f189e9dcb4e713b5c8    = Ibd0c9231ee029200ca39013c839bc4ae;

            Idc3083c3021200345e3edd35a9d4725a = I5a6427c8f18b36d2ea18fe60a0831ef1 + ~I8435e69bc1ff06e7edfabbee7b9aa49e + 1;
            I0fed2eb07a75f701ff7b7ca9dbcddb81 = I2bcab411f9bec1541259751bcb9e0823(Idc3083c3021200345e3edd35a9d4725a);
            I31cee5e2a93635987776b0ea477e6211    = I0fed2eb07a75f701ff7b7ca9dbcddb81;

            I320d4f19a5b18c23ff407508d47caa77 = Icc29441eac6ca7a138d45743d37505e3 + ~Ibfee0b4ad5cdf16e88fcf469c5e031e9 + 1;
            I96140f2ad00cb9a1249b5135ea251bc8 = I2bcab411f9bec1541259751bcb9e0823(I320d4f19a5b18c23ff407508d47caa77);
            I84721f2bc5ae10db78d2e7e07cc28d94    = I96140f2ad00cb9a1249b5135ea251bc8;

            I16becf3c92615d98d5ec51ee9641cc0a = Icc29441eac6ca7a138d45743d37505e3 + ~Ib2afdf9534deaae465d99b7e377788bb + 1;
            I34fecbd6c558b25e7f8d08fb10b224f4 = I2bcab411f9bec1541259751bcb9e0823(I16becf3c92615d98d5ec51ee9641cc0a);
            I6c6d057e910da53aa47441566f95153e    = I34fecbd6c558b25e7f8d08fb10b224f4;

            Ifbfacc3b3a0128119943bcbf80176612 = Icc29441eac6ca7a138d45743d37505e3 + ~Ib6cdbbb765694d822639b7c8fbfc50c4 + 1;
            I8df49bd85a846a4c4c32af63798f3e0e = I2bcab411f9bec1541259751bcb9e0823(Ifbfacc3b3a0128119943bcbf80176612);
            Iecbf70768fbaaab8da98eaa9a2b956ee    = I8df49bd85a846a4c4c32af63798f3e0e;

            I6b4f670c9e8e25984e8891f2440322ab = Icc29441eac6ca7a138d45743d37505e3 + ~I8dddcade21ad3bb330c1c25970c32b73 + 1;
            I05be7b5c657867c4331ed3df72a1aec5 = I2bcab411f9bec1541259751bcb9e0823(I6b4f670c9e8e25984e8891f2440322ab);
            I71b8492d70b423e95938995c07395def    = I05be7b5c657867c4331ed3df72a1aec5;

            I19bf0990a30c72421f231772b8627e8e = Icc29441eac6ca7a138d45743d37505e3 + ~Ib63574478126e6ee30a388d9648cb548 + 1;
            Id47eecb4e17f799da48d80451cb47b5d = I2bcab411f9bec1541259751bcb9e0823(I19bf0990a30c72421f231772b8627e8e);
            Iae469bcbba9598bb46aa7ccf9fa06a37    = Id47eecb4e17f799da48d80451cb47b5d;

            I3ec3eb096ebe3ee8a47e1cba6487b997 = Icc29441eac6ca7a138d45743d37505e3 + ~Ia1aedd38250e76763aaee3de2f832b3c + 1;
            Iedabb8b1ffd46b983fd74b9f6010dcca = I2bcab411f9bec1541259751bcb9e0823(I3ec3eb096ebe3ee8a47e1cba6487b997);
            Ie2e854376f4b6509ec41507401173269    = Iedabb8b1ffd46b983fd74b9f6010dcca;

            I7379ef16405c461ac44b66c4315df831 = Icc29441eac6ca7a138d45743d37505e3 + ~Id5ddf5331aba567aaf5b7eb88b31a52e + 1;
            Ib032a08190a75ceb242a9dc8272b4a02 = I2bcab411f9bec1541259751bcb9e0823(I7379ef16405c461ac44b66c4315df831);
            I7b1401c3c2c389d9bf05658c88ff6b40    = Ib032a08190a75ceb242a9dc8272b4a02;

            I79db45b23d21d533a1f9a6e8f94d403d = Icc29441eac6ca7a138d45743d37505e3 + ~Icb158c031d434cb419c15e0510511231 + 1;
            Ia870db84a0411e463b6e15f502323810 = I2bcab411f9bec1541259751bcb9e0823(I79db45b23d21d533a1f9a6e8f94d403d);
            I88ee95aeb6c744eca0e127e8497b5dc9    = Ia870db84a0411e463b6e15f502323810;

            I0979534730cc2b53547d413dbb6b75f4 = Icc29441eac6ca7a138d45743d37505e3 + ~I79444eef1875b6ad1a0675b66392ff9d + 1;
            I8105600a0847cabdb96310074840bdb7 = I2bcab411f9bec1541259751bcb9e0823(I0979534730cc2b53547d413dbb6b75f4);
            I5573e18ade3430ef3eff5e6d960e44eb    = I8105600a0847cabdb96310074840bdb7;

            I5aa2f9c0667d1a6e871efbd4d2bad3a8 = Icc29441eac6ca7a138d45743d37505e3 + ~Ib88c884e54d6e6ecf5ac015bc304e4f3 + 1;
            I7d6591184fd95d3f288f481734e85c02 = I2bcab411f9bec1541259751bcb9e0823(I5aa2f9c0667d1a6e871efbd4d2bad3a8);
            Id6260fa8a9be077673e82344c736b1c4    = I7d6591184fd95d3f288f481734e85c02;

            Iadb28dc990ccf2dd3099544de16b8f16 = I0e7754dcbc04a4850e052ae4a2fbe328 + ~I31cb0c699cffcd2fedfbed0e1b86490e + 1;
            I69c3d2866b040d67900eeb991b7c2981 = I2bcab411f9bec1541259751bcb9e0823(Iadb28dc990ccf2dd3099544de16b8f16);
            Ic052eadb342350c52d89e73d5fea80bb    = I69c3d2866b040d67900eeb991b7c2981;

            I1f71aebf698788d6ada66891e9ea756f = I0e7754dcbc04a4850e052ae4a2fbe328 + ~I4363ca6b3d9ca9863f70958aa7c23777 + 1;
            Ice61d34abe5e2a9593bfb911da54e959 = I2bcab411f9bec1541259751bcb9e0823(I1f71aebf698788d6ada66891e9ea756f);
            I98b8d024432fc54ebf2f15d99968f2e0    = Ice61d34abe5e2a9593bfb911da54e959;

            Ib234e9cf7e7616a1ebc6ab99df2a7ccb = I0e7754dcbc04a4850e052ae4a2fbe328 + ~I25eb943ea517a4827efb1e797bfdc4f5 + 1;
            I7dfe4eb1588a68b8a35dec39978d06eb = I2bcab411f9bec1541259751bcb9e0823(Ib234e9cf7e7616a1ebc6ab99df2a7ccb);
            I98f54ab8454940141a484332f2a05369    = I7dfe4eb1588a68b8a35dec39978d06eb;

            I297d1edcc583ea4d69da780150f0620c = I0e7754dcbc04a4850e052ae4a2fbe328 + ~I490996026af34eba5bcd8d553af818eb + 1;
            Ica59cc444ecf8f8700bf1ce16a254b89 = I2bcab411f9bec1541259751bcb9e0823(I297d1edcc583ea4d69da780150f0620c);
            I9d94ad2da06ac1fef4da7dcc56abffca    = Ica59cc444ecf8f8700bf1ce16a254b89;

            Ib0a717cbb4fe38a3fc85520ca0826fd9 = I0e7754dcbc04a4850e052ae4a2fbe328 + ~I9d8f8c1792427975a9e7024041f59be9 + 1;
            I0d69f1eb92a8b30d86ffbe0c153197f2 = I2bcab411f9bec1541259751bcb9e0823(Ib0a717cbb4fe38a3fc85520ca0826fd9);
            I51262e3abe460148e3c2d2b74989c2b8    = I0d69f1eb92a8b30d86ffbe0c153197f2;

            I037ecd5945b1f1280b4469d73fe1c7ff = I0e7754dcbc04a4850e052ae4a2fbe328 + ~I452ba61d5fb5c7ead1824dade4bd7801 + 1;
            I5a48ea253b357c8e6441be01918bc57c = I2bcab411f9bec1541259751bcb9e0823(I037ecd5945b1f1280b4469d73fe1c7ff);
            I560583680bb2f5a0b5ede42ceaafcf8b    = I5a48ea253b357c8e6441be01918bc57c;

            I367ff6b11b884e02a3065fc7fe811e15 = I0e7754dcbc04a4850e052ae4a2fbe328 + ~I7e36dcae438a712fca2320117b7e3356 + 1;
            Ic3c81f609bf98f2ded891b55bacbd453 = I2bcab411f9bec1541259751bcb9e0823(I367ff6b11b884e02a3065fc7fe811e15);
            I389f83346ffaffe8186fb0074d71f43c    = Ic3c81f609bf98f2ded891b55bacbd453;

            I6fab19692b512166fe9c74b5e987788d = I0e7754dcbc04a4850e052ae4a2fbe328 + ~Ifc527b6af9486df7f52d7eb9637c671f + 1;
            Ie38b3f5ad91f2c983d519c9b1200559c = I2bcab411f9bec1541259751bcb9e0823(I6fab19692b512166fe9c74b5e987788d);
            Ie89c2a1b3943d12197bb972bd12595b0    = Ie38b3f5ad91f2c983d519c9b1200559c;

            I04dd73af505f618ccdb209b3cf97ceec = I0e7754dcbc04a4850e052ae4a2fbe328 + ~I1062442edb2bff727ca6283c8270bf28 + 1;
            I1e5e2679a0e75104cc0be107ecadd01c = I2bcab411f9bec1541259751bcb9e0823(I04dd73af505f618ccdb209b3cf97ceec);
            Ic7be56919976a2d1088114c21c3c1ffb    = I1e5e2679a0e75104cc0be107ecadd01c;

            If8c559905d4120488d431719c4e8ce24 = I0e7754dcbc04a4850e052ae4a2fbe328 + ~I2959f2dc554e599d675eb6912757e413 + 1;
            I903e174feff2be7109cdb19fa15a63ec = I2bcab411f9bec1541259751bcb9e0823(If8c559905d4120488d431719c4e8ce24);
            Icb5dab0df062ab46bd3d1a73e85ef4c2    = I903e174feff2be7109cdb19fa15a63ec;

            I20ed4f6f14e20ce3f0e106d1b7782fcd = Ia30c019ed8ce395556494a92e7b42a92 + ~I4d4ec5540257040d10182ed478a71918 + 1;
            I6893d09bc4fca46b4ad33c42d1950790 = I2bcab411f9bec1541259751bcb9e0823(I20ed4f6f14e20ce3f0e106d1b7782fcd);
            I27a568cfc2df13cf689d366a25e5d05f    = I6893d09bc4fca46b4ad33c42d1950790;

            Ib10626ffa126188c5bf1fc8399107b26 = Ia30c019ed8ce395556494a92e7b42a92 + ~Ifef870b405335975988b58b2273d4e1a + 1;
            I4ec84e063fb84d278ae90b84751b1bcc = I2bcab411f9bec1541259751bcb9e0823(Ib10626ffa126188c5bf1fc8399107b26);
            Ia6688964078f1ea87b742352877aac45    = I4ec84e063fb84d278ae90b84751b1bcc;

            I29007c52357ac7afbda39d72a5bb60af = Ia30c019ed8ce395556494a92e7b42a92 + ~I9e0a36d0be66b4c02b03e5b75b686226 + 1;
            I33998829023b087dbfa2e568d77291b3 = I2bcab411f9bec1541259751bcb9e0823(I29007c52357ac7afbda39d72a5bb60af);
            I180deab4fe0d03104cf2ee035f6a9b8c    = I33998829023b087dbfa2e568d77291b3;

            I66d367c046611f145e607a90911cf499 = Ia30c019ed8ce395556494a92e7b42a92 + ~If404a00ab81d6ebbc0dbdf4aecdce389 + 1;
            I5bc68432bc0a9ea8cd024d7fc3d3fdc8 = I2bcab411f9bec1541259751bcb9e0823(I66d367c046611f145e607a90911cf499);
            Iff6cd034bb64d13c21910c11bd92266e    = I5bc68432bc0a9ea8cd024d7fc3d3fdc8;

            I9c4c2556f6170a8df61d909855a846ed = Ia30c019ed8ce395556494a92e7b42a92 + ~Ic6f40833f5f6284c9015304fd3fc00f0 + 1;
            Ib84e5271ffa3584148ce87dcf2a4f2a2 = I2bcab411f9bec1541259751bcb9e0823(I9c4c2556f6170a8df61d909855a846ed);
            I7c34057a77f2bdda93c422506959818d    = Ib84e5271ffa3584148ce87dcf2a4f2a2;

            I6fadc3e8d995bb4317bf7b4377c3c2c5 = Ia30c019ed8ce395556494a92e7b42a92 + ~Ib8664a2abe9d6326d6e45bb2a7ad59d0 + 1;
            Ib633998a5fd0df508b47ba9c2f7c390a = I2bcab411f9bec1541259751bcb9e0823(I6fadc3e8d995bb4317bf7b4377c3c2c5);
            I7ff7d3fd63fa67cd72d1591c1a373180    = Ib633998a5fd0df508b47ba9c2f7c390a;

            I99b20e911c189e0616f02376ab736e91 = Ia30c019ed8ce395556494a92e7b42a92 + ~I36ed1a0d0d618f90443fbea17b7c97ec + 1;
            Ie36cfd3519810d325d5cdc5150380fe0 = I2bcab411f9bec1541259751bcb9e0823(I99b20e911c189e0616f02376ab736e91);
            If910e75bf10cf02a5b414cbb4fad1304    = Ie36cfd3519810d325d5cdc5150380fe0;

            I5793c12f5dbdd8245dbb202d550ca960 = Ia30c019ed8ce395556494a92e7b42a92 + ~I397a69dab323c7148b620dd6fe0b0c51 + 1;
            I6ac3755ff9de4d43d0493891b2a5758d = I2bcab411f9bec1541259751bcb9e0823(I5793c12f5dbdd8245dbb202d550ca960);
            I266697a6eca2b73a76fd375a0ad72a05    = I6ac3755ff9de4d43d0493891b2a5758d;

            Id0660e9637cad1ce1a73d37188060154 = Ia30c019ed8ce395556494a92e7b42a92 + ~Ifae488cb68d95ea517376319eb11f1bf + 1;
            I5f0212d2ffe8f85614891882390bbc25 = I2bcab411f9bec1541259751bcb9e0823(Id0660e9637cad1ce1a73d37188060154);
            Iba188abd7715fcbdad3b1f3d985c6fc3    = I5f0212d2ffe8f85614891882390bbc25;

            If5a7af7ca023e1393526e888f4220a44 = Ia30c019ed8ce395556494a92e7b42a92 + ~I10f045edf47784a91a5599494c2d3de2 + 1;
            I1e009fcbec9031954637f055cb9cfe01 = I2bcab411f9bec1541259751bcb9e0823(If5a7af7ca023e1393526e888f4220a44);
            Ic60c640562e3e45c89a1de78af509b6a    = I1e009fcbec9031954637f055cb9cfe01;

            Id043eb50634e803e53adc1168379a5d0 = I9799695ea8244992a6694eaf5c8ae64d + ~If0c2d002c315b21e11ae776bb48c9338 + 1;
            Ia6caeb0fcc8e7486e4d55b72a0d499a5 = I2bcab411f9bec1541259751bcb9e0823(Id043eb50634e803e53adc1168379a5d0);
            I0456494b33e4ec852c123cb3003b9886    = Ia6caeb0fcc8e7486e4d55b72a0d499a5;

            I1f866dd0b129267550aea1a267d9c91e = I9799695ea8244992a6694eaf5c8ae64d + ~Ifbe29365e7035c78af9f42902b0d303e + 1;
            I631e31da7dccd5b9311a4fa73e6a0227 = I2bcab411f9bec1541259751bcb9e0823(I1f866dd0b129267550aea1a267d9c91e);
            I2ed7c217fe3e21fcb27e04f68b95dd6b    = I631e31da7dccd5b9311a4fa73e6a0227;

            I8c4da05c08210fe33139c3d3e5d75d58 = I9799695ea8244992a6694eaf5c8ae64d + ~I6922b510e432e06d209095bcc6297e7e + 1;
            Ib152eea9af905931ab45c4f9d89fa50b = I2bcab411f9bec1541259751bcb9e0823(I8c4da05c08210fe33139c3d3e5d75d58);
            Ifda5780b42bf451a7ce834f17b3fdd20    = Ib152eea9af905931ab45c4f9d89fa50b;

            Ib41f7b823681fdd084b6d8436a407aa8 = I9799695ea8244992a6694eaf5c8ae64d + ~I31bf4597a3b776962f5c820378254065 + 1;
            I94118c50e80e5fed4294d16358d41579 = I2bcab411f9bec1541259751bcb9e0823(Ib41f7b823681fdd084b6d8436a407aa8);
            Iadca92fd39d1fd6032feb8415ca5246f    = I94118c50e80e5fed4294d16358d41579;

            Ic5b50a785b7acac7e3be4095aa92e50a = I9799695ea8244992a6694eaf5c8ae64d + ~Ic3e6e38a2986c7f14fd0db2246367a1c + 1;
            I1269d97f8ab4f5dddc002acf38b4a189 = I2bcab411f9bec1541259751bcb9e0823(Ic5b50a785b7acac7e3be4095aa92e50a);
            I613453382f19dd7eb9bdf51e945a33b0    = I1269d97f8ab4f5dddc002acf38b4a189;

            I3ffbe03796b66d00d47fd918be60ab89 = I9799695ea8244992a6694eaf5c8ae64d + ~Ia1d9dee7a9821283498d17de0cfacb32 + 1;
            I89a793ddaf4887ddb8dbaaba13225d08 = I2bcab411f9bec1541259751bcb9e0823(I3ffbe03796b66d00d47fd918be60ab89);
            Ideafa683e6a3a38848fb8bee22eba11b    = I89a793ddaf4887ddb8dbaaba13225d08;

            Ifc92a916da938ef6164db250be635f88 = I9799695ea8244992a6694eaf5c8ae64d + ~Ibac0851ce1a3c23f18b072d263afff36 + 1;
            I2b4fe952791866aecbbbcf01257d527b = I2bcab411f9bec1541259751bcb9e0823(Ifc92a916da938ef6164db250be635f88);
            Ie4226e7e17c7971f07aaf0cfaeae495a    = I2b4fe952791866aecbbbcf01257d527b;

            I8ccd42508ce7d5bd897c2cf0c54caeb3 = I9799695ea8244992a6694eaf5c8ae64d + ~I53971b75cbd7ebc74b579776a6ea4778 + 1;
            I797321bb9e3c2d7d3727af9a4cf5418b = I2bcab411f9bec1541259751bcb9e0823(I8ccd42508ce7d5bd897c2cf0c54caeb3);
            Ifbbfa268bd4c31c7eed45cd43fe6a405    = I797321bb9e3c2d7d3727af9a4cf5418b;

            I4920e7e82749cc036b58a7cd0a03e327 = I9799695ea8244992a6694eaf5c8ae64d + ~Ibeff607ba15fd8ef504224a9c1d102fc + 1;
            I5eeb78b1511aa7b76765d82328323a4c = I2bcab411f9bec1541259751bcb9e0823(I4920e7e82749cc036b58a7cd0a03e327);
            Ib2d99d95f7a31e4745211c5ff96f851c    = I5eeb78b1511aa7b76765d82328323a4c;

            Ie1040b2aa91f272e4449c4b5f9f8f575 = I9799695ea8244992a6694eaf5c8ae64d + ~I4ae2f2330a8ee7d5626499f2a030c7a5 + 1;
            I55f8232fcfcb929a35717f724f44eb4c = I2bcab411f9bec1541259751bcb9e0823(Ie1040b2aa91f272e4449c4b5f9f8f575);
            I692c0a91b415b400a3640e2d9a40edad    = I55f8232fcfcb929a35717f724f44eb4c;

            I65968fb0f63d52ad96cd8fa270126a1b = I4524cd664b4cb41f642c675fa484c84b + ~I8da7e01f56dc9a70eb6b3f110dc005c2 + 1;
            I7a7705607e93fca1cf1e7b1c92c4e3cc = I2bcab411f9bec1541259751bcb9e0823(I65968fb0f63d52ad96cd8fa270126a1b);
            If8c4dc70212e8873167e1cad8e8e5692    = I7a7705607e93fca1cf1e7b1c92c4e3cc;

            I839ac8ee59f51d4c3de92ba5cb26e788 = I4524cd664b4cb41f642c675fa484c84b + ~I005e8b590924f9486cb23191d35c9797 + 1;
            I7e2e0ffb2b5622ba6e03a47755a9a1dc = I2bcab411f9bec1541259751bcb9e0823(I839ac8ee59f51d4c3de92ba5cb26e788);
            Ib2f75e91bf9e1d32a3f170fc85244139    = I7e2e0ffb2b5622ba6e03a47755a9a1dc;

            I33cd95f1919318a0f3df5df7310d64c6 = I4524cd664b4cb41f642c675fa484c84b + ~Ic1f6842b4f246d624d91daa6ada10ca9 + 1;
            I5f50e835526833015a2087dbdb77686e = I2bcab411f9bec1541259751bcb9e0823(I33cd95f1919318a0f3df5df7310d64c6);
            I3606dc61f24567cb1ace443cea62a43b    = I5f50e835526833015a2087dbdb77686e;

            I4933e8d16fba26cd797b25a9ac2a2de8 = I4524cd664b4cb41f642c675fa484c84b + ~Ief90f8a8efca2b06eff0d4cba1cbb342 + 1;
            I98f32439ec64d796ebb157815b259aa2 = I2bcab411f9bec1541259751bcb9e0823(I4933e8d16fba26cd797b25a9ac2a2de8);
            Ie402c9f793b7306323efb8fe23533250    = I98f32439ec64d796ebb157815b259aa2;

            I218f7578eb748e31d0002052f30c5842 = I4524cd664b4cb41f642c675fa484c84b + ~I0f46a17f14ab18e6338aa3d06678b0a5 + 1;
            Id59ca1b1cff93a8544c54c6d4ee22b2f = I2bcab411f9bec1541259751bcb9e0823(I218f7578eb748e31d0002052f30c5842);
            I54652565023310e2eccfc4cb87c56b43    = Id59ca1b1cff93a8544c54c6d4ee22b2f;

            I2a808d1c42ad758ae3baaaee8129dfb2 = I4524cd664b4cb41f642c675fa484c84b + ~Ia3bfd86e26efbef2cf6bb72be7ac1453 + 1;
            I726538434626c5202d53d29faedddd56 = I2bcab411f9bec1541259751bcb9e0823(I2a808d1c42ad758ae3baaaee8129dfb2);
            I616b7a5987edbc001e0ae1b638f25a39    = I726538434626c5202d53d29faedddd56;

            I4e851fd3c114af87f5e8c68c02594e3a = I4524cd664b4cb41f642c675fa484c84b + ~If6f5efee5e1f9709d86bf28cfb741955 + 1;
            I8ea236c734f7b96620a37750134d3872 = I2bcab411f9bec1541259751bcb9e0823(I4e851fd3c114af87f5e8c68c02594e3a);
            I06604bac478ee906b3fe8ff307cdf046    = I8ea236c734f7b96620a37750134d3872;

            I0da40f88adc46e90f616acdcdb8e0e2c = I4524cd664b4cb41f642c675fa484c84b + ~I60520c850a95b893528569c4069bd677 + 1;
            I259d7244226dbcbd1d02df5ca164afdc = I2bcab411f9bec1541259751bcb9e0823(I0da40f88adc46e90f616acdcdb8e0e2c);
            I135dd8a85aca863db660f2ad4f80ca2e    = I259d7244226dbcbd1d02df5ca164afdc;

            I0dee7767e472a5fd71250ae6c57cc8b5 = I64e959d80af111ed2fcd54a5407d21bf + ~I18e548b082364c75686f2b7ad2ef46ab + 1;
            I086375f289b769938edfc8b9b5146714 = I2bcab411f9bec1541259751bcb9e0823(I0dee7767e472a5fd71250ae6c57cc8b5);
            I8715d73b58270dfa33b903e9cfb50be8    = I086375f289b769938edfc8b9b5146714;

            I9f40be7552b3dd625e5bce0befc5a548 = I64e959d80af111ed2fcd54a5407d21bf + ~I6e4ae763dc4e8aa8afc4599de96c75d3 + 1;
            Icb82f8092f14511d62f7cbe821af9faf = I2bcab411f9bec1541259751bcb9e0823(I9f40be7552b3dd625e5bce0befc5a548);
            I7f60cb59895af6d314f5d0f401c80350    = Icb82f8092f14511d62f7cbe821af9faf;

            I8fdf98ffd757c8845ed6ffa4ddd1a16b = I64e959d80af111ed2fcd54a5407d21bf + ~Ic8759e2f58848b33082bd1b02acc9c0b + 1;
            I7e8df00362c29bd3924ecbe3dd1db23c = I2bcab411f9bec1541259751bcb9e0823(I8fdf98ffd757c8845ed6ffa4ddd1a16b);
            I3e25e6e9de5ee9242a472ce957056762    = I7e8df00362c29bd3924ecbe3dd1db23c;

            I8103b777314a4fa471e0898fde9cde08 = I64e959d80af111ed2fcd54a5407d21bf + ~Ibdaa6d215d34aa0cc27d5234da6fd991 + 1;
            If1014cbbd6e267aaacbcf3c8ba33a98b = I2bcab411f9bec1541259751bcb9e0823(I8103b777314a4fa471e0898fde9cde08);
            I4c5f36517aaf872e7f05de2f7f76a6ce    = If1014cbbd6e267aaacbcf3c8ba33a98b;

            If6c3ee8e0d7dea58043d5be0f4630873 = I64e959d80af111ed2fcd54a5407d21bf + ~I0f9bc36c9d40290f83489aac3d674924 + 1;
            Iae4dfe3ede67923e8b740dd575b216b6 = I2bcab411f9bec1541259751bcb9e0823(If6c3ee8e0d7dea58043d5be0f4630873);
            I0e993e6f98616632f17835a2994f45e3    = Iae4dfe3ede67923e8b740dd575b216b6;

            I711a5171f591f472cdbfc9a0f5e1aa17 = I64e959d80af111ed2fcd54a5407d21bf + ~I9a2bba3f62de5f750dc8161a488dc331 + 1;
            Iccfddf46ea48242ca751b5d53f98d270 = I2bcab411f9bec1541259751bcb9e0823(I711a5171f591f472cdbfc9a0f5e1aa17);
            I281f996740b16568b9d29ca41a3fa50d    = Iccfddf46ea48242ca751b5d53f98d270;

            Ic30bc38184dfbbd694af52640692709d = I64e959d80af111ed2fcd54a5407d21bf + ~I898d1b59aab3d5d4adce8ec3c0e14a0d + 1;
            I804705ac9a613b4107c8ceaac4127386 = I2bcab411f9bec1541259751bcb9e0823(Ic30bc38184dfbbd694af52640692709d);
            I55bbb73d68871d9dbce4d590c029aeab    = I804705ac9a613b4107c8ceaac4127386;

            I422f6fd1d273a3834d04b04ab8e2812d = I64e959d80af111ed2fcd54a5407d21bf + ~Ic92ab3dac1a151d6ff0b4e0c21003eb0 + 1;
            I8f40972503fbfdab92676a32f351dfe6 = I2bcab411f9bec1541259751bcb9e0823(I422f6fd1d273a3834d04b04ab8e2812d);
            Ida491561008f4984480d1b0f09d2fa77    = I8f40972503fbfdab92676a32f351dfe6;

            Ia0fdc60b90ad18b6585ec1ad4e89e80b = I3e0da4bcbab4804b5397fb3aa2c94f51 + ~I3a4a965f22487553dec2a3e8e7836264 + 1;
            I8fc9ec077c7c6ce5e2660a4530a234ae = I2bcab411f9bec1541259751bcb9e0823(Ia0fdc60b90ad18b6585ec1ad4e89e80b);
            I624e237f248d292c0417ff85056857b0    = I8fc9ec077c7c6ce5e2660a4530a234ae;

            I7809fe7a30d041a7e569ffe890242df8 = I3e0da4bcbab4804b5397fb3aa2c94f51 + ~Ie7bf11bab3d601fd0a6e3eb415e263c8 + 1;
            I3e3bf3c2155f584784863ae41cb73c7d = I2bcab411f9bec1541259751bcb9e0823(I7809fe7a30d041a7e569ffe890242df8);
            Ic7c1fd79ba76dbb254c6183017f40b3e    = I3e3bf3c2155f584784863ae41cb73c7d;

            I672b14ec1b3c4797545f266727505a85 = I3e0da4bcbab4804b5397fb3aa2c94f51 + ~I6eaffd980e4d77fdbda5e63bad9489d7 + 1;
            I9cc24d95a0ddbe4145d144003778eebc = I2bcab411f9bec1541259751bcb9e0823(I672b14ec1b3c4797545f266727505a85);
            I546d683af76dc209a5205c6274abe908    = I9cc24d95a0ddbe4145d144003778eebc;

            If9620d20ebaae6245a2c386d9bf5fdb1 = I3e0da4bcbab4804b5397fb3aa2c94f51 + ~Iac4b8906947fc90bfe76cee2f1d4c4ab + 1;
            Ib9b96de1e217660c2ac9f7815249c6a2 = I2bcab411f9bec1541259751bcb9e0823(If9620d20ebaae6245a2c386d9bf5fdb1);
            I7b4bb785489c5bb22c84d9778192fe44    = Ib9b96de1e217660c2ac9f7815249c6a2;

            Ic74e22bffd88f32eefe499cde0fafa8a = I3e0da4bcbab4804b5397fb3aa2c94f51 + ~I612a41511db375f10f3c2b10d13edb24 + 1;
            I2cc498e11d3d487d1e8319df8521ff6d = I2bcab411f9bec1541259751bcb9e0823(Ic74e22bffd88f32eefe499cde0fafa8a);
            Ifc6af7d7aeb7162d554b8604a44f3361    = I2cc498e11d3d487d1e8319df8521ff6d;

            I76d38ce67387bd76ab45c9cba7d18b31 = I3e0da4bcbab4804b5397fb3aa2c94f51 + ~Ia6a78664c080829664158f53ba330312 + 1;
            Iae3d8158d13c8179719cbe12fdd7f9ab = I2bcab411f9bec1541259751bcb9e0823(I76d38ce67387bd76ab45c9cba7d18b31);
            I5b650c4c3291670b480a7f1095093dfb    = Iae3d8158d13c8179719cbe12fdd7f9ab;

            I44413c6f6f6493f8a86abf6eb32604f6 = I3e0da4bcbab4804b5397fb3aa2c94f51 + ~I6a81b4485598387e4656c35e83866209 + 1;
            Ieadf1b0e427ecddd261297ae4054a0bd = I2bcab411f9bec1541259751bcb9e0823(I44413c6f6f6493f8a86abf6eb32604f6);
            I2f5f88cb5e5e4723bd8a83c5fa80cc4c    = Ieadf1b0e427ecddd261297ae4054a0bd;

            I67f632fca617fe06565ddcaaee8fa8b8 = I3e0da4bcbab4804b5397fb3aa2c94f51 + ~Ifb09b84f9681c7bc28ffd562b633ffd9 + 1;
            I8dbe4e03db655e1f691254835fb58798 = I2bcab411f9bec1541259751bcb9e0823(I67f632fca617fe06565ddcaaee8fa8b8);
            Ic174b361182c98486e65b7f87b073274    = I8dbe4e03db655e1f691254835fb58798;

            I3fd38a71ce6aa3db1d7a5a9f8a991e12 = I3740b30d31f3c61d93a14a46e3199c4d + ~Ibed5004d869a01005768ba694c2234d6 + 1;
            I14b22818be28bc385f91920399012555 = I2bcab411f9bec1541259751bcb9e0823(I3fd38a71ce6aa3db1d7a5a9f8a991e12);
            I7ba2f7201745258dbf224de087a25233    = I14b22818be28bc385f91920399012555;

            I63e5718bf7d8771ef90b91be73d73264 = I3740b30d31f3c61d93a14a46e3199c4d + ~I91c2f3cdd7cc98a60090ec6e46d52ae7 + 1;
            Id2878a17128a23eee2272c7e39743bd3 = I2bcab411f9bec1541259751bcb9e0823(I63e5718bf7d8771ef90b91be73d73264);
            I131a4bd335fc23ee10f7ccb1881ab9cd    = Id2878a17128a23eee2272c7e39743bd3;

            Ie385e1aeb2b0dcf6d2454be3d7708b27 = I3740b30d31f3c61d93a14a46e3199c4d + ~Ic902e09b33db1b919c102f7971cdef7b + 1;
            I3701d2d2e74c43b3ae347902c0efff20 = I2bcab411f9bec1541259751bcb9e0823(Ie385e1aeb2b0dcf6d2454be3d7708b27);
            I90cb3e06b42f25956b788a792eef371f    = I3701d2d2e74c43b3ae347902c0efff20;

            Ib2d1b7e105b25b492b45da72536d7578 = I3740b30d31f3c61d93a14a46e3199c4d + ~I1eef40a71c8d1e2da9802929a5347e90 + 1;
            Id6487b559b7ebad725aa43382f09bab3 = I2bcab411f9bec1541259751bcb9e0823(Ib2d1b7e105b25b492b45da72536d7578);
            I56302770a8d56932e7bb5dcff56c71e2    = Id6487b559b7ebad725aa43382f09bab3;

            I588abf5ef4c583f0fec422736a0ce6a0 = I3740b30d31f3c61d93a14a46e3199c4d + ~Id58474582f209a3859f65a447fe99191 + 1;
            Ib6ea830665d44628aef5041b2fa46328 = I2bcab411f9bec1541259751bcb9e0823(I588abf5ef4c583f0fec422736a0ce6a0);
            Id3b8c058b3838c388eb5ddcb31dfc799    = Ib6ea830665d44628aef5041b2fa46328;

            I58bb95c56c7be17c263a2161210d7d8d = I3740b30d31f3c61d93a14a46e3199c4d + ~I1939152ddbede923cde577984e0aa743 + 1;
            Ia6181e1acc2ea46a85626a22983e2662 = I2bcab411f9bec1541259751bcb9e0823(I58bb95c56c7be17c263a2161210d7d8d);
            I7ca8ce63dfb821d10304958bada71737    = Ia6181e1acc2ea46a85626a22983e2662;

            Ifaf0e1f21b3bd7393c475b5126540a72 = I3740b30d31f3c61d93a14a46e3199c4d + ~I4aa98503fc71292d42dba1cab6db952f + 1;
            I8b38fb1f95f036393933d07e0a60b875 = I2bcab411f9bec1541259751bcb9e0823(Ifaf0e1f21b3bd7393c475b5126540a72);
            I06ad44414b45d262f9542015d2dead8d    = I8b38fb1f95f036393933d07e0a60b875;

            I7027db9e0450724a6d417d708f1043f2 = I3740b30d31f3c61d93a14a46e3199c4d + ~I8ce945d9f70bb317064a8d2d4eafd2d3 + 1;
            I33d76ad1185bbf80de5e8ff0ad52b15f = I2bcab411f9bec1541259751bcb9e0823(I7027db9e0450724a6d417d708f1043f2);
            I833ef4acfed17e4699d65cbaa3e7dbd5    = I33d76ad1185bbf80de5e8ff0ad52b15f;

            Iebcb7206d8860b5094459c5d10b4efed = Ibf0a30abfec9031737eada436ac1a0d4 + ~Ica3d4ebff001fb6ee69a66eb898eb5bd + 1;
            If2c522a90684b77b18f0058d1d2b14d8 = I2bcab411f9bec1541259751bcb9e0823(Iebcb7206d8860b5094459c5d10b4efed);
            Ia77e3db939408af719e0a8555dcb68ed    = If2c522a90684b77b18f0058d1d2b14d8;

            I6bbf2b47a7dc50e66a3d8d258d6e31fb = Ibf0a30abfec9031737eada436ac1a0d4 + ~I99ff3922e018c409dc8ce5f3503e3c56 + 1;
            I869e040de179572cdfd9373a4de8b31c = I2bcab411f9bec1541259751bcb9e0823(I6bbf2b47a7dc50e66a3d8d258d6e31fb);
            I57ab4999187992eda55a82bf0f09b31f    = I869e040de179572cdfd9373a4de8b31c;

            I8459abaa907f5afcd11884b1ec8c06c5 = Ibf0a30abfec9031737eada436ac1a0d4 + ~I58a490344f87b4d5bb319e3e85ba9278 + 1;
            I3fb8890ee1f1cb30ecdf50d69e4ac0fa = I2bcab411f9bec1541259751bcb9e0823(I8459abaa907f5afcd11884b1ec8c06c5);
            I21f7b5402ae8e8954d99931bd5108250    = I3fb8890ee1f1cb30ecdf50d69e4ac0fa;

            Ia16ae2f6ef5000d47b6b84ed058252aa = Ibf0a30abfec9031737eada436ac1a0d4 + ~I58361fb97f1b5aff0a2751d35c8da672 + 1;
            I6b60e2478c009889776de20209929ee0 = I2bcab411f9bec1541259751bcb9e0823(Ia16ae2f6ef5000d47b6b84ed058252aa);
            I3627708869b47d460182bc5040092f9a    = I6b60e2478c009889776de20209929ee0;

            Ica32690dbc9ea110fefdce92260b125c = Ibf0a30abfec9031737eada436ac1a0d4 + ~I581eb136fdd08302e02c1fafb5d5c90b + 1;
            Ie6b559c2f0bd388d072b660341eebe31 = I2bcab411f9bec1541259751bcb9e0823(Ica32690dbc9ea110fefdce92260b125c);
            Ifd88f0f0abd1c037434dc16e34550d2a    = Ie6b559c2f0bd388d072b660341eebe31;

            Ic431d9383cce30b1889c92e2be4cb9d0 = Ibf0a30abfec9031737eada436ac1a0d4 + ~I91893028c4409cfeceeb7976815b2d31 + 1;
            Ia46aa3a3e6a01d4690dfe0e7f1eab548 = I2bcab411f9bec1541259751bcb9e0823(Ic431d9383cce30b1889c92e2be4cb9d0);
            I27eec53da48406e7e1202345a0810e08    = Ia46aa3a3e6a01d4690dfe0e7f1eab548;

            Ib9cca4c0e58373c26d5fd9f51f793898 = Ibf0a30abfec9031737eada436ac1a0d4 + ~I19032091a26dfdfffff60818041ec79e + 1;
            Idb7244908662bcd97fe8fe0db4b1abdc = I2bcab411f9bec1541259751bcb9e0823(Ib9cca4c0e58373c26d5fd9f51f793898);
            I682d42afaaf103550ce4fbdba6192c88    = Idb7244908662bcd97fe8fe0db4b1abdc;

            I99bf0bc8ac20832b3724b2753f6ca449 = Ibf0a30abfec9031737eada436ac1a0d4 + ~I563802213afb6abe2f6e8c6f4d1e5b08 + 1;
            If570b3495ea5b3f250cf4873f5dd0bb9 = I2bcab411f9bec1541259751bcb9e0823(I99bf0bc8ac20832b3724b2753f6ca449);
            If225534847db8723768941c3819ed7c0    = If570b3495ea5b3f250cf4873f5dd0bb9;

            Ie701008f3c60c51ed72c5f964a8fc36e = Ibf0a30abfec9031737eada436ac1a0d4 + ~I4ae59dd2f57bda295e11b077e8668f1a + 1;
            I50bbcccc40af5e9700b97e682953c8c9 = I2bcab411f9bec1541259751bcb9e0823(Ie701008f3c60c51ed72c5f964a8fc36e);
            I43a91b2232a47d1f6731bafc15ced5db    = I50bbcccc40af5e9700b97e682953c8c9;

            I3e2d78f8307a1787f8b2eccba94c7557 = Ibf0a30abfec9031737eada436ac1a0d4 + ~If525ac3dc97e3187e036d70e9984939d + 1;
            I5422f11a7e0b646dd4fa254602f91b34 = I2bcab411f9bec1541259751bcb9e0823(I3e2d78f8307a1787f8b2eccba94c7557);
            Ic54026604afd19b0c7c71ea1ac0f1c4e    = I5422f11a7e0b646dd4fa254602f91b34;

            Ic1b4444ab0df9745d29bf893d9b83168 = Id36e8953a02400a5ab1f4dfdb0422e6d + ~I4254f2987cd014ed703ae18e9963e585 + 1;
            Ic5c34f86b03fffdcf723ff4116822e3f = I2bcab411f9bec1541259751bcb9e0823(Ic1b4444ab0df9745d29bf893d9b83168);
            I218bd69f079aa21f0dda241ae6e387ad    = Ic5c34f86b03fffdcf723ff4116822e3f;

            I5f52dbf600656a8f5dc6b6b8a45ccebe = Id36e8953a02400a5ab1f4dfdb0422e6d + ~Id6551b6b053952162b90792ab73a1a49 + 1;
            I2ebd72fb063702a7c36b4b546f4b94b8 = I2bcab411f9bec1541259751bcb9e0823(I5f52dbf600656a8f5dc6b6b8a45ccebe);
            Iaaacca4d06ad0f202d839fd7674f1829    = I2ebd72fb063702a7c36b4b546f4b94b8;

            I7f307af79f45ad4b9511e3961c917078 = Id36e8953a02400a5ab1f4dfdb0422e6d + ~Ied41909cd443432dafadba42672151c1 + 1;
            I6328eca7325eea20ccf30adf8b928edb = I2bcab411f9bec1541259751bcb9e0823(I7f307af79f45ad4b9511e3961c917078);
            Iecddac410bb2121da0df2d73c2d23cb8    = I6328eca7325eea20ccf30adf8b928edb;

            Ie17a5be2a16d2efb98c976d7ee882535 = Id36e8953a02400a5ab1f4dfdb0422e6d + ~I74a7b85ddacad06ab1c6b0db9b084bd3 + 1;
            Ica13fd6daec896ddb0fa6be797edf6bb = I2bcab411f9bec1541259751bcb9e0823(Ie17a5be2a16d2efb98c976d7ee882535);
            I1aabc0c0b7b602297ad592ae48b23452    = Ica13fd6daec896ddb0fa6be797edf6bb;

            I5f19d2adff2f34a4bebe03f929a09c49 = Id36e8953a02400a5ab1f4dfdb0422e6d + ~Ic4501a8a1fb34c30a97e18a0ab189e3a + 1;
            I970c832cf68b5178f3d8111c9fed3b5a = I2bcab411f9bec1541259751bcb9e0823(I5f19d2adff2f34a4bebe03f929a09c49);
            Ida3aaf7237b1383cfe95eeccf3971a8e    = I970c832cf68b5178f3d8111c9fed3b5a;

            I3cd69aeed9e869a2096d6dced5c209a0 = Id36e8953a02400a5ab1f4dfdb0422e6d + ~Idd8643af2515f65fd9a1dfe66494ccf2 + 1;
            I65f78ccc122f96f97fee54955d370288 = I2bcab411f9bec1541259751bcb9e0823(I3cd69aeed9e869a2096d6dced5c209a0);
            Idd2a8ed39edf6697b0988ee4eb4f2d95    = I65f78ccc122f96f97fee54955d370288;

            I359b6a22c9568a13b81670c741281393 = Id36e8953a02400a5ab1f4dfdb0422e6d + ~Ic9e06a355beabfacc053ec48f17f49de + 1;
            I5f77d7804a3e4adb641908be74f3ea19 = I2bcab411f9bec1541259751bcb9e0823(I359b6a22c9568a13b81670c741281393);
            I735c660d5232e03dd8fb129e2ca4b445    = I5f77d7804a3e4adb641908be74f3ea19;

            I24ba99614df383c38bbac50ae8b4487e = Id36e8953a02400a5ab1f4dfdb0422e6d + ~I31d94aae2e3721045fe850d84dd2225a + 1;
            I9263e4ab78ca05f93ff921c4fd9ff787 = I2bcab411f9bec1541259751bcb9e0823(I24ba99614df383c38bbac50ae8b4487e);
            Ia04d6065987df3f007658614406cbc28    = I9263e4ab78ca05f93ff921c4fd9ff787;

            I7498bee46de6b1c946ce95fdcc89f6e5 = Id36e8953a02400a5ab1f4dfdb0422e6d + ~I71da7e172b2b967040b6e6d02ef9949e + 1;
            I6f8f253cfb1fe1c2254e557f732a9b22 = I2bcab411f9bec1541259751bcb9e0823(I7498bee46de6b1c946ce95fdcc89f6e5);
            I7aeddde5b60828ac7f8b6c2addaf220b    = I6f8f253cfb1fe1c2254e557f732a9b22;

            I0f644f42cabf871b71e5a82871bc7b5d = Id36e8953a02400a5ab1f4dfdb0422e6d + ~I3da241c7f221413abfbf1b4384bfca5a + 1;
            I3f247e74edd47e346d3bbb5dc3408844 = I2bcab411f9bec1541259751bcb9e0823(I0f644f42cabf871b71e5a82871bc7b5d);
            I150c28296847348d69cce123f20656c3    = I3f247e74edd47e346d3bbb5dc3408844;

            I71f9e059726a6cac8bdf0efcc0eadd2b = Ica71108a53bfcfd1892b4d03ef68110c + ~I8c5f98353b5b082dc3cf056469945a08 + 1;
            Ie0b33e2c1def11ccdaaae4ed2b042df6 = I2bcab411f9bec1541259751bcb9e0823(I71f9e059726a6cac8bdf0efcc0eadd2b);
            Ib94d38d19b3791fa2d1b42fdfde8435e    = Ie0b33e2c1def11ccdaaae4ed2b042df6;

            I0c9b2c1da30bfab514bbb556ae7bd4c4 = Ica71108a53bfcfd1892b4d03ef68110c + ~If8865fee7dbf593b34ea54692d947f10 + 1;
            I39448514454c92ce93c3b0bc1d0e5d50 = I2bcab411f9bec1541259751bcb9e0823(I0c9b2c1da30bfab514bbb556ae7bd4c4);
            I94865622898b2e481e86a244f7aa2759    = I39448514454c92ce93c3b0bc1d0e5d50;

            I7918b2e37e96aee94fbccca7e0f75fc4 = Ica71108a53bfcfd1892b4d03ef68110c + ~Ib5334df42ee8f1574e41cb30b903fae9 + 1;
            I677e9047c3ede581db9512b4fe072ea9 = I2bcab411f9bec1541259751bcb9e0823(I7918b2e37e96aee94fbccca7e0f75fc4);
            I1a4a432e735367f515ca747cef7d7d04    = I677e9047c3ede581db9512b4fe072ea9;

            I76eebd77eb77e0abcbc727d2c511370a = Ica71108a53bfcfd1892b4d03ef68110c + ~Icbc12ab47f586b12402ae5d4361c967d + 1;
            Ief6fbe6927f26b7a037f8e0bcb7751d8 = I2bcab411f9bec1541259751bcb9e0823(I76eebd77eb77e0abcbc727d2c511370a);
            Ib3a2b744d8f38671a63da6f8f8f1a6a1    = Ief6fbe6927f26b7a037f8e0bcb7751d8;

            Ibb2288e62110bae5b2d3fe901974e5c7 = Ica71108a53bfcfd1892b4d03ef68110c + ~Ie8644d7edbadf19937c399cf275946e5 + 1;
            Ie1e5c12afad8f2d8c2abef26473b7d9c = I2bcab411f9bec1541259751bcb9e0823(Ibb2288e62110bae5b2d3fe901974e5c7);
            I87716ad5a64592abb812ffe041ccc163    = Ie1e5c12afad8f2d8c2abef26473b7d9c;

            I080f931dfef9d8adfb1dc1ee073eb64c = Ica71108a53bfcfd1892b4d03ef68110c + ~I2087576fbc15119bf5d9e8afa2603b69 + 1;
            Ic8f2ae80147ee27c548de195dfefa382 = I2bcab411f9bec1541259751bcb9e0823(I080f931dfef9d8adfb1dc1ee073eb64c);
            I71b259faefbea7ce8f47e0ffb556a0be    = Ic8f2ae80147ee27c548de195dfefa382;

            Ide1106431e3565158bd81ccd6b18f3a1 = Ica71108a53bfcfd1892b4d03ef68110c + ~If1ec4241fd12255369f72b3f3310b6e7 + 1;
            I533eb0729cc85339e2fcd1847930adc9 = I2bcab411f9bec1541259751bcb9e0823(Ide1106431e3565158bd81ccd6b18f3a1);
            I2161b2ff3514dbdbb79d25da87eeec2b    = I533eb0729cc85339e2fcd1847930adc9;

            I63df19931e8d28666cccd79922cbd418 = Ica71108a53bfcfd1892b4d03ef68110c + ~I401ab1ad994f5018061a3f57d3a51ad1 + 1;
            Ic68fd0a9ea4b641913aadb7fe011d8ab = I2bcab411f9bec1541259751bcb9e0823(I63df19931e8d28666cccd79922cbd418);
            I860a3c9fca8d240c68ce3825192353b0    = Ic68fd0a9ea4b641913aadb7fe011d8ab;

            I9a7e4a59447048de90446f877eb06627 = Ica71108a53bfcfd1892b4d03ef68110c + ~I2ba16a10a82c20d54c776a9804ee50e4 + 1;
            Ica1f13759a67176573842e56bcdf09bd = I2bcab411f9bec1541259751bcb9e0823(I9a7e4a59447048de90446f877eb06627);
            Ie4eb18c7e906c9a25c12e9980a9f61cb    = Ica1f13759a67176573842e56bcdf09bd;

            I0917e92ed84363ca92fd2074acd74eba = Ica71108a53bfcfd1892b4d03ef68110c + ~Ib55b0e4c45ebbdb605f0ba9d62bff21c + 1;
            Ifed30886099cbeb5da64d1d0696bb5de = I2bcab411f9bec1541259751bcb9e0823(I0917e92ed84363ca92fd2074acd74eba);
            I20a24846a74af76fa4470d6350546a9a    = Ifed30886099cbeb5da64d1d0696bb5de;

            Ie3eefdf7b5561a90a6ddd9e6aa432509 = I7c97629ec6e594f9b2160815ddd133cc + ~Id8c36004ae8e550569a491f6b514945a + 1;
            I317b34a0f6e16550b4a3e887cdd0c250 = I2bcab411f9bec1541259751bcb9e0823(Ie3eefdf7b5561a90a6ddd9e6aa432509);
            I90d40f6e9721a7d075512b8b81907453    = I317b34a0f6e16550b4a3e887cdd0c250;

            I56eeb10d11e886cff629457a640a1c76 = I7c97629ec6e594f9b2160815ddd133cc + ~I840a1a7c0bf49f4f42499b33f32fa02d + 1;
            I39fa2bacef89a2f523f91b1e7f3cbe90 = I2bcab411f9bec1541259751bcb9e0823(I56eeb10d11e886cff629457a640a1c76);
            Ifc4525a25f38affb399004b057d1318c    = I39fa2bacef89a2f523f91b1e7f3cbe90;

            I7a9eea89c4e76d856df44b6bdc332840 = I7c97629ec6e594f9b2160815ddd133cc + ~Id769d4a92f5f6da262ce0521e5509368 + 1;
            Id01272140c18ae29a8c75e493cf01268 = I2bcab411f9bec1541259751bcb9e0823(I7a9eea89c4e76d856df44b6bdc332840);
            Icc93649a2050b9ded1e625be936b411f    = Id01272140c18ae29a8c75e493cf01268;

            If8d8f4333e893788fcb9ec54256e5b7a = I7c97629ec6e594f9b2160815ddd133cc + ~I19875f52f79482b477f1febaa7e97090 + 1;
            I4d981fbbadbaa97ef98429ac12ca6710 = I2bcab411f9bec1541259751bcb9e0823(If8d8f4333e893788fcb9ec54256e5b7a);
            Ibcc30c960ae0f29c4efb1266c9e490ac    = I4d981fbbadbaa97ef98429ac12ca6710;

            Ie4af0e7e04778d85f5dee73da33376a8 = I7c97629ec6e594f9b2160815ddd133cc + ~I3f2507530dd648814af0964f7da11d35 + 1;
            I2a1672224d3a3c513f2f04bb4dc123e0 = I2bcab411f9bec1541259751bcb9e0823(Ie4af0e7e04778d85f5dee73da33376a8);
            I3b2ffa79fd2227a24c6468a89f2bd989    = I2a1672224d3a3c513f2f04bb4dc123e0;

            I019a4e997adf54f5f5ca651f80b7901b = I7c97629ec6e594f9b2160815ddd133cc + ~I8b5d10c412daccdcb07645bf239d61bd + 1;
            I364afb3546858e133a2bb541798e7886 = I2bcab411f9bec1541259751bcb9e0823(I019a4e997adf54f5f5ca651f80b7901b);
            Ib489a11dfdd8a2b3ad561c965b3d7d2a    = I364afb3546858e133a2bb541798e7886;

            I10294667f09abbfd4e2f757c414072fc = I7c97629ec6e594f9b2160815ddd133cc + ~I3a09554ca009781e28ef1b3ea70d39ad + 1;
            I9908671d65856b8714d43d83f0811a17 = I2bcab411f9bec1541259751bcb9e0823(I10294667f09abbfd4e2f757c414072fc);
            Ifa51cf9f9d3d1b91c72387f5daf05c79    = I9908671d65856b8714d43d83f0811a17;

            Id4e8ab8f15b36bd27d1e4ebc5cbe1495 = I7c97629ec6e594f9b2160815ddd133cc + ~I37e5c3118e8536e37bd797aeaa92476c + 1;
            I3e3f06cade9b6c8ea10e45996449e405 = I2bcab411f9bec1541259751bcb9e0823(Id4e8ab8f15b36bd27d1e4ebc5cbe1495);
            Ifda20d77c574c8f13816620c56fff950    = I3e3f06cade9b6c8ea10e45996449e405;

            I6c93588ca9e7c623d75314da39e89a91 = I7c97629ec6e594f9b2160815ddd133cc + ~Ifbcebda2bb0ce58a0e1764c392a816df + 1;
            I9525b42d4dc80c42608cfa0ea10b8b2d = I2bcab411f9bec1541259751bcb9e0823(I6c93588ca9e7c623d75314da39e89a91);
            I03ce0915d3a170429959221b6c8cd16c    = I9525b42d4dc80c42608cfa0ea10b8b2d;

            I1020412efc78d12a9ebcbaeb83e5dcea = I7c97629ec6e594f9b2160815ddd133cc + ~Iaed105b99eae5b078521e3a94d8a79b7 + 1;
            I94361c7eb9f16c4b20dfcdb7b8ad8cf3 = I2bcab411f9bec1541259751bcb9e0823(I1020412efc78d12a9ebcbaeb83e5dcea);
            I9c2da511df8277b7e61cf8611d04dd32    = I94361c7eb9f16c4b20dfcdb7b8ad8cf3;

            Id0b574f35a83dcfd4481a10043cd1884 = I4823c8239ace86dc399e906c1b5a0d74 + ~I2a2d014f94d7a3b9fb3024a3e9107a73 + 1;
            Idc043493a919ec50417594df96f4d669 = I2bcab411f9bec1541259751bcb9e0823(Id0b574f35a83dcfd4481a10043cd1884);
            Ib8c628f3d97ffdf8a8b5db0fe90bbfa8    = Idc043493a919ec50417594df96f4d669;

            Ifc577e5c2c7288373a8c5e3969ac1589 = I4823c8239ace86dc399e906c1b5a0d74 + ~I9aa11f30712f1779339b985212a7979c + 1;
            I9e051ecfe79c36a913b15a0c7fe27f4d = I2bcab411f9bec1541259751bcb9e0823(Ifc577e5c2c7288373a8c5e3969ac1589);
            I42e0e42ae26723497a1da5e86e855499    = I9e051ecfe79c36a913b15a0c7fe27f4d;

            Id18a1a17c1cf6e8a2492aa73b62898f2 = I4823c8239ace86dc399e906c1b5a0d74 + ~Id15c3bdce785df234c68432ccec8f959 + 1;
            I5479857f4f724aaea25ba124c9edb232 = I2bcab411f9bec1541259751bcb9e0823(Id18a1a17c1cf6e8a2492aa73b62898f2);
            Id7e44a94fcaa2ca22ac9eb6756ecb830    = I5479857f4f724aaea25ba124c9edb232;

            Id8ce8f636723b9f119bb86c25017e6b3 = I4823c8239ace86dc399e906c1b5a0d74 + ~Ia0e77e9544481aa0f56dfdb6eb253137 + 1;
            Id2ed64cae3cb1e0ada8e3fb4ebb2dc78 = I2bcab411f9bec1541259751bcb9e0823(Id8ce8f636723b9f119bb86c25017e6b3);
            Ie91db5e628b828dfaa8c1bd7d614d986    = Id2ed64cae3cb1e0ada8e3fb4ebb2dc78;

            Ic29a18d8d504a2d5280c1d7771346518 = I10ad572ca72c2ea991487c39f7eabd7b + ~Ia4b2db3d48f946b0bfd0be0e32d7518d + 1;
            I16b9849d3f2edd7f9ed7accb138d2c02 = I2bcab411f9bec1541259751bcb9e0823(Ic29a18d8d504a2d5280c1d7771346518);
            I683ebfd7677d9e175d7a86479a5b42c6    = I16b9849d3f2edd7f9ed7accb138d2c02;

            I96a79193aa2956b8f901d5fcc9cf65cf = I10ad572ca72c2ea991487c39f7eabd7b + ~I111ac0aadbdd3e4479ca0786491a7b08 + 1;
            Ibcfe38455aa7aa33ae950172fb915dc5 = I2bcab411f9bec1541259751bcb9e0823(I96a79193aa2956b8f901d5fcc9cf65cf);
            I11090ba16ce17a70438618b474837c33    = Ibcfe38455aa7aa33ae950172fb915dc5;

            I8c97a246c749fbef029f8b1671c772bd = I10ad572ca72c2ea991487c39f7eabd7b + ~I7caf8c7496dd96c1ed08e98b415f5775 + 1;
            Ic9d9832294a3707b4041b2c4d8f92615 = I2bcab411f9bec1541259751bcb9e0823(I8c97a246c749fbef029f8b1671c772bd);
            I845dd61995152e9d39cea7f0370b5a4d    = Ic9d9832294a3707b4041b2c4d8f92615;

            If9ba9d221909ce7499725f6fd7d519f8 = I10ad572ca72c2ea991487c39f7eabd7b + ~Iec0d7ea31e0f1a75b15121090dcf1e11 + 1;
            I3ef9641c53e7aa6a588481b57b865aa3 = I2bcab411f9bec1541259751bcb9e0823(If9ba9d221909ce7499725f6fd7d519f8);
            Ia3e4dff8c98b38b6aebec9094ed26421    = I3ef9641c53e7aa6a588481b57b865aa3;

            I53a7878f44253f0f1a82d9d27b1a44c3 = Ie9f3fd3a6d16316e55addbe0e336519f + ~Icc5d7bcbd7fcdb5092e6d8e18f6de6ec + 1;
            Ie838f76c6fc041e4fa66441094ae477c = I2bcab411f9bec1541259751bcb9e0823(I53a7878f44253f0f1a82d9d27b1a44c3);
            Id69a54dc4854348a482f052c64a736ca    = Ie838f76c6fc041e4fa66441094ae477c;

            Ie0e928125f9d3d17d123d97e00f1fc34 = Ie9f3fd3a6d16316e55addbe0e336519f + ~I27951ef3d612004abdc639662807426b + 1;
            Ice9f8149ed08f537da5e146b417085e0 = I2bcab411f9bec1541259751bcb9e0823(Ie0e928125f9d3d17d123d97e00f1fc34);
            I0f56c52253603ac01a22f3b942429262    = Ice9f8149ed08f537da5e146b417085e0;

            I2bd0f77efeca09eebe82ea234e9fe638 = Ie9f3fd3a6d16316e55addbe0e336519f + ~I6c9ae8b8191507f908c27bbde53bf2d5 + 1;
            I71f6bd2fe34731aab306cfb89a3335ca = I2bcab411f9bec1541259751bcb9e0823(I2bd0f77efeca09eebe82ea234e9fe638);
            I718f82404f82fe0e822ee20d33ad20a2    = I71f6bd2fe34731aab306cfb89a3335ca;

            I94f2e7ef9b3463bd598dc9049f6fb0ef = Ie9f3fd3a6d16316e55addbe0e336519f + ~Ia98bb3648ce3719b1c31ce0f41121c63 + 1;
            I5dd57cfd0d7ce83fcbdb3f560ac713fb = I2bcab411f9bec1541259751bcb9e0823(I94f2e7ef9b3463bd598dc9049f6fb0ef);
            I6c86073aaa32b64a43d06eb1a2d9fba8    = I5dd57cfd0d7ce83fcbdb3f560ac713fb;

            I6dc16510af6b61b79b339d0fce77ac24 = I07965bca84276dd56da1af98e64b0adc + ~I5e0d6b44474a226ab2ce916a6d46072a + 1;
            I239498228bdcb1c2a8b2cbef48e850a6 = I2bcab411f9bec1541259751bcb9e0823(I6dc16510af6b61b79b339d0fce77ac24);
            Ie0c8e27167e6ba97a83dd238086f45e6    = I239498228bdcb1c2a8b2cbef48e850a6;

            Ic655e213ab81f5d61a018d3ed7016b12 = I07965bca84276dd56da1af98e64b0adc + ~I9068cca0de6ecff56ca542d0998fcab2 + 1;
            I82fc4233a3d2840670eb9b9adf6c9215 = I2bcab411f9bec1541259751bcb9e0823(Ic655e213ab81f5d61a018d3ed7016b12);
            I6bb5e8ee16a2bc0c3b77c882cfb659e7    = I82fc4233a3d2840670eb9b9adf6c9215;

            I2ffc4a604025a2f5c4e273c1d070a725 = I07965bca84276dd56da1af98e64b0adc + ~I9cab38b69794ab661e12750cf69c822c + 1;
            Ieb08f6a94aa827632606608d014e26d3 = I2bcab411f9bec1541259751bcb9e0823(I2ffc4a604025a2f5c4e273c1d070a725);
            Ieef625ad664ddadc849be46d1c083748    = Ieb08f6a94aa827632606608d014e26d3;

            I1c76818a9a3b688ca897aa479f7d807f = I07965bca84276dd56da1af98e64b0adc + ~Id9c8055ef530f2cb8096cb7bb2af55a4 + 1;
            Ifdbb9947713ac574738236fcb5c6ae07 = I2bcab411f9bec1541259751bcb9e0823(I1c76818a9a3b688ca897aa479f7d807f);
            Ice91b069200a91b2ad48fbf87bb2e766    = Ifdbb9947713ac574738236fcb5c6ae07;

            I3bfee9d3d88f0569010a4e0101200c19 = Ic2ade31b8bcf68c4dcc1a371ff14074b + ~I5bab5ae46114c487f67b8e779d7461df + 1;
            Ia737ee8f2c01feba1db87fe3e1a2388c = I2bcab411f9bec1541259751bcb9e0823(I3bfee9d3d88f0569010a4e0101200c19);
            I9d4c7c85b4da5f7003ff05ed3a240a2e    = Ia737ee8f2c01feba1db87fe3e1a2388c;

            I5d4738755a26beb6d0f61dd3dec0f804 = Ic2ade31b8bcf68c4dcc1a371ff14074b + ~Ib3ec015a3d43d46e0b7142b21a81cfee + 1;
            I5d8e065dba640832d9d8db3e4338fbb5 = I2bcab411f9bec1541259751bcb9e0823(I5d4738755a26beb6d0f61dd3dec0f804);
            Ia8f1616f8a65025446a5ab4cc1624f9b    = I5d8e065dba640832d9d8db3e4338fbb5;

            I2f3c800091275bcb72d1a2a38fba53f3 = Ic2ade31b8bcf68c4dcc1a371ff14074b + ~Iee0e45914c52a357e1e32922299d6937 + 1;
            I3b3e36ffb1cff2c07bc9a61afdde10c1 = I2bcab411f9bec1541259751bcb9e0823(I2f3c800091275bcb72d1a2a38fba53f3);
            I29848deb21ad480cdf155d849dc7bd48    = I3b3e36ffb1cff2c07bc9a61afdde10c1;

            I378e67cca7c4ff6325683f8346963210 = Ic2ade31b8bcf68c4dcc1a371ff14074b + ~I1684820afb9d9cec38cfdfcd6ca8b36a + 1;
            I2c8137e5ee04a1067858d7bb8d09d65b = I2bcab411f9bec1541259751bcb9e0823(I378e67cca7c4ff6325683f8346963210);
            I1ae69988f89b200bd0e48f640211321c    = I2c8137e5ee04a1067858d7bb8d09d65b;

            I04c8915a7f4bbde003f7facc84435c1a = Ic2ade31b8bcf68c4dcc1a371ff14074b + ~I25888aa2135fc403ca9eac4df634549a + 1;
            I38eb22d29ad9f4192499980fc17898b4 = I2bcab411f9bec1541259751bcb9e0823(I04c8915a7f4bbde003f7facc84435c1a);
            I7ddcc3c9f4d21aacc07d8eb285dee83e    = I38eb22d29ad9f4192499980fc17898b4;

            I3f50b10072f38b6addee6845e6df9118 = Ic2ade31b8bcf68c4dcc1a371ff14074b + ~Ib9081d438413a627f5b16f68c2eabb80 + 1;
            Ib714941df0aaca40e7573e030d97b3f1 = I2bcab411f9bec1541259751bcb9e0823(I3f50b10072f38b6addee6845e6df9118);
            I28f7cf50ea7ac81667ff1353e0e121bd    = Ib714941df0aaca40e7573e030d97b3f1;

            Icc60eb18ba740036d2a17f98f15cfb98 = Ic0edcf240048fbfde4e938c3e4c5e281 + ~I4d908bbe633c193cd9fc93dd33c60bd2 + 1;
            I47bcab5b082a8ce6312244224c162d39 = I2bcab411f9bec1541259751bcb9e0823(Icc60eb18ba740036d2a17f98f15cfb98);
            I09b7dd699ae0c4d34a7d1588efc90452    = I47bcab5b082a8ce6312244224c162d39;

            I1677daa18aa8b226753b1a887b9420d1 = Ic0edcf240048fbfde4e938c3e4c5e281 + ~I65928407b1d5447dbc815cd2d2e7b37d + 1;
            I68ded74f52dbd02ceb1da62a79d619d2 = I2bcab411f9bec1541259751bcb9e0823(I1677daa18aa8b226753b1a887b9420d1);
            Ic937101cc53e67403e56ac85011aa9ba    = I68ded74f52dbd02ceb1da62a79d619d2;

            I36bc2d4c9a4480daa9b0944c08b50738 = Ic0edcf240048fbfde4e938c3e4c5e281 + ~Ic7855ca956651bd368cbdde7ec93ba6d + 1;
            Iaa113fd5f1e0c51d9f47240fe81b5604 = I2bcab411f9bec1541259751bcb9e0823(I36bc2d4c9a4480daa9b0944c08b50738);
            Ib42b03d2f76b8939ff3183008b17a969    = Iaa113fd5f1e0c51d9f47240fe81b5604;

            I38419a6905f50135a6783aacca0384dd = Ic0edcf240048fbfde4e938c3e4c5e281 + ~I7a6ab9e700bd94208ab6528af413f3a9 + 1;
            I907bf413f65fad54303751c054687b29 = I2bcab411f9bec1541259751bcb9e0823(I38419a6905f50135a6783aacca0384dd);
            I4b99f00b1c2cdcee6bf4f1d2e8199ee4    = I907bf413f65fad54303751c054687b29;

            Ib48892dcb0715987289662a14672611e = Ic0edcf240048fbfde4e938c3e4c5e281 + ~I7fc6e2aecff5bd691872d1e10a39103b + 1;
            I7b727f2e9454f90d4fa4ef2cf69ddf23 = I2bcab411f9bec1541259751bcb9e0823(Ib48892dcb0715987289662a14672611e);
            I01e153b020e1349eb66b47de581408df    = I7b727f2e9454f90d4fa4ef2cf69ddf23;

            Icd9c94f929dbc71c9b836fda3019630b = Ic0edcf240048fbfde4e938c3e4c5e281 + ~I9c5bf5451736358f8c84e150004fa5a9 + 1;
            I6fc1f37134064dd7514b46ce7d27ceaa = I2bcab411f9bec1541259751bcb9e0823(Icd9c94f929dbc71c9b836fda3019630b);
            I8ca1a48206ed8f1dc7ca57d77d0331a2    = I6fc1f37134064dd7514b46ce7d27ceaa;

            I5d0249d9a772805b3fba3f3c7f5d35bd = I8b42e89ff5f780d4ef8cd1cd5c99ef61 + ~I83cec264bd378f1dc23f87e439e7310e + 1;
            I7856585e0374651fc5f9921f69706a0b = I2bcab411f9bec1541259751bcb9e0823(I5d0249d9a772805b3fba3f3c7f5d35bd);
            I40e8430f50206db37e500c22f461b0c7    = I7856585e0374651fc5f9921f69706a0b;

            Ie97341deb6fb24d49eb8b96bd0fd3f35 = I8b42e89ff5f780d4ef8cd1cd5c99ef61 + ~Ib83242b57ab050b0e5f9bdf91fa118fb + 1;
            I79b1967c2128c611ee4fe0d14bced1f4 = I2bcab411f9bec1541259751bcb9e0823(Ie97341deb6fb24d49eb8b96bd0fd3f35);
            I521128b7d945e025ded04037494c850a    = I79b1967c2128c611ee4fe0d14bced1f4;

            I17dd788f9d8e91307b6b1ab7488f9ce2 = I8b42e89ff5f780d4ef8cd1cd5c99ef61 + ~I8ab7efc436a0f2cc3efbc299a0ddf914 + 1;
            Ib8aeaf62789d1d7a5a23d7492ff551b2 = I2bcab411f9bec1541259751bcb9e0823(I17dd788f9d8e91307b6b1ab7488f9ce2);
            Ic24dbb1a30bb9a32c1992afcba90d4fb    = Ib8aeaf62789d1d7a5a23d7492ff551b2;

            I92ae370022ed107b152b10fd0aa3d2b7 = I8b42e89ff5f780d4ef8cd1cd5c99ef61 + ~I9b1390839ee2b9ba591e3873e967c8e2 + 1;
            I9a8e8c3ce2c6323acee0877d445a2268 = I2bcab411f9bec1541259751bcb9e0823(I92ae370022ed107b152b10fd0aa3d2b7);
            I06cc903106b42e397fa7c4bc6c5edea4    = I9a8e8c3ce2c6323acee0877d445a2268;

            Iebb39f0d19ec1208bbfba6cf67a3bfc7 = I8b42e89ff5f780d4ef8cd1cd5c99ef61 + ~Iec936eeebd1f8c95307bd8705e6def81 + 1;
            I701a3c05ad8e6ac5cea30b78707e77d1 = I2bcab411f9bec1541259751bcb9e0823(Iebb39f0d19ec1208bbfba6cf67a3bfc7);
            I765dff22de01d419a6626919d23850f2    = I701a3c05ad8e6ac5cea30b78707e77d1;

            I81861f6bb8bbbab6e93407cfb4a852b8 = I8b42e89ff5f780d4ef8cd1cd5c99ef61 + ~I377933518c3807edb71f648c65ad5c85 + 1;
            I75fefd09122859510021931c16051262 = I2bcab411f9bec1541259751bcb9e0823(I81861f6bb8bbbab6e93407cfb4a852b8);
            Ie9538b63a057a50371de2d17898d3ad7    = I75fefd09122859510021931c16051262;

            I217b2e3ca0a534fc5b1910adf3c1b57d = I70b1b8521b36920707e95fc9418eb8a9 + ~I0c53d8d6a5b92960e29fc31cf456c23b + 1;
            I2779af0ff280ea511af850df795d1fb6 = I2bcab411f9bec1541259751bcb9e0823(I217b2e3ca0a534fc5b1910adf3c1b57d);
            If93a5596528db9017b8783fa0cf1dbc2    = I2779af0ff280ea511af850df795d1fb6;

            I8429b08891dc56af24c72ce1b7725457 = I70b1b8521b36920707e95fc9418eb8a9 + ~Ice4f4ba8bb3381c8846941d5d5fe4534 + 1;
            I2eb84b0b6b12b9269bb791ae03e5094d = I2bcab411f9bec1541259751bcb9e0823(I8429b08891dc56af24c72ce1b7725457);
            I68016caaf170fbe2734c5b6aaf089894    = I2eb84b0b6b12b9269bb791ae03e5094d;

            If96747262303f6c5c6b129e39224bd23 = I70b1b8521b36920707e95fc9418eb8a9 + ~I2b0b168ce4fe8aa4a2e7cb69fe532aa3 + 1;
            Ie42cb87efb2b87d88eed6139132bb23e = I2bcab411f9bec1541259751bcb9e0823(If96747262303f6c5c6b129e39224bd23);
            I169b0fac6d01a713986b636bf8dfc3fb    = Ie42cb87efb2b87d88eed6139132bb23e;

            If7012457af15c405baeaa1710319b541 = I70b1b8521b36920707e95fc9418eb8a9 + ~I2e14fb1e667e967ab4c116e0c7438aec + 1;
            Id2e2722999e300df1bc7ea89dbf5689d = I2bcab411f9bec1541259751bcb9e0823(If7012457af15c405baeaa1710319b541);
            Iddb14d68b464d04fe9e0b4e62789601a    = Id2e2722999e300df1bc7ea89dbf5689d;

            Ia0a0229ef71b85195352bb664ea4e4e3 = I70b1b8521b36920707e95fc9418eb8a9 + ~I24180fba17c21bacefa8a4514e4b685c + 1;
            I2b7e1a65c52821f3f7e194a443b0117d = I2bcab411f9bec1541259751bcb9e0823(Ia0a0229ef71b85195352bb664ea4e4e3);
            Ie5b71f77beb734a6ab7f7be6c6f9c252    = I2b7e1a65c52821f3f7e194a443b0117d;

            I42aeb7c23accc2ca874c7f8221c3af93 = I70b1b8521b36920707e95fc9418eb8a9 + ~Icec98d794a64752081fadfa74308fad3 + 1;
            I8b31aa4edbc800c99628c5851cad8770 = I2bcab411f9bec1541259751bcb9e0823(I42aeb7c23accc2ca874c7f8221c3af93);
            I59f9fa0b81ca88915c338ece1d1e08d5    = I8b31aa4edbc800c99628c5851cad8770;

            I7df6a95bf51f40693c439c6df36510d4 = I4fb1c32a62cbbaeb585c6564a3c938f9 + ~I45373bff54eccf8137da2931d841934e + 1;
            Id40d461c28ecc2017d9b7d2eadf5ea44 = I2bcab411f9bec1541259751bcb9e0823(I7df6a95bf51f40693c439c6df36510d4);
            I4f27922ccb21b65dcfe2dc0fcc97cdf3    = Id40d461c28ecc2017d9b7d2eadf5ea44;

            I8fe65f9c344d7ec8657f192abefc3fb6 = I4fb1c32a62cbbaeb585c6564a3c938f9 + ~I3934ed7170967ff3852944cc39ba1de9 + 1;
            I4b8f58440e6848610f2e7e06efbc64fe = I2bcab411f9bec1541259751bcb9e0823(I8fe65f9c344d7ec8657f192abefc3fb6);
            Idd7ae55ba748fb36e49684037212936d    = I4b8f58440e6848610f2e7e06efbc64fe;

            I4d75c95d34d8d8aeeb528456bbe136e1 = I4fb1c32a62cbbaeb585c6564a3c938f9 + ~I17e818b67440efaba9a5d19e7467bf85 + 1;
            Ica1d5cc8dc277e91787ec1bf0f2ed65c = I2bcab411f9bec1541259751bcb9e0823(I4d75c95d34d8d8aeeb528456bbe136e1);
            Ib8da505d1572487e814e7b0682e6dfa9    = Ica1d5cc8dc277e91787ec1bf0f2ed65c;

            I43746054a38c9521f8da9db9d0e91f99 = I4fb1c32a62cbbaeb585c6564a3c938f9 + ~Ia5b779ef95333736b08f63770900e275 + 1;
            Ie5d481ac7a371e1fd3c48c5cf9649a67 = I2bcab411f9bec1541259751bcb9e0823(I43746054a38c9521f8da9db9d0e91f99);
            Idedb59a6fa2f6ad049f81ac652c645d8    = Ie5d481ac7a371e1fd3c48c5cf9649a67;

            I0430ac2a4b2b2e2fc7f8154bf946553c = I4fb1c32a62cbbaeb585c6564a3c938f9 + ~I83bbe6fa947f9f909e1a6785ab31901f + 1;
            I9786bf468ba8540d7e75d762fc832709 = I2bcab411f9bec1541259751bcb9e0823(I0430ac2a4b2b2e2fc7f8154bf946553c);
            I7d50b49718ab2007accda67ac77a65d0    = I9786bf468ba8540d7e75d762fc832709;

            I25dc807fd55b81c9f24fd0d1edcaa758 = I4fb1c32a62cbbaeb585c6564a3c938f9 + ~I7bbe4d0a7d61d3f7da346de71b9a3a5f + 1;
            Ib093fabefab0a1b46d2199c1c948abc8 = I2bcab411f9bec1541259751bcb9e0823(I25dc807fd55b81c9f24fd0d1edcaa758);
            I27e0600689451a7475a36143f0eb1079    = Ib093fabefab0a1b46d2199c1c948abc8;

            I7881184f1779b9fd4fdf329c5f7664da = Iefc37daeec14e14ef2fe0716f73109dc + ~Ib14733d3585dbf7f196cfc068e9508f0 + 1;
            I9b53bbb22003297175c6c4655ef83c93 = I2bcab411f9bec1541259751bcb9e0823(I7881184f1779b9fd4fdf329c5f7664da);
            Iba6724b61ecb74552b9bb3cab96480c6    = I9b53bbb22003297175c6c4655ef83c93;

            I8e6de2d692a307ee8a5a4b2a9265a633 = Iefc37daeec14e14ef2fe0716f73109dc + ~I3e8d26ea83937cae01aadf1092c59bdf + 1;
            I9df2a441fadba7dc49effc5eecf4b0e8 = I2bcab411f9bec1541259751bcb9e0823(I8e6de2d692a307ee8a5a4b2a9265a633);
            I0abb44bd896fbc695e880fee67fb0c42    = I9df2a441fadba7dc49effc5eecf4b0e8;

            I54b2b18ab051b468808a3d0fc4bc893f = Iefc37daeec14e14ef2fe0716f73109dc + ~I0fb60c4f56f6d7b4007cf0dae39f4573 + 1;
            I102372ac8a06119e5d827d83f172bbd2 = I2bcab411f9bec1541259751bcb9e0823(I54b2b18ab051b468808a3d0fc4bc893f);
            Ifd714548110aa979e735cc6e13d3ef57    = I102372ac8a06119e5d827d83f172bbd2;

            I37ee86e2ca32832862cb57efe76bbedf = Iefc37daeec14e14ef2fe0716f73109dc + ~If3bdbb4c20efca0c5af78614b4271ed1 + 1;
            I5cad4cd564b0956b08f22cd42d594b01 = I2bcab411f9bec1541259751bcb9e0823(I37ee86e2ca32832862cb57efe76bbedf);
            Ieeb6c7cdf1379ee3d2933d81bc812dbc    = I5cad4cd564b0956b08f22cd42d594b01;

            Ic95f2fc697574803c0f7fa35c2609f0c = Iefc37daeec14e14ef2fe0716f73109dc + ~I632ffd09a9091335b3aa91ab2a8f1cce + 1;
            Id685ced1c37d97c75b49b2f790dbabad = I2bcab411f9bec1541259751bcb9e0823(Ic95f2fc697574803c0f7fa35c2609f0c);
            Id682af5250edce8e3811d418ecf2dd10    = Id685ced1c37d97c75b49b2f790dbabad;

            I933a30c52c9bec5172530b2d739a3b63 = Iefc37daeec14e14ef2fe0716f73109dc + ~I197c05f74bf7fb8d44124d40bd7c6563 + 1;
            I219e400c87948e7b2bf715745a4b152c = I2bcab411f9bec1541259751bcb9e0823(I933a30c52c9bec5172530b2d739a3b63);
            I1d02127e28fb2e9aaf352815627960e7    = I219e400c87948e7b2bf715745a4b152c;

            I7bbd7df18f85197c22fe8cfe37312af6 = Ibd15f164f6d2ac9e5721a21464bc2c5c + ~Ied7e494fb288f78d110ed06662f1926a + 1;
            I3372567dacc350adf991928753209605 = I2bcab411f9bec1541259751bcb9e0823(I7bbd7df18f85197c22fe8cfe37312af6);
            Ibee34260749dc92b8523e83cd64d6a40    = I3372567dacc350adf991928753209605;

            I50d5ada7c91c7af16492c6b41151b68f = Ibd15f164f6d2ac9e5721a21464bc2c5c + ~Iefe423653d454e21324a6857b52f98ac + 1;
            Ibf50476ac553bceaedcb121b28093394 = I2bcab411f9bec1541259751bcb9e0823(I50d5ada7c91c7af16492c6b41151b68f);
            Ie9a2a59c7b3571194198dca0c679c5f6    = Ibf50476ac553bceaedcb121b28093394;

            I32c8e7996b3473d4906c40018799a16b = Ibd15f164f6d2ac9e5721a21464bc2c5c + ~Ice8a82bdd966719098a8d5f2a826f73d + 1;
            I5d20fcccde5844e36b83d7fd7034c413 = I2bcab411f9bec1541259751bcb9e0823(I32c8e7996b3473d4906c40018799a16b);
            Ie4b5a941feb385e88498a98e5f8ddc01    = I5d20fcccde5844e36b83d7fd7034c413;

            Ic0eacd5a4812ad7ae3fa251ab2db4694 = Ibd15f164f6d2ac9e5721a21464bc2c5c + ~I3a47540f34ce47bcfa1da66cc4e6e088 + 1;
            I47e720341773b3a11f4c71b4e9644525 = I2bcab411f9bec1541259751bcb9e0823(Ic0eacd5a4812ad7ae3fa251ab2db4694);
            I30b2b34a0cecfdbdeecba5f286befccd    = I47e720341773b3a11f4c71b4e9644525;

            Ideecf8ab87d28a840cd93851169ab05b = Ibd15f164f6d2ac9e5721a21464bc2c5c + ~I49321308413cb4dbe5e6c01ba5b9023c + 1;
            I0251d8ecec82a24878ce494f0b417ce3 = I2bcab411f9bec1541259751bcb9e0823(Ideecf8ab87d28a840cd93851169ab05b);
            I8ce739ddc344cacb2de7f2c88a882170    = I0251d8ecec82a24878ce494f0b417ce3;

            I1ac6775eb38457b7962241d2e7336b0d = Ibd15f164f6d2ac9e5721a21464bc2c5c + ~I92acc55d81ec6e02880337b0a451ae21 + 1;
            Ibeef795b2235c98439628da8d7c094e0 = I2bcab411f9bec1541259751bcb9e0823(I1ac6775eb38457b7962241d2e7336b0d);
            I8b00260bb93e928e66e9d4aaeb0d9b55    = Ibeef795b2235c98439628da8d7c094e0;

            I2ecaa89698604fddd863d7e28d643a57 = I951dfff9507bb70214d48e03a0ebb3a7 + ~Ib16c6096ce80e2f15a5ccea145e28510 + 1;
            I61769f7c08a0b9cf78068455410b6bb2 = I2bcab411f9bec1541259751bcb9e0823(I2ecaa89698604fddd863d7e28d643a57);
            I9c1ca916654bad308af37d040b486cf8    = I61769f7c08a0b9cf78068455410b6bb2;

            I273e0fe9c51c8549c8dfff393ca2e4e1 = I951dfff9507bb70214d48e03a0ebb3a7 + ~Ic57a2627a194099105a2908a41feddfb + 1;
            I77fe52c685b1075c294ac3c0a5b0d63a = I2bcab411f9bec1541259751bcb9e0823(I273e0fe9c51c8549c8dfff393ca2e4e1);
            I05749703a8a131453c563ed2264680a7    = I77fe52c685b1075c294ac3c0a5b0d63a;

            Ifb1fc76002f6920a1f44c7b1bbcd0020 = I951dfff9507bb70214d48e03a0ebb3a7 + ~I4481555c402ba99bee05658ba6017984 + 1;
            Ia688029a35b4a62417906c9aa1cd7719 = I2bcab411f9bec1541259751bcb9e0823(Ifb1fc76002f6920a1f44c7b1bbcd0020);
            I4b76fe5f9863a41733b76decf9867d16    = Ia688029a35b4a62417906c9aa1cd7719;

            Idf6d4e3aa753aa396a9bffb27732f851 = I951dfff9507bb70214d48e03a0ebb3a7 + ~I9c68bfa3b888b6a6d41e38e674578284 + 1;
            Ifaaab2c6f368b133936a7295eeb9b45d = I2bcab411f9bec1541259751bcb9e0823(Idf6d4e3aa753aa396a9bffb27732f851);
            I2805bb16fd574a64de548b39a532cd8a    = Ifaaab2c6f368b133936a7295eeb9b45d;

            If14ca1f5d1c2977f9da79eaebaad1bf9 = I951dfff9507bb70214d48e03a0ebb3a7 + ~I6332af145d560e3f22a4a88106749f98 + 1;
            Ifbe064ac0a5f4bbf6caae486064a983d = I2bcab411f9bec1541259751bcb9e0823(If14ca1f5d1c2977f9da79eaebaad1bf9);
            Ide6a696c06f17f455d56bb28cad98bd0    = Ifbe064ac0a5f4bbf6caae486064a983d;

            If8f1505d9f10e30bd3320f500d34932f = I951dfff9507bb70214d48e03a0ebb3a7 + ~I35c0ca76b28cd2f9355276b5d2f29ad4 + 1;
            I439ac39c831e0ca87a40f49e439ce24f = I2bcab411f9bec1541259751bcb9e0823(If8f1505d9f10e30bd3320f500d34932f);
            I39bce1f71ede4663c187ddfd6501eda1    = I439ac39c831e0ca87a40f49e439ce24f;

            Id32aa77c6406b35a00168bb5452b12fb = Ie78e30b2a2eda75d0df7d10fd67b5e36 + ~I8cb171677016e4309034dc5d83981a48 + 1;
            I5c616021ebd98fc8e0fcf5b19732175c = I2bcab411f9bec1541259751bcb9e0823(Id32aa77c6406b35a00168bb5452b12fb);
            Id0e769bee61ae0a90c167fab061f5965    = I5c616021ebd98fc8e0fcf5b19732175c;

            I9a73686acefeb361337511f6943b036b = Ie78e30b2a2eda75d0df7d10fd67b5e36 + ~I4d1ba6ee8fb9505ba3b58b2b7553245b + 1;
            Id3a6c8114a92efaf5f6c280f897bef71 = I2bcab411f9bec1541259751bcb9e0823(I9a73686acefeb361337511f6943b036b);
            I83e03af8657a4a237641a9da7922e502    = Id3a6c8114a92efaf5f6c280f897bef71;

            Ib6eb7ce5a070f3a87bcf0e18be8c855d = Ie78e30b2a2eda75d0df7d10fd67b5e36 + ~Ib849494e5087777f646ee0947b4f634a + 1;
            I854d4e2867b459da2e2fc06c438e6077 = I2bcab411f9bec1541259751bcb9e0823(Ib6eb7ce5a070f3a87bcf0e18be8c855d);
            I7565e071282ca6e77bb469afc522f1a2    = I854d4e2867b459da2e2fc06c438e6077;

            If69b0b717c35d33fc8c0e59b07eb9edc = Ie78e30b2a2eda75d0df7d10fd67b5e36 + ~I283331db80e6d0891b13dc55e6a7d76c + 1;
            I3b334e8064cbfe97e70a0f4055496f04 = I2bcab411f9bec1541259751bcb9e0823(If69b0b717c35d33fc8c0e59b07eb9edc);
            I5d0dc5d40385ab67bc7f540f212b6a97    = I3b334e8064cbfe97e70a0f4055496f04;

            Ibb0d73078b779585e6b0e228391ecb96 = Ie78e30b2a2eda75d0df7d10fd67b5e36 + ~I0c1e4d400520935c5c78b792a9d554ba + 1;
            Iff92d12470884efa033800c88e1983e3 = I2bcab411f9bec1541259751bcb9e0823(Ibb0d73078b779585e6b0e228391ecb96);
            I548cac395730b8386670cc4c7a64319a    = Iff92d12470884efa033800c88e1983e3;

            I2894546e399fe3e33d7579772a1310df = Ie78e30b2a2eda75d0df7d10fd67b5e36 + ~I29da0e5661f29bd8493c19885c998582 + 1;
            I3d167f5af41902dc0a6477d55cf0abfd = I2bcab411f9bec1541259751bcb9e0823(I2894546e399fe3e33d7579772a1310df);
            Ic6d9bbbfb7890540edd10aa5758b0c4b    = I3d167f5af41902dc0a6477d55cf0abfd;

            I97f99a266267859aed199b278a430417 = Ia0b83a372dd4115dc4d61eb8ff0811b9 + ~If5b3850da967f6f3d7a71d680341ad1c + 1;
            Iaa7edba3767735cad1ec76479b5548b0 = I2bcab411f9bec1541259751bcb9e0823(I97f99a266267859aed199b278a430417);
            I7beb1f915a881a302f93c869d81417d1    = Iaa7edba3767735cad1ec76479b5548b0;

            Ie18cc792329941a3654322376a937d8d = Ia0b83a372dd4115dc4d61eb8ff0811b9 + ~Ic690477b1672dea4905a5e1c92b47366 + 1;
            Ifaa7aff0fb2af9d3e04b2641b13cf884 = I2bcab411f9bec1541259751bcb9e0823(Ie18cc792329941a3654322376a937d8d);
            I5fc389bbc1ce31f7b326da719dc576d4    = Ifaa7aff0fb2af9d3e04b2641b13cf884;

            Ie914a99f08d60b74c3c36a632a4ca9b0 = Ia0b83a372dd4115dc4d61eb8ff0811b9 + ~Ifa67d343acc6f3ec50c2b01fc26b4374 + 1;
            Ia78b9e9a1faddb38b4a1472f5eea3939 = I2bcab411f9bec1541259751bcb9e0823(Ie914a99f08d60b74c3c36a632a4ca9b0);
            I922e6f05f7c6e0f6f0b1a5c9548df238    = Ia78b9e9a1faddb38b4a1472f5eea3939;

            I82916e9dc3894ad88e12de01a68d6aa5 = Ia0b83a372dd4115dc4d61eb8ff0811b9 + ~Id27560fb44b4f2fda98d47e9f20d6898 + 1;
            I367d25430d8ec417123931f9534f3eba = I2bcab411f9bec1541259751bcb9e0823(I82916e9dc3894ad88e12de01a68d6aa5);
            I8c6bb234a1ca3deba637adf746672194    = I367d25430d8ec417123931f9534f3eba;

            I6cbf576b3d652e34c0221f8316b5a392 = Ia0b83a372dd4115dc4d61eb8ff0811b9 + ~I0807a826e91f92ef279ccf0b6512a428 + 1;
            I38a19bd51c6ee4fcb38493d869b7808a = I2bcab411f9bec1541259751bcb9e0823(I6cbf576b3d652e34c0221f8316b5a392);
            Ide24ebd7423d4c4f43577b019f2e30e4    = I38a19bd51c6ee4fcb38493d869b7808a;

            I9141b2516d7f855cd186472780af7b67 = Ia0b83a372dd4115dc4d61eb8ff0811b9 + ~I9426c8c1b4d988d5cd7d89a7aed4f8fc + 1;
            I0fe662c7d5cce9cf3cac56b6125852ff = I2bcab411f9bec1541259751bcb9e0823(I9141b2516d7f855cd186472780af7b67);
            Ifc412122eab7560c9021a17d7f8700c4    = I0fe662c7d5cce9cf3cac56b6125852ff;

            I07bf32ed72de9c02abf700c64853af61 = If5c5bcbbea01aa22f242b913f0d01929 + ~I7be8b2f8a9fe8e13001c2a1fce4a8a3f + 1;
            I6867bb41ee0a7f4c6ae0071e7975526d = I2bcab411f9bec1541259751bcb9e0823(I07bf32ed72de9c02abf700c64853af61);
            Ia5a56ed2c6b98e72002c6c5f946e7264    = I6867bb41ee0a7f4c6ae0071e7975526d;

            I52663a2999fb9571834d517538691b6f = If5c5bcbbea01aa22f242b913f0d01929 + ~I90a4190941651d885d04deb86a163365 + 1;
            I74d3dc7b6116f47b27dbfd112d7afd5d = I2bcab411f9bec1541259751bcb9e0823(I52663a2999fb9571834d517538691b6f);
            Ia888ed8885f66084b777f66e25cef1e7    = I74d3dc7b6116f47b27dbfd112d7afd5d;

            I8dcb88c94506367aabe8d7ed62cc56c2 = If5c5bcbbea01aa22f242b913f0d01929 + ~I24b4c998d19ae97f7178e37f75c77d06 + 1;
            I13440021cb8441969d3242de4fc6a0b5 = I2bcab411f9bec1541259751bcb9e0823(I8dcb88c94506367aabe8d7ed62cc56c2);
            I248229aecef00b87a70ce88920e407f5    = I13440021cb8441969d3242de4fc6a0b5;

            Ie676a4bee61154145391d9cc473fe91d = If5c5bcbbea01aa22f242b913f0d01929 + ~I0c121fa3e9e6e0e2e8291a594d6b4ceb + 1;
            Id3c71879c307df1390bbc60c55a5f249 = I2bcab411f9bec1541259751bcb9e0823(Ie676a4bee61154145391d9cc473fe91d);
            I3d162a0ec918f220a7d5f4efdf89cb58    = Id3c71879c307df1390bbc60c55a5f249;

            I9502c8fbf6b48749bf9f84a89a937dfe = If5c5bcbbea01aa22f242b913f0d01929 + ~I4319fa23d59f4e690e31fb7e3a823d17 + 1;
            I2e1fa8e49bf48184e6a669d18f5c8ced = I2bcab411f9bec1541259751bcb9e0823(I9502c8fbf6b48749bf9f84a89a937dfe);
            I1ca0372f60e48f2f803778c9017023c0    = I2e1fa8e49bf48184e6a669d18f5c8ced;

            I0c91e540e7106f32ae59491d8ed1853e = If5c5bcbbea01aa22f242b913f0d01929 + ~Ibd010f15e36194cbd2ce9f01c98a2b6f + 1;
            Ibc9c9339a0bcbc6addcce833051a8cd0 = I2bcab411f9bec1541259751bcb9e0823(I0c91e540e7106f32ae59491d8ed1853e);
            Ieb9693d54f0808b0ba463fd3c316a80e    = Ibc9c9339a0bcbc6addcce833051a8cd0;

            Iddfb8a8e261389eb4a2a10880c19446a = Iccba58cd3519fb4cc75a61b50da1d562 + ~I223151b6414d9979d71023053dd3f5e2 + 1;
            I2c0a2ad9eef6e84c60d1a6503aa836db = I2bcab411f9bec1541259751bcb9e0823(Iddfb8a8e261389eb4a2a10880c19446a);
            I63da03315d7e51fcacb0bc0298e506ed    = I2c0a2ad9eef6e84c60d1a6503aa836db;

            If0d55f861d4b3f0970c529024ca142d5 = Iccba58cd3519fb4cc75a61b50da1d562 + ~I6d6a242cdfadfc97fe656510bef73adc + 1;
            I3b06c3a23b2068e8f45870524c4af870 = I2bcab411f9bec1541259751bcb9e0823(If0d55f861d4b3f0970c529024ca142d5);
            I918f5a12e96bb96941f019940f27a5be    = I3b06c3a23b2068e8f45870524c4af870;

            Ib054f5d3f5cbb29a053d0e50c23cb3a8 = Iccba58cd3519fb4cc75a61b50da1d562 + ~I338400586daa58006c0a3dcd82ea8f4a + 1;
            I87d44c01b261e9c13add415e6b3cc5ba = I2bcab411f9bec1541259751bcb9e0823(Ib054f5d3f5cbb29a053d0e50c23cb3a8);
            Ib4fb115f442ff544fa3d21b4e9d3f075    = I87d44c01b261e9c13add415e6b3cc5ba;

            I1d65e9f97e93de8cc2a5dd532f8e482a = Iccba58cd3519fb4cc75a61b50da1d562 + ~I202c385beeccee309104b66f8f096b2c + 1;
            Ifc15e0dd91741676f23cc20fc542ec14 = I2bcab411f9bec1541259751bcb9e0823(I1d65e9f97e93de8cc2a5dd532f8e482a);
            I387403482432a3196109484d1120d584    = Ifc15e0dd91741676f23cc20fc542ec14;

            I3bdeab8c87325d46e45d9e2d44756934 = Iccba58cd3519fb4cc75a61b50da1d562 + ~I05a812cd935867d1e417c64c26ea0952 + 1;
            I50fdfffb4e2dbcf33282b3653f595ad0 = I2bcab411f9bec1541259751bcb9e0823(I3bdeab8c87325d46e45d9e2d44756934);
            I619af17eaa4a56726d6ab322a74dd0a4    = I50fdfffb4e2dbcf33282b3653f595ad0;

            If9228f7ecf19c41f4bbd8dabd0d5816c = Iccba58cd3519fb4cc75a61b50da1d562 + ~I7e86ab53e6d9647b230a94e076831ba2 + 1;
            I4e9786ec39d388cdce110c86bb436ae3 = I2bcab411f9bec1541259751bcb9e0823(If9228f7ecf19c41f4bbd8dabd0d5816c);
            I7a67ed3bb370520d0d25ce407ab8cd8b    = I4e9786ec39d388cdce110c86bb436ae3;

            I9e3edee214c4937d2aa462d3cffa624b = Ibc0999e4d0b3cc2650f9348b8c204b14 + ~I0e7ca2d6470b9bfc6a1ca6143b468507 + 1;
            I47cb30eb341ae7ce99042a16cd109f26 = I2bcab411f9bec1541259751bcb9e0823(I9e3edee214c4937d2aa462d3cffa624b);
            I7629b35ca548190a81021a2c13d8919b    = I47cb30eb341ae7ce99042a16cd109f26;

            I9fcbbd2e81b006b50e2d35ed2627bf83 = Ibc0999e4d0b3cc2650f9348b8c204b14 + ~I0aa5522190c741b7df4c4d7d34e46987 + 1;
            If004fa1c4e6bbe1f458c2d2a4f1f6e03 = I2bcab411f9bec1541259751bcb9e0823(I9fcbbd2e81b006b50e2d35ed2627bf83);
            I004851d3828f135ebe4d2e6ab83936bf    = If004fa1c4e6bbe1f458c2d2a4f1f6e03;

            Ie16f3d50ad5e5581ca099549db7232d2 = Ibc0999e4d0b3cc2650f9348b8c204b14 + ~Icf7630b6002db2f9b59d5323d6cc8105 + 1;
            I7c9910ade59c54e170c4f10822b5aff4 = I2bcab411f9bec1541259751bcb9e0823(Ie16f3d50ad5e5581ca099549db7232d2);
            I0e2c382b2e62ed43b76697230e34b719    = I7c9910ade59c54e170c4f10822b5aff4;

            I6345e93f3fa7f5eb2008dd41742afc2d = Ibc0999e4d0b3cc2650f9348b8c204b14 + ~Ia0ecfaedbc1d546d484978fd50096d10 + 1;
            I98939499dd98e583a4788cacc66c7fc4 = I2bcab411f9bec1541259751bcb9e0823(I6345e93f3fa7f5eb2008dd41742afc2d);
            I36dac27d10701db70fb2b5996a3f038f    = I98939499dd98e583a4788cacc66c7fc4;

            I698b93e10073b5d29357cde4bcac9dbe = I2aeff1fb4b839a581acaf26f90f9113c + ~Ib9322ec1d3866ba3cb42e96b5ff5cfb2 + 1;
            Ic530781e13180026815873e12550e405 = I2bcab411f9bec1541259751bcb9e0823(I698b93e10073b5d29357cde4bcac9dbe);
            I51d62ebd160eb0d073a7efb64d20079a    = Ic530781e13180026815873e12550e405;

            Ie7ced910d84655790823e6173a5a314a = I2aeff1fb4b839a581acaf26f90f9113c + ~If4d030e5858f325debc6f37abf4a7d6c + 1;
            Iba43927cdbcb6a80953fced163686073 = I2bcab411f9bec1541259751bcb9e0823(Ie7ced910d84655790823e6173a5a314a);
            Ib3545a88d68631af1c94ca2cb1f379af    = Iba43927cdbcb6a80953fced163686073;

            If6e3b6fd1810f6964e9024329d7cb3e3 = I2aeff1fb4b839a581acaf26f90f9113c + ~Ic35d5ac4dac46d47b2796bbac6452161 + 1;
            I29aefee3f95a7d2838ec5068515f69b0 = I2bcab411f9bec1541259751bcb9e0823(If6e3b6fd1810f6964e9024329d7cb3e3);
            I81ad7b044118734f4dc32a1a4e8eba31    = I29aefee3f95a7d2838ec5068515f69b0;

            If1045908c6d7476bd5507e57d08c406c = I2aeff1fb4b839a581acaf26f90f9113c + ~I27098cbe2d4fdd634385d771cc290c2b + 1;
            Ib964c4dd0a0ce2553766251b73018699 = I2bcab411f9bec1541259751bcb9e0823(If1045908c6d7476bd5507e57d08c406c);
            I5ad8c235d46349b6d310d0f175f84288    = Ib964c4dd0a0ce2553766251b73018699;

            I4d4f6705ed77a16ff31b34bae0d8b6d9 = I7d60d53f883f8187700c4e78b4c22f1c + ~Idfcf7f3240d92bfc87d44833bc00ff9d + 1;
            Ifd870cf74e7e3e5b348ad55af7242c27 = I2bcab411f9bec1541259751bcb9e0823(I4d4f6705ed77a16ff31b34bae0d8b6d9);
            Ibc00920378e2427df2a63a47dc3eaded    = Ifd870cf74e7e3e5b348ad55af7242c27;

            I70a492396580ac1143d8a2f4b181e873 = I7d60d53f883f8187700c4e78b4c22f1c + ~I73d2731c1b1ae5ef73ce0eb9c8995912 + 1;
            Ic4ba744721cdd747affca302b2b926d4 = I2bcab411f9bec1541259751bcb9e0823(I70a492396580ac1143d8a2f4b181e873);
            Ic5195bbaa69d95059cca6e152dc9f705    = Ic4ba744721cdd747affca302b2b926d4;

            I2fade32b5bdf245fa15289620dae2670 = I7d60d53f883f8187700c4e78b4c22f1c + ~Ia0caf6693d441ac622f416a86b665166 + 1;
            Id381e35622a3ac2c549a8c9b702ec020 = I2bcab411f9bec1541259751bcb9e0823(I2fade32b5bdf245fa15289620dae2670);
            Ia01f20e0bcf35c2ee4963e9c392c1004    = Id381e35622a3ac2c549a8c9b702ec020;

            Ie0dc166f57fea074496241a32cdb6015 = I7d60d53f883f8187700c4e78b4c22f1c + ~I5d7a0739e447775e00115799c52b11dd + 1;
            If49e3943165e2782c928a7da86847145 = I2bcab411f9bec1541259751bcb9e0823(Ie0dc166f57fea074496241a32cdb6015);
            I9f6f48fea88d1cd73ef2b24c7e819964    = If49e3943165e2782c928a7da86847145;

            If6a2518891412caa6d6d507082501f1e = Id6fcf4b7af4a37c854a12e2ae80851fa + ~Idd5b362dab4f93bba0c39af78c4c5981 + 1;
            Ie4d85aa4951d1a918d698c9e411b1ab2 = I2bcab411f9bec1541259751bcb9e0823(If6a2518891412caa6d6d507082501f1e);
            I847feea780cc8a06caea2d2ea79ad281    = Ie4d85aa4951d1a918d698c9e411b1ab2;

            Ic9912e5a838a377b26a19d22148a64df = Id6fcf4b7af4a37c854a12e2ae80851fa + ~I2a4b3573ae7c3b38ec34591f20c1d076 + 1;
            Iff6a8d4bc8f5f37d0ccc2d41f469ca86 = I2bcab411f9bec1541259751bcb9e0823(Ic9912e5a838a377b26a19d22148a64df);
            I7ef6f4aeda7fd6775839c068c681f9bc    = Iff6a8d4bc8f5f37d0ccc2d41f469ca86;

            Ibc0fca22d16444bc17877106ca772c31 = Id6fcf4b7af4a37c854a12e2ae80851fa + ~Ibb6e54edb9d277242c06d386a9a75a26 + 1;
            I6bed9b6e8b499c11d719f869467d2322 = I2bcab411f9bec1541259751bcb9e0823(Ibc0fca22d16444bc17877106ca772c31);
            I0645e741da20a4957747188273a655b1    = I6bed9b6e8b499c11d719f869467d2322;

            Ie4291d233597d5d676a80fd62d9bd208 = Id6fcf4b7af4a37c854a12e2ae80851fa + ~Ie95793e09085b6de1383a37cc7fc41ac + 1;
            Id1db54a136ab42fe675fa77b2b7fd2de = I2bcab411f9bec1541259751bcb9e0823(Ie4291d233597d5d676a80fd62d9bd208);
            I71125dffdd2d37e44dbb46143c1e8d9a    = Id1db54a136ab42fe675fa77b2b7fd2de;

            Ifc13b798d76aa70ec1877c275fb31d36 = Ifa5e5f7d753964f14f0f16dbe552fd85 + ~I627e4bdc8061c69e3fcac17535b9f1e0 + 1;
            Ia6ed9442d22d3228ce14749ffdacfab2 = I2bcab411f9bec1541259751bcb9e0823(Ifc13b798d76aa70ec1877c275fb31d36);
            I50c166f958b22ce866cd40334918274c    = Ia6ed9442d22d3228ce14749ffdacfab2;

            I57d6637f0bdab578a790e4a12ccaa16b = Ifa5e5f7d753964f14f0f16dbe552fd85 + ~I28ea268c5b51ac1d9249e96599bb6b0d + 1;
            I32e0c22a86e88cadc6a956c213ff992c = I2bcab411f9bec1541259751bcb9e0823(I57d6637f0bdab578a790e4a12ccaa16b);
            Icd225144fd331b870847044b4d02bed0    = I32e0c22a86e88cadc6a956c213ff992c;

            If8ea04fe685b4f20cdaf9a84984d56fe = Ifa5e5f7d753964f14f0f16dbe552fd85 + ~Ib97b2670a6cd88b2327f07f62d887900 + 1;
            I1b0dcddcb3e0a398857f038d3a52e719 = I2bcab411f9bec1541259751bcb9e0823(If8ea04fe685b4f20cdaf9a84984d56fe);
            I5e876482090ce6007c2a2f2101c24654    = I1b0dcddcb3e0a398857f038d3a52e719;

            Ie0c86f20c28bcbe410b191b90d29bf76 = Ifa5e5f7d753964f14f0f16dbe552fd85 + ~I134a734d93e62f6ac6635015fe3a2096 + 1;
            I8c6bcabb8814607901102aca5f820293 = I2bcab411f9bec1541259751bcb9e0823(Ie0c86f20c28bcbe410b191b90d29bf76);
            I026ded06f56d9ca93f47fd85aec4f7ad    = I8c6bcabb8814607901102aca5f820293;

            I3dc5d3f66726e15968a70cbf3d3b656a = Ifa5e5f7d753964f14f0f16dbe552fd85 + ~Ib24b68cb35da39a743e1d90bba3f0836 + 1;
            I731089de22b5becf3621097ed7a81b7e = I2bcab411f9bec1541259751bcb9e0823(I3dc5d3f66726e15968a70cbf3d3b656a);
            Iec596e94ec168a564bccbbaa7df833c9    = I731089de22b5becf3621097ed7a81b7e;

            Id674686e7ac37fd6f63846f9a9cede19 = I900d471b087cf5a436c2ad66a84d8280 + ~I5ca15c7da1f49580ddedd9ff8ba822c0 + 1;
            Ifb3674681315fa8cf6739996b823a7aa = I2bcab411f9bec1541259751bcb9e0823(Id674686e7ac37fd6f63846f9a9cede19);
            Ib514e01c261e43a725582a10596eed32    = Ifb3674681315fa8cf6739996b823a7aa;

            Ie2ed9668d13d219c60f2e0614488cd42 = I900d471b087cf5a436c2ad66a84d8280 + ~I6aba8ca0e4b20a6355b43a70f19d9d8c + 1;
            I2d5ef5bf9c28065a2a4ab718fbc8ba3e = I2bcab411f9bec1541259751bcb9e0823(Ie2ed9668d13d219c60f2e0614488cd42);
            Ic19a62cdecb2329370f7e11c48d3738d    = I2d5ef5bf9c28065a2a4ab718fbc8ba3e;

            I98abc995ff89934534543be93c6e3ffa = I900d471b087cf5a436c2ad66a84d8280 + ~Ie9a316de516ec4fb828a614c67e38b2a + 1;
            I7c5f9c301a0bdbf642f7b3f33e9bfc66 = I2bcab411f9bec1541259751bcb9e0823(I98abc995ff89934534543be93c6e3ffa);
            Ib2f5691baa59adfbaad62f6ffc71fb05    = I7c5f9c301a0bdbf642f7b3f33e9bfc66;

            I579cf9386ab7b08efa204d735335e462 = I900d471b087cf5a436c2ad66a84d8280 + ~I745187336b8a5ae4eac66e90539752cf + 1;
            I7bde3bcef8556c1b1e4c7d2192196e00 = I2bcab411f9bec1541259751bcb9e0823(I579cf9386ab7b08efa204d735335e462);
            I9bdfaca6112385deb86e24ad7e45bbaa    = I7bde3bcef8556c1b1e4c7d2192196e00;

            I9efa4d729d10a6b7cc335fb765ed032c = I900d471b087cf5a436c2ad66a84d8280 + ~Id4cdd72193e90dddd211af73d7f3634a + 1;
            Id13f3a39b334d8a80b7c8286b09bd1e1 = I2bcab411f9bec1541259751bcb9e0823(I9efa4d729d10a6b7cc335fb765ed032c);
            I0e647bb8351cfe7828423e7099525585    = Id13f3a39b334d8a80b7c8286b09bd1e1;

            If9191ebc8e88d4e75f0f35897ebb1421 = I6d1434907f0292ea2ee47cbc5b52bfb9 + ~I276c2ce5d3a1b7551c2790971071b094 + 1;
            Ie6443f42260e0a2983927d0940c82a06 = I2bcab411f9bec1541259751bcb9e0823(If9191ebc8e88d4e75f0f35897ebb1421);
            I185b758fb3e50bcfb1464fe2ab593cfe    = Ie6443f42260e0a2983927d0940c82a06;

            I3511287cfe69d5cedc5a8fbcad708437 = I6d1434907f0292ea2ee47cbc5b52bfb9 + ~I77fd8001d879fc9e9117464fba27902d + 1;
            I43003b2ef41b34363169f004a6668a59 = I2bcab411f9bec1541259751bcb9e0823(I3511287cfe69d5cedc5a8fbcad708437);
            Ie25e944f9e3100c39b69bb38dffca177    = I43003b2ef41b34363169f004a6668a59;

            I91812179d44cb675b90d477f33ec48ad = I6d1434907f0292ea2ee47cbc5b52bfb9 + ~I6d0d098e6d47dea04d6d7be67b648a0d + 1;
            Ic385923d90d69cd387eb9fb5f62fd9ba = I2bcab411f9bec1541259751bcb9e0823(I91812179d44cb675b90d477f33ec48ad);
            I8e77032a54376578b3d16799e30c97f7    = Ic385923d90d69cd387eb9fb5f62fd9ba;

            Idb04a1aae91fdc477ca38ed66789ee88 = I6d1434907f0292ea2ee47cbc5b52bfb9 + ~Ic3c59a5167cb83fd76ec6236572b1f3d + 1;
            I2f642acd0cb0bd30177bc0d65751ed99 = I2bcab411f9bec1541259751bcb9e0823(Idb04a1aae91fdc477ca38ed66789ee88);
            I4cd2a7f8f8ec378200b00d03e447ac92    = I2f642acd0cb0bd30177bc0d65751ed99;

            I566054aece562960590ee28b157e4a3e = I6d1434907f0292ea2ee47cbc5b52bfb9 + ~Iccab4c19a9190689f90a42160e2379de + 1;
            If1064670adff5b00cbf7809e2621cfd5 = I2bcab411f9bec1541259751bcb9e0823(I566054aece562960590ee28b157e4a3e);
            I1b3c55aca0da232cf3f81d6d0914729f    = If1064670adff5b00cbf7809e2621cfd5;

            I7b2ffb762cd9ef7aa8ba224efb75c46c = I938bef7ba7ae1739d8e6a6a7c117a1b1 + ~Iff777b2c4a3939e330c4cbb36cbe1ac5 + 1;
            I72311a2c7557be2b6cb95b3bc6f511a5 = I2bcab411f9bec1541259751bcb9e0823(I7b2ffb762cd9ef7aa8ba224efb75c46c);
            I34c76f1a126120c4474e750e9b51e034    = I72311a2c7557be2b6cb95b3bc6f511a5;

            Id90bbb642b0f4434d8a148a28b6b2f65 = I938bef7ba7ae1739d8e6a6a7c117a1b1 + ~Iedf37dac8b3a5331277ae4f0176968aa + 1;
            I79ee4c7277f713aa710ae8cf7c470aa1 = I2bcab411f9bec1541259751bcb9e0823(Id90bbb642b0f4434d8a148a28b6b2f65);
            I0edb624c344787066a2267757052196b    = I79ee4c7277f713aa710ae8cf7c470aa1;

            Ia4e297e35d484b15adce7e1d67f582b0 = I938bef7ba7ae1739d8e6a6a7c117a1b1 + ~I3f6fad8bb0fba790fcdb1612b6fa7712 + 1;
            I32bfef7a7ecaa533e3bf92fb560e657b = I2bcab411f9bec1541259751bcb9e0823(Ia4e297e35d484b15adce7e1d67f582b0);
            Ia8443f199838742595ac114f35c00143    = I32bfef7a7ecaa533e3bf92fb560e657b;

            I84996b1d03b692f6f736fb04c7f91e83 = I938bef7ba7ae1739d8e6a6a7c117a1b1 + ~Idc549661d6694035874a3366704801c7 + 1;
            If4a6b6a8b44d2c55c93b111d20525ec6 = I2bcab411f9bec1541259751bcb9e0823(I84996b1d03b692f6f736fb04c7f91e83);
            Ib25b8a538c9d64880e114bf4a80ca42e    = If4a6b6a8b44d2c55c93b111d20525ec6;

            I83078cc7857fc17b30f640854a4d6be5 = I938bef7ba7ae1739d8e6a6a7c117a1b1 + ~I275ea08a3dc0600d8ccb6300eb7f2a6b + 1;
            I7d41f27ff64d549b7e5df6b172969d8a = I2bcab411f9bec1541259751bcb9e0823(I83078cc7857fc17b30f640854a4d6be5);
            I25f6a3d7bb869082e4dbbd0ee8574c95    = I7d41f27ff64d549b7e5df6b172969d8a;

            I94bb467129904032736fb13dd636c600 = I6384a9416b2d1da01df1b2d7b16c5390 + ~I0a9cb91319cc0d0c1c4d0020cce321d7 + 1;
            Ie3a2d4d85d4e4ac011887cbd329bd9b7 = I2bcab411f9bec1541259751bcb9e0823(I94bb467129904032736fb13dd636c600);
            If96057023747a1538d9f06966af48bc2    = Ie3a2d4d85d4e4ac011887cbd329bd9b7;

            Ifa76758b50f439170ecd6d86ff898bc4 = I6384a9416b2d1da01df1b2d7b16c5390 + ~I9dff504e40aaddefedbb7b0f822c844a + 1;
            I3bc9fcec69ab6a1efb2d86e03804415c = I2bcab411f9bec1541259751bcb9e0823(Ifa76758b50f439170ecd6d86ff898bc4);
            I199e995390462e06853b1f5cdbd46e0a    = I3bc9fcec69ab6a1efb2d86e03804415c;

            I9d831dd976e8cd5d8f6a6818601e6424 = I6384a9416b2d1da01df1b2d7b16c5390 + ~Id9edc6ac95a260bf5af3de25f00e9e9c + 1;
            I9ee16e46a399d1445fcdf251757a5e43 = I2bcab411f9bec1541259751bcb9e0823(I9d831dd976e8cd5d8f6a6818601e6424);
            Iec6325d585ddd0a9f86bb5cd0229960d    = I9ee16e46a399d1445fcdf251757a5e43;

            I474774ae149804412ed4aaf1cdcaba88 = I6384a9416b2d1da01df1b2d7b16c5390 + ~If0676ef300628c4097565b13ef2d8854 + 1;
            I45cf986a60a429a68051f76beb8188fb = I2bcab411f9bec1541259751bcb9e0823(I474774ae149804412ed4aaf1cdcaba88);
            I4be1ccfec148a522fbf5b8375245cbb3    = I45cf986a60a429a68051f76beb8188fb;

            I964cdcb4e6b49a62d30c2a2540851317 = I6384a9416b2d1da01df1b2d7b16c5390 + ~I1b53098a7240d2b5dc1f5c5c3b4bcc11 + 1;
            I4e48461fcd58a133a09d856852887a4f = I2bcab411f9bec1541259751bcb9e0823(I964cdcb4e6b49a62d30c2a2540851317);
            I074386ff6a3d8d644f4b2501c69f26c7    = I4e48461fcd58a133a09d856852887a4f;

            I6df268bc9f85ce88674a9165664ea84a = I5097a79e7cf7a30d38ba198d1407119c + ~I1cff7306aaf303bb3342ea3d72048908 + 1;
            I901714025da5b89ee929ea2859f3e6c7 = I2bcab411f9bec1541259751bcb9e0823(I6df268bc9f85ce88674a9165664ea84a);
            I83b378e5534c553b57beb22c5178a3ce    = I901714025da5b89ee929ea2859f3e6c7;

            I74fdcbe9f49f7bce1f5e31d956c5883c = I5097a79e7cf7a30d38ba198d1407119c + ~I2d839c10960739097d449efab58b9fd4 + 1;
            I976786b0539b07b056dad0f050eeb53f = I2bcab411f9bec1541259751bcb9e0823(I74fdcbe9f49f7bce1f5e31d956c5883c);
            I14f79d67f75af6a495d6eb2986210cda    = I976786b0539b07b056dad0f050eeb53f;

            I4a1b8453cb7a21745d5f74ad05653ed2 = I5097a79e7cf7a30d38ba198d1407119c + ~I080832c25509f7003ed50d71210bc7f7 + 1;
            I8e1ad4f44dcac3e770dd862413b25a4e = I2bcab411f9bec1541259751bcb9e0823(I4a1b8453cb7a21745d5f74ad05653ed2);
            Iacd805413ec1eb001b3083554f187554    = I8e1ad4f44dcac3e770dd862413b25a4e;

            I9c53b478b2011fac0615a152fe60d5b6 = I5097a79e7cf7a30d38ba198d1407119c + ~Idb73eba1bd4ce25a6109e296f51e7dc4 + 1;
            Iaf5caa6558f0a98b91fb72db734bbec4 = I2bcab411f9bec1541259751bcb9e0823(I9c53b478b2011fac0615a152fe60d5b6);
            I3e61e09fcc81a0011a79f5c5ce77bc46    = Iaf5caa6558f0a98b91fb72db734bbec4;

            Id75dbed8f1a5befda32c60b994681013 = I5097a79e7cf7a30d38ba198d1407119c + ~I278659ca1a0b093fc883d01987989dc0 + 1;
            I7b37d3b1b23f09c6ac46a94cf2c4ead7 = I2bcab411f9bec1541259751bcb9e0823(Id75dbed8f1a5befda32c60b994681013);
            I6e6cbb7dba8eb3c02b5b4e4469e23cea    = I7b37d3b1b23f09c6ac46a94cf2c4ead7;

            I378a59323b74623c5524f854d6e11226 = Ib113c26c8dcf49c972c41a938059a787 + ~Id033e7adfcfb0420cc592a1fb6c297b6 + 1;
            Ief8b577d924f257ae5e1dd47009b0db2 = I2bcab411f9bec1541259751bcb9e0823(I378a59323b74623c5524f854d6e11226);
            I8b25822c33f7d506ef69216af3fdab44    = Ief8b577d924f257ae5e1dd47009b0db2;

            I080bf885464a0cc948a4450e9f7d1d26 = Ib113c26c8dcf49c972c41a938059a787 + ~Ia443284a35e0873de59b3ae55b7f809d + 1;
            Ie59366fcd6132a48f3e9be1bb5b600c6 = I2bcab411f9bec1541259751bcb9e0823(I080bf885464a0cc948a4450e9f7d1d26);
            I06fd642cbc8aa2f65197801d7459cfa2    = Ie59366fcd6132a48f3e9be1bb5b600c6;

            If769e73adea227de1fd85c2e89d0ba08 = Ib113c26c8dcf49c972c41a938059a787 + ~I2b807c16cfc6d65cb2a7f28ffa837974 + 1;
            I273c1e28c3ed897b7d0f6b36a3a8def9 = I2bcab411f9bec1541259751bcb9e0823(If769e73adea227de1fd85c2e89d0ba08);
            I22202e6c3de9b06c04ce9514af28933e    = I273c1e28c3ed897b7d0f6b36a3a8def9;

            Ifa6a34b83225e9d9b28b14874c4444e3 = Ib113c26c8dcf49c972c41a938059a787 + ~Ie467c5fde1d123da4e9587b5a56748a0 + 1;
            I64b507fe58b933919d0766631985a74e = I2bcab411f9bec1541259751bcb9e0823(Ifa6a34b83225e9d9b28b14874c4444e3);
            Ib991cdbb91133cb82e154c575e00a174    = I64b507fe58b933919d0766631985a74e;

            I584b1d4d6fb7ee4f20ad9c96715cdf90 = Ib113c26c8dcf49c972c41a938059a787 + ~If92e66cba66732798dd19f968a5ef8ce + 1;
            I7c0376cbc3660f3d82a5da22806ef5e3 = I2bcab411f9bec1541259751bcb9e0823(I584b1d4d6fb7ee4f20ad9c96715cdf90);
            I5590364df6874420e169aa444ab520b9    = I7c0376cbc3660f3d82a5da22806ef5e3;

            I265f9b91fbb62164e589dcf96818c4f5 = I970c4a25a8bce82a9d2846679029fcab + ~I4ba05e74c2f63e2f4c59268775d549aa + 1;
            I3884d561185660e7e0f461b3487fdfd4 = I2bcab411f9bec1541259751bcb9e0823(I265f9b91fbb62164e589dcf96818c4f5);
            I43a9e393037fb4aa84741dca22648459    = I3884d561185660e7e0f461b3487fdfd4;

            I3d59a47c88227734cf6fc0d6fd30db11 = I970c4a25a8bce82a9d2846679029fcab + ~I8289bfc08a5d8979ec26825bcb6e3d18 + 1;
            I4b991f90354e3f74d105a64929a97d6f = I2bcab411f9bec1541259751bcb9e0823(I3d59a47c88227734cf6fc0d6fd30db11);
            Ibb4d8301d90c66fdfac92b3fbc53c019    = I4b991f90354e3f74d105a64929a97d6f;

            I6144b6df2c87ea0948d730343b42129f = I970c4a25a8bce82a9d2846679029fcab + ~I2b32537c9178028493af165398a60875 + 1;
            I9534939768f7d2532ca4e6757dfafb72 = I2bcab411f9bec1541259751bcb9e0823(I6144b6df2c87ea0948d730343b42129f);
            Ibae217fa4b808e4accbeb8f4a9a976ab    = I9534939768f7d2532ca4e6757dfafb72;

            Ia7ca7400e36ea572fba8e19bcc81ecbd = I970c4a25a8bce82a9d2846679029fcab + ~I18d0dd7a10d6533f721a2392d4ad2d02 + 1;
            I090228a60e5919fa88d842b1638ee296 = I2bcab411f9bec1541259751bcb9e0823(Ia7ca7400e36ea572fba8e19bcc81ecbd);
            Ia8bd7a3594f7084a57e64da023bf784c    = I090228a60e5919fa88d842b1638ee296;

            I302e61b49accf5db556b87517f2341f5 = I970c4a25a8bce82a9d2846679029fcab + ~I784c4e9fb75c314f271477e0621aaf7c + 1;
            I8994d511d611a3c1b7a8122cd3d2825e = I2bcab411f9bec1541259751bcb9e0823(I302e61b49accf5db556b87517f2341f5);
            I3ce4b9d41f5472bf60ed2802a2ab10eb    = I8994d511d611a3c1b7a8122cd3d2825e;

            I5d9af1abff6efe3a55c6568d936b6ec7 = Ibe2af096ad2db26e54d8b4b3bb05175c + ~I299b37fd45c6ee2031fb2c74caac73be + 1;
            I43d14ec8853bfd211aa6b887c7ebdd5a = I2bcab411f9bec1541259751bcb9e0823(I5d9af1abff6efe3a55c6568d936b6ec7);
            I93ec9bc6fbd056e7e52496546493e727    = I43d14ec8853bfd211aa6b887c7ebdd5a;

            I8cde0aa611c476b5112edeb8f17f15bf = Ibe2af096ad2db26e54d8b4b3bb05175c + ~Ib8603cb82ceb97c2f35bf8209306a457 + 1;
            Icd810cceba64ffbb087600155338911c = I2bcab411f9bec1541259751bcb9e0823(I8cde0aa611c476b5112edeb8f17f15bf);
            I2374b90dde1cf481baa40af31e1a43e3    = Icd810cceba64ffbb087600155338911c;

            Icaa40ec40d6d26cdf70bb5ae7d492e47 = Ibe2af096ad2db26e54d8b4b3bb05175c + ~I18916d0023ca275d84c52af07dcc5ca2 + 1;
            I33ddd4cdef0a0704f204f4fdb14fd859 = I2bcab411f9bec1541259751bcb9e0823(Icaa40ec40d6d26cdf70bb5ae7d492e47);
            I0cee595f488a909ade8a3b4c90dbb0c7    = I33ddd4cdef0a0704f204f4fdb14fd859;

            I8346f15d822cacfeecbe5d75412cb53f = Ibe2af096ad2db26e54d8b4b3bb05175c + ~Ic7d5fe6c4b1dcb97d10ba3de2f95d1df + 1;
            I0c87f78f08ac77246d7b3b8604dfd700 = I2bcab411f9bec1541259751bcb9e0823(I8346f15d822cacfeecbe5d75412cb53f);
            Iba4c3d91d492b000ab1de7add9f171a9    = I0c87f78f08ac77246d7b3b8604dfd700;

            I5ee364aab320ab40c0f65feda6f53b18 = Ibe2af096ad2db26e54d8b4b3bb05175c + ~I3d3aafdd4d9d3e9fdab1f487c48a0ea9 + 1;
            I54745c58c61eba829e4717cd842d519d = I2bcab411f9bec1541259751bcb9e0823(I5ee364aab320ab40c0f65feda6f53b18);
            I2b4152aa4c51cc1c1ffabac78cea267c    = I54745c58c61eba829e4717cd842d519d;

            I1f0ecba054900f96cd7100741191c5f4 = Ie48569c467fba0c1291f71d6080ebedc + ~I26bdcc44692db066911c8d5b0a1aae0c + 1;
            I9e278d7b6cccaa39163d0867427709ed = I2bcab411f9bec1541259751bcb9e0823(I1f0ecba054900f96cd7100741191c5f4);
            Ie4c3dd5c191aff00a6d62006223c2b76    = I9e278d7b6cccaa39163d0867427709ed;

            I4faf2caf62966416118a54015908c889 = Ie48569c467fba0c1291f71d6080ebedc + ~I8d26e73fafa909f1e26e329828cf4888 + 1;
            I3e5d8af6fed6b47aebf2eef7010afa8b = I2bcab411f9bec1541259751bcb9e0823(I4faf2caf62966416118a54015908c889);
            Ie4c0ba9510f9b924999bb5f432137271    = I3e5d8af6fed6b47aebf2eef7010afa8b;

            Idd0329980a36f87859150530ab44b52d = Ie48569c467fba0c1291f71d6080ebedc + ~I2c72d6c5fa6968dffa6517cf81219875 + 1;
            Ie96538fd32c8f8d7a3144012d10b29a5 = I2bcab411f9bec1541259751bcb9e0823(Idd0329980a36f87859150530ab44b52d);
            I5bad544a17b384973d5672acbe0ac0d5    = Ie96538fd32c8f8d7a3144012d10b29a5;

            Ie66bc10dde27f08813d4d347fd7cf6ce = Ie48569c467fba0c1291f71d6080ebedc + ~I05aabdf73200996b7bea8db700fa8930 + 1;
            I050a226112c903de442358e2d5be8274 = I2bcab411f9bec1541259751bcb9e0823(Ie66bc10dde27f08813d4d347fd7cf6ce);
            I231bfb8e19e1d9c4bbd29a0bd75c1ed3    = I050a226112c903de442358e2d5be8274;

            Ie1d8b3ea7c6603cebf2f9adb776910b7 = Ie48569c467fba0c1291f71d6080ebedc + ~Idb4c722992139f39914af7085378c6cc + 1;
            I4df410c6a7eea67fd73cc33c791e7aa0 = I2bcab411f9bec1541259751bcb9e0823(Ie1d8b3ea7c6603cebf2f9adb776910b7);
            I1ecf87e33de04d02db9e64590bcaffde    = I4df410c6a7eea67fd73cc33c791e7aa0;

            Ia37488e9a50cf5cc08de74ade676db96 = I90e7ded06617b49cdb8b5301fe9c6a20 + ~Iaee91a5e94c3f174682f72a1ebfd0021 + 1;
            Id7e318f124e0534c8e0538f99616ed01 = I2bcab411f9bec1541259751bcb9e0823(Ia37488e9a50cf5cc08de74ade676db96);
            I60c97bf58193f004e3fcfdbd6a03ce6e    = Id7e318f124e0534c8e0538f99616ed01;

            I08aa45211cab01d567cd5eb172fd2f0c = I90e7ded06617b49cdb8b5301fe9c6a20 + ~Ibc1a16427d8dfa5ee20dac15327a53ea + 1;
            I66ba7e48a07f5fdfe16d23b0dc243514 = I2bcab411f9bec1541259751bcb9e0823(I08aa45211cab01d567cd5eb172fd2f0c);
            Ib71065a3fe70d3ab5f05b0c393278631    = I66ba7e48a07f5fdfe16d23b0dc243514;

            If4ff0c63ec1deb46412858e496451a01 = I90e7ded06617b49cdb8b5301fe9c6a20 + ~Ic1120eb027841908cd64fe5c7274da14 + 1;
            I62e6e8be411f12cd5c4d63f1825521f3 = I2bcab411f9bec1541259751bcb9e0823(If4ff0c63ec1deb46412858e496451a01);
            I984074a5c77445ad266463e20d77899e    = I62e6e8be411f12cd5c4d63f1825521f3;

            Ife7bfd15fc4c392b5d2288d9a4e879b3 = I90e7ded06617b49cdb8b5301fe9c6a20 + ~I4ee3f608cc8f8df27345949f1a3713a7 + 1;
            I2f94d5aad80c081124e3efa3804af183 = I2bcab411f9bec1541259751bcb9e0823(Ife7bfd15fc4c392b5d2288d9a4e879b3);
            I50bb40691aa09c42e0b64a076b50a971    = I2f94d5aad80c081124e3efa3804af183;

            I24ac26debafd03c7333d174e8725afd6 = I90e7ded06617b49cdb8b5301fe9c6a20 + ~I63c9deb7e6a4b400e0aff6887a09e647 + 1;
            I7a91b23716bf81bea4956eafb467c96a = I2bcab411f9bec1541259751bcb9e0823(I24ac26debafd03c7333d174e8725afd6);
            I753bff437b6c563f5fddf19685405504    = I7a91b23716bf81bea4956eafb467c96a;

            I99d80ad68e2563d0f78a0e3bb82c5328 = I4920014f5d017f4e840dc3b88526955f + ~Iaed26e1c4a2578d16b111d15d31339d2 + 1;
            I17572136bb435e84505c016523a6ec88 = I2bcab411f9bec1541259751bcb9e0823(I99d80ad68e2563d0f78a0e3bb82c5328);
            I21f2ec69bcc507756e2a5f85d3ead3e8    = I17572136bb435e84505c016523a6ec88;

            I9943733ef305983c629565c881054bbf = I4920014f5d017f4e840dc3b88526955f + ~Ifc52604a4f9f9de392a35f2f9fe885b8 + 1;
            I9b0ac56afa21022e8bc69f5d20d17b66 = I2bcab411f9bec1541259751bcb9e0823(I9943733ef305983c629565c881054bbf);
            Iddec4486996054e475499d370016a685    = I9b0ac56afa21022e8bc69f5d20d17b66;

            I7cb4420bc55c03a6500f5228d31fe43c = I4920014f5d017f4e840dc3b88526955f + ~I4037f1b207aa101f354e59eddd7c9eb4 + 1;
            Id9468cba18d4c67a84cb2b16d2cf495e = I2bcab411f9bec1541259751bcb9e0823(I7cb4420bc55c03a6500f5228d31fe43c);
            I3d3edd06f8907f4369b825062348da87    = Id9468cba18d4c67a84cb2b16d2cf495e;

            Ic4d19dec464359c0a9fa75148fe90c73 = I4920014f5d017f4e840dc3b88526955f + ~Ic0a580f94f3d03f72e3a487f84bf6612 + 1;
            I2bda0265c40a5cedc359dee75fb15b4c = I2bcab411f9bec1541259751bcb9e0823(Ic4d19dec464359c0a9fa75148fe90c73);
            I72467ef10ecced8395a6870a39525787    = I2bda0265c40a5cedc359dee75fb15b4c;

            I44993416e1d22613dbd78402c37a934d = I4920014f5d017f4e840dc3b88526955f + ~Ie6f67c6e4c5e2b8357c0a902979e8722 + 1;
            I318ebdf91ab8e83b80a880395879fc77 = I2bcab411f9bec1541259751bcb9e0823(I44993416e1d22613dbd78402c37a934d);
            I9b74b672f55e7bf7560ba4dd2d0c79fd    = I318ebdf91ab8e83b80a880395879fc77;

            Ibc9b94a9dea471805cb442ac6904bc97 = I03b70553f1c501609400574ae7cd73f5 + ~Ibafedcf9f2990ed9c1efa973a0b1d81d + 1;
            I8ac8dbc25a20c0c27e09240a5cd1bfd2 = I2bcab411f9bec1541259751bcb9e0823(Ibc9b94a9dea471805cb442ac6904bc97);
            I285b012d2fb5e2279a79cf8edca24ac8    = I8ac8dbc25a20c0c27e09240a5cd1bfd2;

            I917d9f9b144d3bffafc77bddae7fba6b = I03b70553f1c501609400574ae7cd73f5 + ~Icf4405d4a4063448a2be8ad0354ab1a8 + 1;
            Id8c4e5d6318622bd8ec2974684f542b6 = I2bcab411f9bec1541259751bcb9e0823(I917d9f9b144d3bffafc77bddae7fba6b);
            I8faf911a7d1ea8b0abe54f6688068ca0    = Id8c4e5d6318622bd8ec2974684f542b6;

            Ibc91c6c3d56bb8a14e22909c43ffec51 = I03b70553f1c501609400574ae7cd73f5 + ~I778fbaea65beeb6de599490daf3b7e3c + 1;
            I8df19e0871c18890419c593410596b59 = I2bcab411f9bec1541259751bcb9e0823(Ibc91c6c3d56bb8a14e22909c43ffec51);
            I3dca974bf2d5631a47ebf8b945efab20    = I8df19e0871c18890419c593410596b59;

            If7c2d3eddd96b47b6c2aea8b27c8c7f4 = I03b70553f1c501609400574ae7cd73f5 + ~I1d7a4f99e3975fd01bfe5a9a1da84765 + 1;
            Ifb977d4c5bac50b9d7f2f814a500f0f2 = I2bcab411f9bec1541259751bcb9e0823(If7c2d3eddd96b47b6c2aea8b27c8c7f4);
            I12141c45d147b058a9e392f3b7d7d06e    = Ifb977d4c5bac50b9d7f2f814a500f0f2;

            I4df093ed94d26b058e97db550e347e3c = I63c9bf68b43ed66c51b0f4c0ed92e9ab + ~Ie3c88bc240576aa220f0f110b13bfdd3 + 1;
            Id9a1f5bd846dc7d093ed9392722317be = I2bcab411f9bec1541259751bcb9e0823(I4df093ed94d26b058e97db550e347e3c);
            Ia527c96e30b782f837bc6206961400e4    = Id9a1f5bd846dc7d093ed9392722317be;

            Ie90303b0326bee4ab203a8cf1e643da9 = I63c9bf68b43ed66c51b0f4c0ed92e9ab + ~Ibc8679379ddc43ee4bc508a1f577eb2c + 1;
            Ic886ecf946cd5c297012444cb34980ab = I2bcab411f9bec1541259751bcb9e0823(Ie90303b0326bee4ab203a8cf1e643da9);
            I6adbdb64422a08be9bf9e538db97463b    = Ic886ecf946cd5c297012444cb34980ab;

            I19030d352fd059156ee42c66f9270beb = I63c9bf68b43ed66c51b0f4c0ed92e9ab + ~Id66798f8ea67e74a67f264fe6b4503a3 + 1;
            I37085a233f195dce1a76d05b0157fcac = I2bcab411f9bec1541259751bcb9e0823(I19030d352fd059156ee42c66f9270beb);
            I958cdf5367c7b0bd58b70b763d3af8aa    = I37085a233f195dce1a76d05b0157fcac;

            I36767a902c53a384128ae1443cf88963 = I63c9bf68b43ed66c51b0f4c0ed92e9ab + ~I059d847e09f5aa3f6a8147062f4b13bf + 1;
            Ia2812d1ba8ca6831a2f059eb23384b38 = I2bcab411f9bec1541259751bcb9e0823(I36767a902c53a384128ae1443cf88963);
            I91b7b8e8887b5dd9853297463c55b78d    = Ia2812d1ba8ca6831a2f059eb23384b38;

            I868dffa3f07407f7996bb5bc596939b7 = If408dfead07757878cc878131bc7d6a3 + ~I4ed5da534afbfe9ecbc10ef4cc649a55 + 1;
            Id176f2681568337762559e78cde29ba6 = I2bcab411f9bec1541259751bcb9e0823(I868dffa3f07407f7996bb5bc596939b7);
            I6162978f0c57958ad0403246fb0530dd    = Id176f2681568337762559e78cde29ba6;

            I7d928be164d0dce8b1322ff230c053e9 = If408dfead07757878cc878131bc7d6a3 + ~Ie2e3d64640c339dc51512979dbd6a173 + 1;
            Ia0c4e9942a4b08f69c2a027a712c9e39 = I2bcab411f9bec1541259751bcb9e0823(I7d928be164d0dce8b1322ff230c053e9);
            I508142e70fd04513977130556aa574ef    = Ia0c4e9942a4b08f69c2a027a712c9e39;

            I98be4971a8a9a08abb3ebe474d7f0c6d = If408dfead07757878cc878131bc7d6a3 + ~I772e844c41387e7079259875e0ba3fa0 + 1;
            I2da299005fed6f2b710e25acd48ebe91 = I2bcab411f9bec1541259751bcb9e0823(I98be4971a8a9a08abb3ebe474d7f0c6d);
            I2afab673e4b803ffd888f187de47fa49    = I2da299005fed6f2b710e25acd48ebe91;

            I779e70dea33201e9237f29681ffd5e27 = If408dfead07757878cc878131bc7d6a3 + ~I48e5256ade4d061a3b5ba08a53252bc3 + 1;
            Ia1038e3b807e16a30f6f4564509ddd30 = I2bcab411f9bec1541259751bcb9e0823(I779e70dea33201e9237f29681ffd5e27);
            I7a56f81596920126a9ea2c9fb3a19285    = Ia1038e3b807e16a30f6f4564509ddd30;

            Ie2262914042172ab7e08599278f36af5 = Ia0857d63d309807789b6ff4f6028f1b3 + ~Ice8765807beffd3acf59fa137ee0baac + 1;
            I25d94516522c19c0e53b5f52f4480216 = I2bcab411f9bec1541259751bcb9e0823(Ie2262914042172ab7e08599278f36af5);
            Ic6252de2c819f2243476ddf82e22d137    = I25d94516522c19c0e53b5f52f4480216;

            I4001323da8f7956cdd480ac2d56df929 = Ia0857d63d309807789b6ff4f6028f1b3 + ~I6e4786234b286b12c83e06e93c628534 + 1;
            I4b96be53e3d059113bb74b27ffe30179 = I2bcab411f9bec1541259751bcb9e0823(I4001323da8f7956cdd480ac2d56df929);
            Ieea8672b2f23711c6ba893de5c5d8bc2    = I4b96be53e3d059113bb74b27ffe30179;

            Ib1cd6731034887a0a55e405c9db3e8de = Ia0857d63d309807789b6ff4f6028f1b3 + ~I3e8e280553edaa5c8555ace81ecc10e0 + 1;
            Ic091d8daff9f609c53cb191ed6b6ddeb = I2bcab411f9bec1541259751bcb9e0823(Ib1cd6731034887a0a55e405c9db3e8de);
            I3a4dbdf517b8f9c93b567f91870e6160    = Ic091d8daff9f609c53cb191ed6b6ddeb;

            I51aa496e8c03944c28a908102514e6f8 = Ia0857d63d309807789b6ff4f6028f1b3 + ~I635fb29c55e0fb5cff0b6f443c2e3de5 + 1;
            I2468caeaf9733c8bc6a485542b6b263f = I2bcab411f9bec1541259751bcb9e0823(I51aa496e8c03944c28a908102514e6f8);
            I4731ee7a0e08c69e2bd2a8bcea0838c2    = I2468caeaf9733c8bc6a485542b6b263f;

            I6415f3996318472532e161510ccc8ca3 = I53921b825c5e434b63bee0e1ecb7a517 + ~Ic2f450f7ab60ba57dfc1406c92c0f077 + 1;
            I6611d1fa58dd253fe6344a41584d7e22 = I2bcab411f9bec1541259751bcb9e0823(I6415f3996318472532e161510ccc8ca3);
            I1b6cbbcf01a65cd1c2f1e241f849c904    = I6611d1fa58dd253fe6344a41584d7e22;

            Ia11b671b59240988737979328c472812 = I53921b825c5e434b63bee0e1ecb7a517 + ~I529eaa7e5eeb6d0a1aba78df5d5a2fa0 + 1;
            I8afb33eced17e8675a8e2bd90d16030b = I2bcab411f9bec1541259751bcb9e0823(Ia11b671b59240988737979328c472812);
            I663aee79f824c854f57c19e87207529b    = I8afb33eced17e8675a8e2bd90d16030b;

            Id4fabe0165a117a402dc14f2f3ec626a = I53921b825c5e434b63bee0e1ecb7a517 + ~I839895c8614ff28df83314c44824900b + 1;
            Idac55755226133905d3250273b1eccb8 = I2bcab411f9bec1541259751bcb9e0823(Id4fabe0165a117a402dc14f2f3ec626a);
            I34ff7299c9d83affa4512b7da302c199    = Idac55755226133905d3250273b1eccb8;

            I57238f501ab7278b308d76211ced8cf7 = I53921b825c5e434b63bee0e1ecb7a517 + ~Iede5d56e52612e083407888da49470e5 + 1;
            I4cd564459b8d65976195b2994e7d44f2 = I2bcab411f9bec1541259751bcb9e0823(I57238f501ab7278b308d76211ced8cf7);
            I70ca6c9d0a5c99e0036479f7b5dd760a    = I4cd564459b8d65976195b2994e7d44f2;

            I9b257f8556ca4e5402637f01081b78e1 = I53921b825c5e434b63bee0e1ecb7a517 + ~I088c5b971a2def57248769a33b7d2a2d + 1;
            I2280162ee1c08ccc9f0c17d1ca0e3628 = I2bcab411f9bec1541259751bcb9e0823(I9b257f8556ca4e5402637f01081b78e1);
            I835bb7345787eaadc41816858e0a71a1    = I2280162ee1c08ccc9f0c17d1ca0e3628;

            I2e093412a9fa3972cea01664389d8c27 = I5e68f84e123c37f19a03c13892c77e19 + ~Id144785da9b171f1e2d0e9182d693e31 + 1;
            I28b3ba64175358f277427fd790a9228b = I2bcab411f9bec1541259751bcb9e0823(I2e093412a9fa3972cea01664389d8c27);
            I3c7f6fdd0e9cc7426df76027912d1ccb    = I28b3ba64175358f277427fd790a9228b;

            I17907fd8c6975c8c642535ff929221a6 = I5e68f84e123c37f19a03c13892c77e19 + ~I439c7c302b535bfd7db655c3c607d71f + 1;
            I6c03138440f9bd0cb2cfe12abf619c10 = I2bcab411f9bec1541259751bcb9e0823(I17907fd8c6975c8c642535ff929221a6);
            I9ff512085174a7720705d0fb37c4ec34    = I6c03138440f9bd0cb2cfe12abf619c10;

            I3c6577b04ad56d864bbaa2c048323c11 = I5e68f84e123c37f19a03c13892c77e19 + ~I2a0dc4ed573a544cb13544e049514903 + 1;
            Ib3709eb9dfc3a594d38ea5a0ef0cd444 = I2bcab411f9bec1541259751bcb9e0823(I3c6577b04ad56d864bbaa2c048323c11);
            I6a69cdf2bae1ea68c9be56dcc4e76a59    = Ib3709eb9dfc3a594d38ea5a0ef0cd444;

            I6f0c341c05eaa8f35bbce4521f6e8f94 = I5e68f84e123c37f19a03c13892c77e19 + ~I39d9044227c161f0163e58dd82aadc90 + 1;
            I44cf5ba18d7d029df13f446f09191b2c = I2bcab411f9bec1541259751bcb9e0823(I6f0c341c05eaa8f35bbce4521f6e8f94);
            I855ddead34ac131137ba644afbfea2b7    = I44cf5ba18d7d029df13f446f09191b2c;

            Ib72ba950ecf9ae2668374f6633a67ca7 = I5e68f84e123c37f19a03c13892c77e19 + ~Ide22394fce1658f9e7002bdb30d03c2f + 1;
            I6aa1e5acf0c2b01c94438bd1cff484c6 = I2bcab411f9bec1541259751bcb9e0823(Ib72ba950ecf9ae2668374f6633a67ca7);
            Ib1a463388daf270eb0ce698d7b5ded4b    = I6aa1e5acf0c2b01c94438bd1cff484c6;

            I3d7c72d725f4563bb562e2992093cb02 = Id5270b57c6fb4b18db3bbd0a523e467e + ~I0cd8a6e719305ee3fbe8228081993957 + 1;
            Ia23629f3881e4119c36576f7da58ceaa = I2bcab411f9bec1541259751bcb9e0823(I3d7c72d725f4563bb562e2992093cb02);
            I74e4bb7530c02073f9b15a6389659d4b    = Ia23629f3881e4119c36576f7da58ceaa;

            I813c881ac61a59041be3be78f6a466c8 = Id5270b57c6fb4b18db3bbd0a523e467e + ~I583c6d23506c7d7b84403bfe977ec1ec + 1;
            I2f12d1fa0b815564cefafc28ceb3de82 = I2bcab411f9bec1541259751bcb9e0823(I813c881ac61a59041be3be78f6a466c8);
            I6721b13abeddc76139bdc7380434cc2a    = I2f12d1fa0b815564cefafc28ceb3de82;

            I866510e7dc721fa5aac312bc5ab5ba0a = Id5270b57c6fb4b18db3bbd0a523e467e + ~Ia422fbdf8f318ff3ddc049d1374e7939 + 1;
            Ib09ac099bcf61b09922b353403b29987 = I2bcab411f9bec1541259751bcb9e0823(I866510e7dc721fa5aac312bc5ab5ba0a);
            I84fba239c5705bcd92096e204cc9438c    = Ib09ac099bcf61b09922b353403b29987;

            Ib4432359f97849dff6ad3e0f044157bd = Id5270b57c6fb4b18db3bbd0a523e467e + ~I8efad9622c05177563ab8a2747879044 + 1;
            I3c2b6da8e286d0a7b628ba1071f29424 = I2bcab411f9bec1541259751bcb9e0823(Ib4432359f97849dff6ad3e0f044157bd);
            I4d46e4d50176768fda897949545e2125    = I3c2b6da8e286d0a7b628ba1071f29424;

            Ic86aa6eb1b4dcc2520309089b43292e6 = Id5270b57c6fb4b18db3bbd0a523e467e + ~I9ff276a14d3205b98174a8a736f79774 + 1;
            I550630b507ceec38b960ab2a86a57f1a = I2bcab411f9bec1541259751bcb9e0823(Ic86aa6eb1b4dcc2520309089b43292e6);
            I57086cfab3b163c3911c3cf7bfb3141a    = I550630b507ceec38b960ab2a86a57f1a;

            I0731115afe5c15bcf131f7ef4f05802b = I3c18a84617eb21472d53e598700d7f4c + ~Ic566fe27ccaf2220101cbc49fc187a6b + 1;
            I795c1c91cb6b7870b7efb07d67085be1 = I2bcab411f9bec1541259751bcb9e0823(I0731115afe5c15bcf131f7ef4f05802b);
            Ice174debd5dc911fdf5d5756cff8d731    = I795c1c91cb6b7870b7efb07d67085be1;

            Ib080b8fd34385aa7986dace4afd95267 = I3c18a84617eb21472d53e598700d7f4c + ~I618363a8ac413dd0ee52eb658940eaed + 1;
            I531b70d12349f3bc67e6a3ec53368d97 = I2bcab411f9bec1541259751bcb9e0823(Ib080b8fd34385aa7986dace4afd95267);
            Ie369670edc5b602d305904f3a4a4381f    = I531b70d12349f3bc67e6a3ec53368d97;

            I134890b77451d0b78afc7402a6a28048 = I3c18a84617eb21472d53e598700d7f4c + ~I1d648ed8f07f0743a6d616584270c513 + 1;
            Id8a109043bc922b718c203bd5d60a999 = I2bcab411f9bec1541259751bcb9e0823(I134890b77451d0b78afc7402a6a28048);
            I41f66f79339962ef42fab3b88e571170    = Id8a109043bc922b718c203bd5d60a999;

            I956da75f13433c1dd7a3cbd3b78922c1 = I3c18a84617eb21472d53e598700d7f4c + ~I03038b940be8bd21bd26b150b28754a6 + 1;
            Ic126109499ee1dc2787ab05b404e7ae2 = I2bcab411f9bec1541259751bcb9e0823(I956da75f13433c1dd7a3cbd3b78922c1);
            I5cbd2fad4d90bd77ba3d2448a37ac60f    = Ic126109499ee1dc2787ab05b404e7ae2;

            I440b26c9f1b9ccf70f97c9d5f732d38e = I3c18a84617eb21472d53e598700d7f4c + ~I123255637493b9c7924e3a72d1b86ee9 + 1;
            I1cd8ba53b876e2436901749e355f354b = I2bcab411f9bec1541259751bcb9e0823(I440b26c9f1b9ccf70f97c9d5f732d38e);
            Id86a2869148e2885633d9e277f7041c3    = I1cd8ba53b876e2436901749e355f354b;

            I5e3a441faca44bffc4368d96d8fb0bfd = Id36663e7a01fff3170833ecfecac1321 + ~I2133d362ba45ceb3dceaa84e95ace1e6 + 1;
            I4e8ff51a6f70f8ca6a17a1dea8caf0a9 = I2bcab411f9bec1541259751bcb9e0823(I5e3a441faca44bffc4368d96d8fb0bfd);
            Ifb7b585189db23efabfb522c9b45bede    = I4e8ff51a6f70f8ca6a17a1dea8caf0a9;

            I21d7ba25247a87a1a9c245d0d1f553b0 = Id36663e7a01fff3170833ecfecac1321 + ~Ib43383830037df764b48c637a28ab6b5 + 1;
            Ic1a27480c9acc1684f3fed116d74cb5f = I2bcab411f9bec1541259751bcb9e0823(I21d7ba25247a87a1a9c245d0d1f553b0);
            I7763f0d28d8065d8c94ef8df96b2ab06    = Ic1a27480c9acc1684f3fed116d74cb5f;

            I55aafa8162cfc4fccfae68cf78cd1c2b = Id36663e7a01fff3170833ecfecac1321 + ~If2ce7b8d2573494564393f7d426fa47f + 1;
            I0df7a888610865486aa1aaa2703dd041 = I2bcab411f9bec1541259751bcb9e0823(I55aafa8162cfc4fccfae68cf78cd1c2b);
            I115ba88588187c7115977e95bd26ee5a    = I0df7a888610865486aa1aaa2703dd041;

            Ib99c25f0d8d6493cac4d5c816884c704 = Id36663e7a01fff3170833ecfecac1321 + ~Ied4ddedaf801fbd7238d8a55c17c8090 + 1;
            If6448c72403a3d0bd904beac87f8aa96 = I2bcab411f9bec1541259751bcb9e0823(Ib99c25f0d8d6493cac4d5c816884c704);
            I6e7f2bdd0c8231a3689893ef4877fdba    = If6448c72403a3d0bd904beac87f8aa96;

            Iee7c9f0a0e8ca127efee008b4874edbd = Id36663e7a01fff3170833ecfecac1321 + ~I87e6ef84894cfc86b94e19c9d3065bc6 + 1;
            Iecf45496b391208d62e88544b5d2ca49 = I2bcab411f9bec1541259751bcb9e0823(Iee7c9f0a0e8ca127efee008b4874edbd);
            I546c513d5357ac1a6fe669888dfaf717    = Iecf45496b391208d62e88544b5d2ca49;

            I17b4a3baae65161387f472037ffc6fc4 = I8d3be15109c7007a79fecaac0d891626 + ~I768afe193d9d79b136736abc6846d945 + 1;
            Ib0fd0a839c85f3da5ae7b221f6e623d6 = I2bcab411f9bec1541259751bcb9e0823(I17b4a3baae65161387f472037ffc6fc4);
            Ib3e12c614471912d0b276cb9f0382b1b    = Ib0fd0a839c85f3da5ae7b221f6e623d6;

            Ie7b7b202a968fe73f6b1e02a044414c5 = I8d3be15109c7007a79fecaac0d891626 + ~I0aa93075086164fdbab3814d60633141 + 1;
            Ie045750c9289c899860823f90a306f3c = I2bcab411f9bec1541259751bcb9e0823(Ie7b7b202a968fe73f6b1e02a044414c5);
            I7187a2499e3319da90b6d6fc64411b46    = Ie045750c9289c899860823f90a306f3c;

            I479ab5c0e483c36267d8248340006666 = I8d3be15109c7007a79fecaac0d891626 + ~I32c35da92922c5b477f8aba837fa6d92 + 1;
            I1627b19e0ca42f9c264b626809fb37b7 = I2bcab411f9bec1541259751bcb9e0823(I479ab5c0e483c36267d8248340006666);
            I9b46582473bb4dd5541a35ac708486f4    = I1627b19e0ca42f9c264b626809fb37b7;

            I777bfe165e25d7fde4fc950f23db7b84 = I8d3be15109c7007a79fecaac0d891626 + ~Ibf547f8a5e1059ffaabeb3f447904dcf + 1;
            Ic9593f3fe23f258c2ab4ddcadaa8ca4c = I2bcab411f9bec1541259751bcb9e0823(I777bfe165e25d7fde4fc950f23db7b84);
            I929796fe327ee9c8a05e6bb683ae5d7c    = Ic9593f3fe23f258c2ab4ddcadaa8ca4c;

            I146d505a34ddb8d65e0a1769f623a7fd = I8d3be15109c7007a79fecaac0d891626 + ~I4c32900878260a261bc5403e8abd6258 + 1;
            Idc0085a6595a7de7e2bc87c789b7d935 = I2bcab411f9bec1541259751bcb9e0823(I146d505a34ddb8d65e0a1769f623a7fd);
            Ib6638da8b69373c2026d3f5305825cde    = Idc0085a6595a7de7e2bc87c789b7d935;

            Ia85239bddc04bf50bcf037ed2f76d7ac = I92169cc57291f20d336a479e392ec271 + ~I54166b387c02e12374d6febc425bfb7a + 1;
            Id029b4c310acea870263d3715689e729 = I2bcab411f9bec1541259751bcb9e0823(Ia85239bddc04bf50bcf037ed2f76d7ac);
            I28c26bf4cf9693d1807818b2ca7883ac    = Id029b4c310acea870263d3715689e729;

            Ia7306bacf3c2b180d3261a5c1f0f4a30 = I92169cc57291f20d336a479e392ec271 + ~If06a1563b9d7348de03a98d31bd85b06 + 1;
            Iec123ddb8d1e623d03d85a667c97ef31 = I2bcab411f9bec1541259751bcb9e0823(Ia7306bacf3c2b180d3261a5c1f0f4a30);
            I291fc4eef4b80d1020c96488b869727e    = Iec123ddb8d1e623d03d85a667c97ef31;

            I2018147b86e47af5842c4f29d047d157 = I92169cc57291f20d336a479e392ec271 + ~I3e466d40a4447a23953d96d2e6d61d47 + 1;
            I89f0b0713e165a454e187fa51e89c642 = I2bcab411f9bec1541259751bcb9e0823(I2018147b86e47af5842c4f29d047d157);
            I53006ed50f6211439681aa7659647e35    = I89f0b0713e165a454e187fa51e89c642;

            Id17a85459845f8a8be694c4bf1fc29c9 = I92169cc57291f20d336a479e392ec271 + ~I3b2739319710681986b9d3f8cd04f619 + 1;
            Id812cf3919ed50a5e3897d129eeb4b8d = I2bcab411f9bec1541259751bcb9e0823(Id17a85459845f8a8be694c4bf1fc29c9);
            I47fe32973727237ae0cd4c306c7efbfb    = Id812cf3919ed50a5e3897d129eeb4b8d;

            Ic012b15584d9d25af38f83d0526503da = I92169cc57291f20d336a479e392ec271 + ~Ifc100357ae3f754fb0e3863334bcc764 + 1;
            I2d65b5115be2a22ed1e29426be3f0d15 = I2bcab411f9bec1541259751bcb9e0823(Ic012b15584d9d25af38f83d0526503da);
            Ic3e0c7d71f13a56a9a63e158c7f2cfa8    = I2d65b5115be2a22ed1e29426be3f0d15;

            I7f09bd4a45143a036ce04af11b9927f9 = I6178b220b469b40dac39168057023a1c + ~Icb2805685607d5fedd0300c9d800f863 + 1;
            I47c8671569e2c5c2a21f27aff2d1f4b8 = I2bcab411f9bec1541259751bcb9e0823(I7f09bd4a45143a036ce04af11b9927f9);
            If383f241447cbea4e18f4f79fcdbf144    = I47c8671569e2c5c2a21f27aff2d1f4b8;

            Ica32f94af6e6f3eaf2b724a2173fa463 = I6178b220b469b40dac39168057023a1c + ~I28fa295ebd90c2b7255d48ca9ffcfcf3 + 1;
            Iaf2144dab2167cd2629067e40bea3053 = I2bcab411f9bec1541259751bcb9e0823(Ica32f94af6e6f3eaf2b724a2173fa463);
            Ia05354d3b4f61299d5897832639df2c2    = Iaf2144dab2167cd2629067e40bea3053;

            Ib750bb83ddfbbad2a2be8d1c8392b4ff = I6178b220b469b40dac39168057023a1c + ~I4fd45670f88265e5d7aa6582f3ad3ff8 + 1;
            I4c2b80e4bbbd4c5e8d0da28c5d0f681e = I2bcab411f9bec1541259751bcb9e0823(Ib750bb83ddfbbad2a2be8d1c8392b4ff);
            I9faec40665477e8b3237773d606af2f0    = I4c2b80e4bbbd4c5e8d0da28c5d0f681e;

            I3906ece39480f96020717c6243e8ba4c = I6178b220b469b40dac39168057023a1c + ~I5f607bdc9b276fdf07a17a11a20a6720 + 1;
            I6300fbbd385ad9280c751076bc68d70c = I2bcab411f9bec1541259751bcb9e0823(I3906ece39480f96020717c6243e8ba4c);
            Id231ab3133d4bed02aad7e5f560ee5f0    = I6300fbbd385ad9280c751076bc68d70c;

            Ie68ce21ade07fa53c30ebf27216b03f9 = I6178b220b469b40dac39168057023a1c + ~Iefe9e5376010997c0ee52eeb28e57a25 + 1;
            Iea078843b3c5139a395997c54462850a = I2bcab411f9bec1541259751bcb9e0823(Ie68ce21ade07fa53c30ebf27216b03f9);
            I13616c8c7be221cf4d2c13ae87c38bed    = Iea078843b3c5139a395997c54462850a;

            I6cc6fa167c0d2b4b62ddbeecea175ed2 = I55342938216a0ea0889f96c2f6c05ce5 + ~Ieca5b21b91e150c9d509964bdcea500d + 1;
            I654debf65019f2748e631a051f3b17ca = I2bcab411f9bec1541259751bcb9e0823(I6cc6fa167c0d2b4b62ddbeecea175ed2);
            I8793bc728a4d423fb96a88c83bb9746f    = I654debf65019f2748e631a051f3b17ca;

            Ibddf3468ae7c27d5a4b1388e524aa9c2 = I55342938216a0ea0889f96c2f6c05ce5 + ~Icaeb9a2ec8ec5822658fa85b88cca04b + 1;
            I1e88b57c19a1ddfc1c1f0e168b60f814 = I2bcab411f9bec1541259751bcb9e0823(Ibddf3468ae7c27d5a4b1388e524aa9c2);
            I2fb6af0f152232550a3cadd55656df20    = I1e88b57c19a1ddfc1c1f0e168b60f814;

            Iadcb2b3acaac2e1bb505c65d3cbe4235 = I55342938216a0ea0889f96c2f6c05ce5 + ~I76e4c55148effeba62a4837cd19c5e51 + 1;
            Ibaf7ab7333434b0d7e76e436ee40a406 = I2bcab411f9bec1541259751bcb9e0823(Iadcb2b3acaac2e1bb505c65d3cbe4235);
            I5144918fcd4ce1a061644240730fc52a    = Ibaf7ab7333434b0d7e76e436ee40a406;

            I37cd96b8b0a4939d9a70098fd8bcf452 = I55342938216a0ea0889f96c2f6c05ce5 + ~Ie6060acdcb16b6fa6aeeb649ed621053 + 1;
            I1af14572832bd6d6b5890b8340b79ec7 = I2bcab411f9bec1541259751bcb9e0823(I37cd96b8b0a4939d9a70098fd8bcf452);
            I1821eb21cdf8208ff6c2f28d963f7bd6    = I1af14572832bd6d6b5890b8340b79ec7;

            Ib34b169dcc76daee2d1aa2b2a7513af3 = Idf28431c76a84a48dd895979d2b11a63 + ~I6b7a8ba12de5b44817ec99faebe54617 + 1;
            I652d3ed935b39f8fda8d84296456d633 = I2bcab411f9bec1541259751bcb9e0823(Ib34b169dcc76daee2d1aa2b2a7513af3);
            I80471575b1d4b69ef073056f798394ea    = I652d3ed935b39f8fda8d84296456d633;

            If36fc316d6ec7c7e09eae77807b37099 = Idf28431c76a84a48dd895979d2b11a63 + ~I58416287b268462d28f55c6c2705e613 + 1;
            I5e33cad360aae934f418852541f5f2bd = I2bcab411f9bec1541259751bcb9e0823(If36fc316d6ec7c7e09eae77807b37099);
            I890bf9b72cc3c71351547178d72796e5    = I5e33cad360aae934f418852541f5f2bd;

            Ifd214c332218ac5c0fe5aded4b952711 = Idf28431c76a84a48dd895979d2b11a63 + ~I2d636a246d815a4d12c478794860dd40 + 1;
            If950e448e3cba7cc9aa7aff7718775f7 = I2bcab411f9bec1541259751bcb9e0823(Ifd214c332218ac5c0fe5aded4b952711);
            Icc9d28b84fa91028ae96cc9b8bae7555    = If950e448e3cba7cc9aa7aff7718775f7;

            Idcd0fc8f86e2b6f03606b818b8346e5a = Idf28431c76a84a48dd895979d2b11a63 + ~I46c2b923860b0d1c01b9475f4467f280 + 1;
            I9adf8836419a1c85b146e5e36de68af5 = I2bcab411f9bec1541259751bcb9e0823(Idcd0fc8f86e2b6f03606b818b8346e5a);
            I0b0d167c415f8c14594bd61907d46d80    = I9adf8836419a1c85b146e5e36de68af5;

            If486aa8ac2cfb46f936714812cc760df = I1ef61124c8d62e8f6a82a729fb091694 + ~I9b8cfdb69b76453a3ac687a1e098417f + 1;
            I0f2bcdf124dff4219fd1a35ed1db7937 = I2bcab411f9bec1541259751bcb9e0823(If486aa8ac2cfb46f936714812cc760df);
            I9577d49a74520355e53a1818f479db0e    = I0f2bcdf124dff4219fd1a35ed1db7937;

            I2d8e5b5fdbda7d599423c38aaace6658 = I1ef61124c8d62e8f6a82a729fb091694 + ~Ib2963b82260024e1853d297798d88d3c + 1;
            Iae82e5de28b12f962bd7c5e221317ac2 = I2bcab411f9bec1541259751bcb9e0823(I2d8e5b5fdbda7d599423c38aaace6658);
            Ie6e888d582ba9e600e91b119e2804642    = Iae82e5de28b12f962bd7c5e221317ac2;

            I6d0878fb7ec75c0a26be4dbba62f80dc = I1ef61124c8d62e8f6a82a729fb091694 + ~Id59cf860d9f4aff11b205b8970d93df3 + 1;
            Ia7b3cb9de8e18f41561c2a46dda8696a = I2bcab411f9bec1541259751bcb9e0823(I6d0878fb7ec75c0a26be4dbba62f80dc);
            Iccfac3d489b4b110d6b6e005a5ba45d8    = Ia7b3cb9de8e18f41561c2a46dda8696a;

            I16a16ff0e8a6685a09803634da429fd2 = I1ef61124c8d62e8f6a82a729fb091694 + ~I38b4eceb159ecb0dda3920290a21a02a + 1;
            Id0119672c8b017bce6fdba53d4dccf8b = I2bcab411f9bec1541259751bcb9e0823(I16a16ff0e8a6685a09803634da429fd2);
            I69a67481ca8fd01dc5400dbe887b4f83    = Id0119672c8b017bce6fdba53d4dccf8b;

            Idb211abaa54ac26e7379c64a63f7d07c = Ib8bb96f0372323e6a8072ca56fb9396d + ~Ibf9f6d7baed9e761b69fb41442761ac6 + 1;
            I4aaef2f654ba03b1dc05719c81d5da69 = I2bcab411f9bec1541259751bcb9e0823(Idb211abaa54ac26e7379c64a63f7d07c);
            I1f36f045becec7f0528f4a935d3da2ff    = I4aaef2f654ba03b1dc05719c81d5da69;

            I351205eb71acb31b59d2b4470f0ba28c = Ib8bb96f0372323e6a8072ca56fb9396d + ~Ie945349d77442536992d9ad52ce84218 + 1;
            Ia6355e548635a4107a11c7952aa8b3d9 = I2bcab411f9bec1541259751bcb9e0823(I351205eb71acb31b59d2b4470f0ba28c);
            I530fe7720e3bcda35e940aa4973a7da4    = Ia6355e548635a4107a11c7952aa8b3d9;

            If5660c495bf7690252783d888d1ad6e8 = Ib8bb96f0372323e6a8072ca56fb9396d + ~I3bc01b072987a0c980615abbc2251e5f + 1;
            I0bd950eee6abde9d1eaaabbe902fff5d = I2bcab411f9bec1541259751bcb9e0823(If5660c495bf7690252783d888d1ad6e8);
            I03069dda9fa863172d8747408800eeba    = I0bd950eee6abde9d1eaaabbe902fff5d;

            I3a5229cb8e44a15560b5c7bef96e65cc = Ib8bb96f0372323e6a8072ca56fb9396d + ~Ic45561ffe1837c3d5bb42c695a377f82 + 1;
            I93caf487f67a2adce04a7b2cd7fff358 = I2bcab411f9bec1541259751bcb9e0823(I3a5229cb8e44a15560b5c7bef96e65cc);
            Ie7f36ee89f2b092555fbf8031d2347d9    = I93caf487f67a2adce04a7b2cd7fff358;

            I889b9b0828e97fe44d8366c5ef71a8f2 = I432f74dda4f6b1cebdf5ad59c659080b + ~I67534b68fee8f76ac0c5e64cd02aba42 + 1;
            If68a9cc5609ea7d87062bad2ebddb1a8 = I2bcab411f9bec1541259751bcb9e0823(I889b9b0828e97fe44d8366c5ef71a8f2);
            I18af7980562b28c537be3bea8dc5252b    = If68a9cc5609ea7d87062bad2ebddb1a8;

            Ie23062e00e39ead706f5b6ead233747d = I432f74dda4f6b1cebdf5ad59c659080b + ~Ic79072d9e42dbc9974231f1d642b3f12 + 1;
            If201a7afedfd1c329b55048e6bbad629 = I2bcab411f9bec1541259751bcb9e0823(Ie23062e00e39ead706f5b6ead233747d);
            I22ec20f9396d28ed39c5fc4bf060c44a    = If201a7afedfd1c329b55048e6bbad629;

            I8a2589544c75ecfdc31d28912c639695 = I432f74dda4f6b1cebdf5ad59c659080b + ~If08adda7d796da7c7849e472a73282a3 + 1;
            I1f8936599ead5ce1cd85132e382533f1 = I2bcab411f9bec1541259751bcb9e0823(I8a2589544c75ecfdc31d28912c639695);
            I105eac4e38f4661c7c7ca32161e42baa    = I1f8936599ead5ce1cd85132e382533f1;

            I5c21c59147e9c3a74c7cbbb6f2a23919 = I432f74dda4f6b1cebdf5ad59c659080b + ~I3db0adb3457cb22c755f5d29a8fe7ed8 + 1;
            I37eb148270af62adba8341c83411f9f2 = I2bcab411f9bec1541259751bcb9e0823(I5c21c59147e9c3a74c7cbbb6f2a23919);
            I5030734bfa54065cbef20c1350cd647d    = I37eb148270af62adba8341c83411f9f2;

            Idacd78e24408e432abbbfb0c447fdde5 = I432f74dda4f6b1cebdf5ad59c659080b + ~I3e76abc721bf7ed186f4d0f8f4bbf4e3 + 1;
            Ie4729048b95fede1806dbd006de01338 = I2bcab411f9bec1541259751bcb9e0823(Idacd78e24408e432abbbfb0c447fdde5);
            Ieccf25e3abd6bae7dcf08baf815f3439    = Ie4729048b95fede1806dbd006de01338;

            I0e8b171fe5080485a7f4fef83f1f1528 = Idc689442305acd00f0f32416d8fb3773 + ~I277d7065150714e33d8ba64875d18190 + 1;
            I02330d212434a6e8c303db2c3d36a3e5 = I2bcab411f9bec1541259751bcb9e0823(I0e8b171fe5080485a7f4fef83f1f1528);
            I600c21fca7901299f8e95e8fa0ea0eb0    = I02330d212434a6e8c303db2c3d36a3e5;

            Ib22c2bd76e6c29cc2f1440885bf24b7b = Idc689442305acd00f0f32416d8fb3773 + ~I9bb4d58b1fe80549451b00c4ed2b3885 + 1;
            Id89498cf205e0cdef4886afd878c48f6 = I2bcab411f9bec1541259751bcb9e0823(Ib22c2bd76e6c29cc2f1440885bf24b7b);
            Ic4363dfd133124dd45ec2211499d0788    = Id89498cf205e0cdef4886afd878c48f6;

            I149559fccd9def4ec1ead1fdcff3c7fd = Idc689442305acd00f0f32416d8fb3773 + ~Ie335e68643fd2b0a53351f4bd45c3475 + 1;
            I547ae5055196f12eeeb36d69c325b84d = I2bcab411f9bec1541259751bcb9e0823(I149559fccd9def4ec1ead1fdcff3c7fd);
            I7c0bc779c09847e3beb0a139e8826511    = I547ae5055196f12eeeb36d69c325b84d;

            Icfa8fed3239748abca27a5fc17de79c0 = Idc689442305acd00f0f32416d8fb3773 + ~I32679702c19eab37b46d13bb372967ea + 1;
            I4871ccbe2f182791243b7bdcc9b8e286 = I2bcab411f9bec1541259751bcb9e0823(Icfa8fed3239748abca27a5fc17de79c0);
            If64db4386bf8f7d07292f14e3b313520    = I4871ccbe2f182791243b7bdcc9b8e286;

            I2ff115fa483f080d93bada49a9566b33 = Idc689442305acd00f0f32416d8fb3773 + ~I1afb4061458e9d2f5799afa1f2373bd2 + 1;
            I12fd829f22ba908180290432320a3660 = I2bcab411f9bec1541259751bcb9e0823(I2ff115fa483f080d93bada49a9566b33);
            Ibf51e537b992c4b4c0539dda9948f45c    = I12fd829f22ba908180290432320a3660;

            Ibee4f3cd2f516c29ab68e07a640ab65e = Ida03738adc101c03c2229756bed2469d + ~I0b6cdfa1dbfa774fc9a12d856e61cddb + 1;
            I8f967710d03870e026564db0df46d146 = I2bcab411f9bec1541259751bcb9e0823(Ibee4f3cd2f516c29ab68e07a640ab65e);
            I9f83063bdc3c352024f702cb9dc71ce8    = I8f967710d03870e026564db0df46d146;

            Ie495ab560f59ad038992c573de7d2f5b = Ida03738adc101c03c2229756bed2469d + ~I5160de2c5ce4782d8f8be10dc740694b + 1;
            Ia347d80a70a49605c51d19bc2e696aef = I2bcab411f9bec1541259751bcb9e0823(Ie495ab560f59ad038992c573de7d2f5b);
            I72127f6d422ec68dcd47126b87b3d3b1    = Ia347d80a70a49605c51d19bc2e696aef;

            Ibd812def78c3a9c02f9ba45cc0413711 = Ida03738adc101c03c2229756bed2469d + ~I3319313fe1d2b4ec2626711b187b4a5a + 1;
            I730db85d3d11d8327c6d48b8b87a00a4 = I2bcab411f9bec1541259751bcb9e0823(Ibd812def78c3a9c02f9ba45cc0413711);
            I0b4a1b48d110b820d8d87f6e94d32988    = I730db85d3d11d8327c6d48b8b87a00a4;

            I98166634dc80201b0cefb01d9559c228 = Ida03738adc101c03c2229756bed2469d + ~I85dd6a9634284c22027b4241551ea628 + 1;
            I5c6a3ec08cb17d6646bb3e63411a9698 = I2bcab411f9bec1541259751bcb9e0823(I98166634dc80201b0cefb01d9559c228);
            I2e3aeede695007fabe0d6247a93ed403    = I5c6a3ec08cb17d6646bb3e63411a9698;

            Ic2f03a980b5f0b042853ca746abab22b = Ida03738adc101c03c2229756bed2469d + ~I18bb9a781a4c314fe6bd990e4c275f67 + 1;
            I7b5baeec7b11eca457dcd9d2b2b64ac5 = I2bcab411f9bec1541259751bcb9e0823(Ic2f03a980b5f0b042853ca746abab22b);
            I8c5ea3dc59fdcdea1c5f503dde1e815f    = I7b5baeec7b11eca457dcd9d2b2b64ac5;

            I2807a88097d2683ebdb9e0e785e3af02 = I4d14c75f28f3e516c259ea288996131b + ~Idadf072247b351cf51d718f797c3b375 + 1;
            Ic4c7a9d491c560d7b6c410d8216f59bf = I2bcab411f9bec1541259751bcb9e0823(I2807a88097d2683ebdb9e0e785e3af02);
            I873c4dbe95220e40d7388870520261bd    = Ic4c7a9d491c560d7b6c410d8216f59bf;

            I8bebbb3a676c8506af0768516abcd740 = I4d14c75f28f3e516c259ea288996131b + ~If4d63635a5f99c4dc9e5b57712830c20 + 1;
            I2151735079b41a7f8cbfe2b93f1b7470 = I2bcab411f9bec1541259751bcb9e0823(I8bebbb3a676c8506af0768516abcd740);
            I561fa67a9bfbedffcb04e7a4d6b76a64    = I2151735079b41a7f8cbfe2b93f1b7470;

            I31d380f34691c9fe9022035f233b77e2 = I4d14c75f28f3e516c259ea288996131b + ~I75aaeab4f372e28a8e51453540f9c6b2 + 1;
            Ia69e34af60619fa04e8478e2d04768bb = I2bcab411f9bec1541259751bcb9e0823(I31d380f34691c9fe9022035f233b77e2);
            Ia55752d6c4f20378ff570a661ab31d9a    = Ia69e34af60619fa04e8478e2d04768bb;

            I1ffb5675c98ab5b3c62b24eb23441473 = I4d14c75f28f3e516c259ea288996131b + ~I51b1cd475d0e389326b182cbe680a402 + 1;
            I7f9984597d0e7bcda92f13fbb8805687 = I2bcab411f9bec1541259751bcb9e0823(I1ffb5675c98ab5b3c62b24eb23441473);
            Ia13307be43e9155ed0333df62ccc8bf2    = I7f9984597d0e7bcda92f13fbb8805687;

            If56424546ec4f3445853538207ea864e = I4d14c75f28f3e516c259ea288996131b + ~I49d7342f105c4502377abd23db973752 + 1;
            I342ef25fefdb6a326dac80d76052bbd9 = I2bcab411f9bec1541259751bcb9e0823(If56424546ec4f3445853538207ea864e);
            I07b3d1451487a55fbbedda48b0cb6c73    = I342ef25fefdb6a326dac80d76052bbd9;

            I31a49be4a34d9bac2e0d815097439772 = I6e6cbbf430d57f347a0d70558af143d8 + ~I6fcb3b133a6a654b69f41468a713d922 + 1;
            Id1414254ab35ee805c4010432eb24243 = I2bcab411f9bec1541259751bcb9e0823(I31a49be4a34d9bac2e0d815097439772);
            I9f8cf1a6cd0182fba35a49bd232f062a    = Id1414254ab35ee805c4010432eb24243;

            I6b96a2498078953e87de223aa2236d50 = I6e6cbbf430d57f347a0d70558af143d8 + ~I5eaa11e26f19b94dcb7eaee7f09d24b4 + 1;
            I8db7cc6cb4bf55131bee6b00e76baf46 = I2bcab411f9bec1541259751bcb9e0823(I6b96a2498078953e87de223aa2236d50);
            Ie2e488a8589559deeec8598cf6726f1f    = I8db7cc6cb4bf55131bee6b00e76baf46;

            I79bf36e298a85a42c7432f877055f0b4 = I6e6cbbf430d57f347a0d70558af143d8 + ~I586aaa5c55efd37996b01febd3bc60a4 + 1;
            I355aec2468fa96e2f32c8c324c48c5f5 = I2bcab411f9bec1541259751bcb9e0823(I79bf36e298a85a42c7432f877055f0b4);
            I9118ee5ff8c9ba9b125e5baa07bf52e0    = I355aec2468fa96e2f32c8c324c48c5f5;

            I90c070b9bde5da05e8a5d25d2de3ba6b = I6e6cbbf430d57f347a0d70558af143d8 + ~Id5cedaa397ebfc2567efcc2f8a648db5 + 1;
            Ic45ea6e09fd20a2285b7e6e2507910f4 = I2bcab411f9bec1541259751bcb9e0823(I90c070b9bde5da05e8a5d25d2de3ba6b);
            I13b894057e2deae2c00787385de252a8    = Ic45ea6e09fd20a2285b7e6e2507910f4;

            I28d0e4e6d772dd58d845d91952ada300 = I6e6cbbf430d57f347a0d70558af143d8 + ~Ieeb12d463444ca36af1ecf2e09504c06 + 1;
            I288b192ad6d04370df8084511c7f44ce = I2bcab411f9bec1541259751bcb9e0823(I28d0e4e6d772dd58d845d91952ada300);
            I7797a3ea5b97b514a797243cf9fe890a    = I288b192ad6d04370df8084511c7f44ce;

            I7232b4e277acc6f1acefcb606ca24508 = Ib7487df45118e44acec6b9d07bbd5969 + ~I8613cac4ccd4f956e8a0ae7b627f5be2 + 1;
            I4d589e9479ee494636d90a910e530863 = I2bcab411f9bec1541259751bcb9e0823(I7232b4e277acc6f1acefcb606ca24508);
            I3af78697aacc410108d0be7fd13c686b    = I4d589e9479ee494636d90a910e530863;

            I32da124c433c55f692ffa4734d0dc8fc = Ib7487df45118e44acec6b9d07bbd5969 + ~I7d85b73e85379bf3a480e954c05516f3 + 1;
            Ib8fcb6e6569d34c67145861431ad5334 = I2bcab411f9bec1541259751bcb9e0823(I32da124c433c55f692ffa4734d0dc8fc);
            I871cb63247618a543b444aa3f888fffe    = Ib8fcb6e6569d34c67145861431ad5334;

            I56e487db14eeb8d93f494d2f11b57a49 = Ib7487df45118e44acec6b9d07bbd5969 + ~I2266afbacf1ba750ce18f296aba1181d + 1;
            I5405b3c646988338f12191bb8cb02205 = I2bcab411f9bec1541259751bcb9e0823(I56e487db14eeb8d93f494d2f11b57a49);
            I124404013f8fc6b302661900b9ad8ed8    = I5405b3c646988338f12191bb8cb02205;

            I94d3c02bd5b8e84926d4b3c2f56efeac = Ib7487df45118e44acec6b9d07bbd5969 + ~If12366160fdc899bd71cb0de5bcfd84d + 1;
            I371946ff4a809b62ceed2334a9656787 = I2bcab411f9bec1541259751bcb9e0823(I94d3c02bd5b8e84926d4b3c2f56efeac);
            I8e413271c9d13748a1aa2d1a018ff28f    = I371946ff4a809b62ceed2334a9656787;

            I0c35b2e9176f9a06e26ca67d036411b4 = Ib7487df45118e44acec6b9d07bbd5969 + ~I17525df1798fa2c1c4bbc4a1ddcdd0a5 + 1;
            I6d5be8ddd471c1ddf781949169bd9807 = I2bcab411f9bec1541259751bcb9e0823(I0c35b2e9176f9a06e26ca67d036411b4);
            I4d799e93b4dfcabd69977ddb25634a69    = I6d5be8ddd471c1ddf781949169bd9807;

            Ia6ee7b70d0b7fe7c346760b1784e50b9 = I492f382fea500462b3d0866240fb91b2 + ~Ia5c77c9be26d62b026f24ee5a5e25fb8 + 1;
            I499f6bbf3456d23378ff02b6f65a5ae4 = I2bcab411f9bec1541259751bcb9e0823(Ia6ee7b70d0b7fe7c346760b1784e50b9);
            I1487f0027b7d16f4bc85bb00e537cbaf    = I499f6bbf3456d23378ff02b6f65a5ae4;

            I7ce57c278c683ad045526e49bcc47412 = I492f382fea500462b3d0866240fb91b2 + ~Ib5c8d91204a2d313c9c23110a53cd0cf + 1;
            I0c81821914371a777679053e2aa5a55e = I2bcab411f9bec1541259751bcb9e0823(I7ce57c278c683ad045526e49bcc47412);
            I1a5cdaa10022adf0ffbbc0f58b3e690a    = I0c81821914371a777679053e2aa5a55e;

            Ie3d3e681cac0bb919946ac27057409e2 = I492f382fea500462b3d0866240fb91b2 + ~Ife3bb8945e14d8746c82b66886293997 + 1;
            Ief591e9d4759a4b1059574bb624e4ce6 = I2bcab411f9bec1541259751bcb9e0823(Ie3d3e681cac0bb919946ac27057409e2);
            I98246759d003e9bc6676ceb2d093a06b    = Ief591e9d4759a4b1059574bb624e4ce6;

            I8ea0a8cdd6506c982ad75f23136bcebe = I492f382fea500462b3d0866240fb91b2 + ~I887911fd9466f4d4fa7f50642d610d88 + 1;
            Ie40648c85ed87c979a54dfc1f85d1cc8 = I2bcab411f9bec1541259751bcb9e0823(I8ea0a8cdd6506c982ad75f23136bcebe);
            Ia3c2dfb3c4a45091be7cfecfad11f3ec    = Ie40648c85ed87c979a54dfc1f85d1cc8;

            Ic812f8bc775c5ee6a83e2b9aeb22b2a4 = I492f382fea500462b3d0866240fb91b2 + ~I90c44c31fa7903a81826c1c568597362 + 1;
            I36956634f94d6053aa455b29bc0b7a0f = I2bcab411f9bec1541259751bcb9e0823(Ic812f8bc775c5ee6a83e2b9aeb22b2a4);
            I74cda651bcb24472a7697ba017f831a4    = I36956634f94d6053aa455b29bc0b7a0f;

            I0f0adf7fe957b9a68772bd8a1bc163d4 = I3fb3ebddaf28efb56092d19a1b4695de + ~Ic4af6c9097257c9b22a57ce4b79b40fe + 1;
            I05a652e83a9b8c2c38de64de6a70f8bc = I2bcab411f9bec1541259751bcb9e0823(I0f0adf7fe957b9a68772bd8a1bc163d4);
            Id7ba55b14ac0f471142011dc2d57cc4b    = I05a652e83a9b8c2c38de64de6a70f8bc;

            If09562f8d82bc1dea7c38ed51523a889 = I3fb3ebddaf28efb56092d19a1b4695de + ~Ieb7b388ff89e352dd239e0ccbe7b9ecc + 1;
            Iaefa87388884b85eed690e9917bc9d5b = I2bcab411f9bec1541259751bcb9e0823(If09562f8d82bc1dea7c38ed51523a889);
            I5890643c88c4255a0e5efd45f8af3ee2    = Iaefa87388884b85eed690e9917bc9d5b;

            Ib0fd21d66cd89c4e5c95fbc9c7680b62 = I3fb3ebddaf28efb56092d19a1b4695de + ~I89f75107ea95f207b9e664a1f4f0746a + 1;
            I98836c38732b8da439946aa5fcbbd963 = I2bcab411f9bec1541259751bcb9e0823(Ib0fd21d66cd89c4e5c95fbc9c7680b62);
            I4f53e4955e9e506a7169ae810da5dde6    = I98836c38732b8da439946aa5fcbbd963;

            I5a2b2bfadc638fe3fdc31136a8f09a8d = I3fb3ebddaf28efb56092d19a1b4695de + ~I6a86b03402bd2e35208d3fc74601f9cf + 1;
            I8ff116e234a1007cc47989f3fdcf88d6 = I2bcab411f9bec1541259751bcb9e0823(I5a2b2bfadc638fe3fdc31136a8f09a8d);
            Ifc7c1ea337b122fb720767f1890f1a6a    = I8ff116e234a1007cc47989f3fdcf88d6;

            Ica914d8c556285d6b90b35747065a6e5 = I3fb3ebddaf28efb56092d19a1b4695de + ~I3997cf122743b612f49cd5dd125a9201 + 1;
            I53dfee31709f8eca30897d6bf1618418 = I2bcab411f9bec1541259751bcb9e0823(Ica914d8c556285d6b90b35747065a6e5);
            Id40d6f3a8dd09678b25b3e579dd5fb68    = I53dfee31709f8eca30897d6bf1618418;

            I00c5d739bccb0ab6d05da70fe51aafea = I22a26b7f0b1c8c16b00597732ce2ab23 + ~I4a403449a9ba75243369032e1cca1a0d + 1;
            I3ac389b6b81baf93095cc3e9e9c3d8ef = I2bcab411f9bec1541259751bcb9e0823(I00c5d739bccb0ab6d05da70fe51aafea);
            I7002830b0a5f40ba2a2fe7a00c7b6d58    = I3ac389b6b81baf93095cc3e9e9c3d8ef;

            I18e448761bc014ce490b766183350312 = I22a26b7f0b1c8c16b00597732ce2ab23 + ~I886750aaf8d2040c3f12ff113294f658 + 1;
            Ief52e91e9170809b980aa881bf76957a = I2bcab411f9bec1541259751bcb9e0823(I18e448761bc014ce490b766183350312);
            I3f377e8994959ef8182a08538e393d9a    = Ief52e91e9170809b980aa881bf76957a;

            I1b5920f488e9469bd416a6af3072a30b = I22a26b7f0b1c8c16b00597732ce2ab23 + ~I0e52c25aa840402d944cbd81f73c1ffe + 1;
            Iebf813928bcad8ee3b6911057c59752b = I2bcab411f9bec1541259751bcb9e0823(I1b5920f488e9469bd416a6af3072a30b);
            I71bf29f3519e3238cec112ef97ce0579    = Iebf813928bcad8ee3b6911057c59752b;

            I70b41ffed4b6d88ddff219c567b8e968 = I22a26b7f0b1c8c16b00597732ce2ab23 + ~I1112c4267582ddb8148ee40d9529beee + 1;
            I57ae0d331753595cd56d45a28cd5c790 = I2bcab411f9bec1541259751bcb9e0823(I70b41ffed4b6d88ddff219c567b8e968);
            Iaa4bc2f51984f383479b597e6cd4c873    = I57ae0d331753595cd56d45a28cd5c790;

            I935e083b4561da7d015e98ca7f02854e = I2ac08a2d8c917ecb37fbaf5325cb0473 + ~Ic2159627df2efa5e677fa6f4498bdd31 + 1;
            Ibd173152b9400b4c8011451d68b07e4c = I2bcab411f9bec1541259751bcb9e0823(I935e083b4561da7d015e98ca7f02854e);
            I9066a5cf776f80ebf89bdac1f2edb4ac    = Ibd173152b9400b4c8011451d68b07e4c;

            Iaca9ef263bf220d786242b88c994fd21 = I2ac08a2d8c917ecb37fbaf5325cb0473 + ~I58a7c7b05b84d292cd06d68e96ecb9f8 + 1;
            Idc21b018b7b6f2e0bc627e8968e06eda = I2bcab411f9bec1541259751bcb9e0823(Iaca9ef263bf220d786242b88c994fd21);
            I7319203d7231bebb6d6e52422cce5ed2    = Idc21b018b7b6f2e0bc627e8968e06eda;

            I92169291959eb33452b79bfd32618cbc = I2ac08a2d8c917ecb37fbaf5325cb0473 + ~I20c4e393929b875521e5316f4d8e2d42 + 1;
            I783423950d0e0229826b2249f5cfdf5c = I2bcab411f9bec1541259751bcb9e0823(I92169291959eb33452b79bfd32618cbc);
            I4e8309976fd6011d78728cef935dc3c1    = I783423950d0e0229826b2249f5cfdf5c;

            I126dabc3ebb9c4157adf62b57f217bd0 = I2ac08a2d8c917ecb37fbaf5325cb0473 + ~I21c207af859b94634d3750482b42a2ca + 1;
            I6b8fc6d29fb4549e3f191f913bccff9e = I2bcab411f9bec1541259751bcb9e0823(I126dabc3ebb9c4157adf62b57f217bd0);
            I5ed502118c175d5bdb4607973554a3a3    = I6b8fc6d29fb4549e3f191f913bccff9e;

            If4433b1ef2eb963cd301946958b69884 = I50ff8f51e75fb9ce3db983c2a0f57196 + ~Id5b4ee69444e5b499476c05a7f1d6e60 + 1;
            Idc98380b110c22495027a7cdb6f2029d = I2bcab411f9bec1541259751bcb9e0823(If4433b1ef2eb963cd301946958b69884);
            If457f80b3d29b60b840f886fa928297c    = Idc98380b110c22495027a7cdb6f2029d;

            I67ac5b9b794787b3c4738c3366689871 = I50ff8f51e75fb9ce3db983c2a0f57196 + ~Ia308e09137af1cb50167562efb5da628 + 1;
            Ieb72df81e325eda4d80a237454fa9dbd = I2bcab411f9bec1541259751bcb9e0823(I67ac5b9b794787b3c4738c3366689871);
            I7e0f785ec7554540c9a4a413a3afa75f    = Ieb72df81e325eda4d80a237454fa9dbd;

            I4f022d70078c412bdbef158f750d3da3 = I50ff8f51e75fb9ce3db983c2a0f57196 + ~I2418ae211f327ed45cc70c42078180dc + 1;
            If70e7ed8d4989cd75d37af1dc5d185ed = I2bcab411f9bec1541259751bcb9e0823(I4f022d70078c412bdbef158f750d3da3);
            Id3662bbe1b5191995d1656045fe6b6a6    = If70e7ed8d4989cd75d37af1dc5d185ed;

            I6be6165385f6a77aeedb88f2baaa9cab = I50ff8f51e75fb9ce3db983c2a0f57196 + ~I2ff2421bd86bf9ec110724460f1171e9 + 1;
            Ifc99661bc592c2c43bae53db10c8d472 = I2bcab411f9bec1541259751bcb9e0823(I6be6165385f6a77aeedb88f2baaa9cab);
            Idf922fab93bc2357ac1f66f73f3ead0b    = Ifc99661bc592c2c43bae53db10c8d472;

            Id1f7fe91547e158e1d39edffb1421ff3 = I444bc340ffb7ef7b72d4d2e761d58872 + ~I48b39ee498563e23c3a4be079b6100d8 + 1;
            Ic8860cc8d323e5a4c68233109ed70512 = I2bcab411f9bec1541259751bcb9e0823(Id1f7fe91547e158e1d39edffb1421ff3);
            I780371393ef898aa144c5bc36e74c654    = Ic8860cc8d323e5a4c68233109ed70512;

            I7a51924134902612db53941390891245 = I444bc340ffb7ef7b72d4d2e761d58872 + ~Iddf65ccb4396288264a400ba37cbb655 + 1;
            I439288f09536ca87fa0feb5f6436716e = I2bcab411f9bec1541259751bcb9e0823(I7a51924134902612db53941390891245);
            I79696cd10cffa4c0181a2089da6b3262    = I439288f09536ca87fa0feb5f6436716e;

            I45128b9e29dd2fdd94a78fc5ffdff2b1 = I444bc340ffb7ef7b72d4d2e761d58872 + ~If29fcea810adbdb1c4d8a4ace1d8081b + 1;
            I66c4beb8fe2d9f363c8e153a12f216ca = I2bcab411f9bec1541259751bcb9e0823(I45128b9e29dd2fdd94a78fc5ffdff2b1);
            I073155ab0359a13b77f730653dcfc08d    = I66c4beb8fe2d9f363c8e153a12f216ca;

            I7f1082408c8ebb5be18e8f71ff9510e5 = I444bc340ffb7ef7b72d4d2e761d58872 + ~I6ba5c453b17e4b33c61caf5d70041c4a + 1;
            Ib2a96d55b1f7bf9b89286de32e59fad3 = I2bcab411f9bec1541259751bcb9e0823(I7f1082408c8ebb5be18e8f71ff9510e5);
            I1b44f781d81438654f69bb7fbdb94011    = Ib2a96d55b1f7bf9b89286de32e59fad3;

            I655ebf19c2f4b3dde716668f9ce12e59 = I039c6cac5830759529595a958b7f65c9 + ~Iac8cb32c2d86b975f51a2ed605002e51 + 1;
            I3028dabd706c9e5768eac56c66463955 = I2bcab411f9bec1541259751bcb9e0823(I655ebf19c2f4b3dde716668f9ce12e59);
            Id68f1a0ec8ff80da3190fe517bd935e3    = I3028dabd706c9e5768eac56c66463955;

            Ibc9d493a507122d92af42d858cdc4c61 = I039c6cac5830759529595a958b7f65c9 + ~I88a325547ccfe4eabf90792abd60e356 + 1;
            I265f3da3571d2ddb786b98ba3959823b = I2bcab411f9bec1541259751bcb9e0823(Ibc9d493a507122d92af42d858cdc4c61);
            I3704464d41956032b779eebe27511815    = I265f3da3571d2ddb786b98ba3959823b;

            Ib3d3103e5ee4feb160a97c7e26f7102b = I039c6cac5830759529595a958b7f65c9 + ~I0722ec4e9d400f8eaeacd060e42de79c + 1;
            If8d81c152d863660081339144b37a052 = I2bcab411f9bec1541259751bcb9e0823(Ib3d3103e5ee4feb160a97c7e26f7102b);
            Ie6756ee9631791940ffc6fddb223b4d0    = If8d81c152d863660081339144b37a052;

            I6cc56b119e72175df3b7ce64dc3d9305 = I039c6cac5830759529595a958b7f65c9 + ~I08318099725fbe033ab8d5427eb8b278 + 1;
            Ie9cba6422546d378655d0ef98ef974fb = I2bcab411f9bec1541259751bcb9e0823(I6cc56b119e72175df3b7ce64dc3d9305);
            I085151dfc2e773a7a485f5ef1b7cd6bd    = Ie9cba6422546d378655d0ef98ef974fb;

            I57cf4a9378f1cdd94a1a5608dc57e05f = I0584de7d919236ab138e288a27d08ff1 + ~If85d9a95c1c02ce2da1dc3486b53eb81 + 1;
            Iaddf6de71a6329eb536f54e3d18d43d6 = I2bcab411f9bec1541259751bcb9e0823(I57cf4a9378f1cdd94a1a5608dc57e05f);
            I2654e83fff153df7760c341f59a23396    = Iaddf6de71a6329eb536f54e3d18d43d6;

            I4160ab1aa18e8151c0a5c23b9edeb907 = I0584de7d919236ab138e288a27d08ff1 + ~Iae21bdea20a6266d3f69aa680b6b2817 + 1;
            I280ed7bf157554fcad915f0e7fa12653 = I2bcab411f9bec1541259751bcb9e0823(I4160ab1aa18e8151c0a5c23b9edeb907);
            Iee3eec7a9d7a3a5c22281545ec143e50    = I280ed7bf157554fcad915f0e7fa12653;

            Ia1f183f2d904d006e46399424e06c614 = I0584de7d919236ab138e288a27d08ff1 + ~Ic6a7a82d16e6106071934ba79d3698cd + 1;
            I0ca797b233dcdac8e390e1e41d99b196 = I2bcab411f9bec1541259751bcb9e0823(Ia1f183f2d904d006e46399424e06c614);
            Ied2b9ca07a6d498abada30fb0726df24    = I0ca797b233dcdac8e390e1e41d99b196;

            If979702738671323995e56108bc9376c = I0584de7d919236ab138e288a27d08ff1 + ~If36cb462cdf20b0b1758cd6417e524fa + 1;
            I150792edd72cc07cf8242d787cb52056 = I2bcab411f9bec1541259751bcb9e0823(If979702738671323995e56108bc9376c);
            If95315702519e7a08386a870e599aab0    = I150792edd72cc07cf8242d787cb52056;

            Ibc96fe0a6bf1f95036f97c7d44fab575 = I086402c82ec67ae09a9e6360c58904b4 + ~I59fba74472ded0a985cb237104ac127f + 1;
            I186c13747ff5a1ee6e562ad9e5faabd9 = I2bcab411f9bec1541259751bcb9e0823(Ibc96fe0a6bf1f95036f97c7d44fab575);
            I1091064aef7d915ba8fb6cbded069102    = I186c13747ff5a1ee6e562ad9e5faabd9;

            I755a38220a693ba43701d30e7e9508ad = I086402c82ec67ae09a9e6360c58904b4 + ~I77e1f5f504a794edbb89c66cf1ffcf66 + 1;
            I6fb8240f8c68b71cafe4c2c43ac7db33 = I2bcab411f9bec1541259751bcb9e0823(I755a38220a693ba43701d30e7e9508ad);
            I40685c7d2c8be12698f734ec6213b5b4    = I6fb8240f8c68b71cafe4c2c43ac7db33;

            I896fb82baa9647a14f4b5b1ecfa70a15 = I086402c82ec67ae09a9e6360c58904b4 + ~I3cc30aaba3dcd3eda262a19e85e53117 + 1;
            I166f5cab59c2a66117f2287d2b11c096 = I2bcab411f9bec1541259751bcb9e0823(I896fb82baa9647a14f4b5b1ecfa70a15);
            Icc7775fe34c162006b93662530fd4944    = I166f5cab59c2a66117f2287d2b11c096;

            I23d1c973d7a2048353fbb68e4a294c08 = I086402c82ec67ae09a9e6360c58904b4 + ~I40e8463645b1122b7cb224770fa00447 + 1;
            Ie896986a747c1cd8ccad7117125c6e0d = I2bcab411f9bec1541259751bcb9e0823(I23d1c973d7a2048353fbb68e4a294c08);
            I2e6f1a5695ad23b8ca282b344832ee8e    = Ie896986a747c1cd8ccad7117125c6e0d;

            If9fd1e08af14f2fd4ca363383f48580a = I1cefdc831c146187c77f861b3e2d1af0 + ~Id6105518ade80c89d4f20222a2382efb + 1;
            I0c829f14ef188ff7ae1417e28903f2b3 = I2bcab411f9bec1541259751bcb9e0823(If9fd1e08af14f2fd4ca363383f48580a);
            I016ce894bebdaa7e56af9deb1ccfb3f5    = I0c829f14ef188ff7ae1417e28903f2b3;

            I8f3782f78d88a5c3bc93709564999b30 = I1cefdc831c146187c77f861b3e2d1af0 + ~I8493e2dac01f009db1d2d5504b49d135 + 1;
            I3591d4f320f8401ef8ad8f92d2d89bf6 = I2bcab411f9bec1541259751bcb9e0823(I8f3782f78d88a5c3bc93709564999b30);
            Iad2dd0815c1107160992e5070632f76c    = I3591d4f320f8401ef8ad8f92d2d89bf6;

            I986d61d79ce31f4677f3293339db6ad2 = I1cefdc831c146187c77f861b3e2d1af0 + ~I106d0e71b7378d110b0a624e5cbf0d6e + 1;
            I3816895f23a1381e42aaeb64dd158fda = I2bcab411f9bec1541259751bcb9e0823(I986d61d79ce31f4677f3293339db6ad2);
            Iefaba2acd282081b9a0a98ed057ca85e    = I3816895f23a1381e42aaeb64dd158fda;

            Ica4d93d9fad21316002008ade5106a9d = I1cefdc831c146187c77f861b3e2d1af0 + ~Ide386e751e06dd5df0c042cd76f0f800 + 1;
            Ic9c34a36b2fde9649064680904ec9150 = I2bcab411f9bec1541259751bcb9e0823(Ica4d93d9fad21316002008ade5106a9d);
            Id4ef94eb8d5db8810bca4c9d669f0b7f    = Ic9c34a36b2fde9649064680904ec9150;

            If77592d5d8bed32477fd690341e543d0 = Ida9c16ae57d17b6faee8a54838860447 + ~I185085cbf8da6df921ba32442b28bcca + 1;
            If7eb75eccc5a6384c80d99b64d534fca = I2bcab411f9bec1541259751bcb9e0823(If77592d5d8bed32477fd690341e543d0);
            I04e845e6a5ed71978b636593dd749b12    = If7eb75eccc5a6384c80d99b64d534fca;

            I25b70c6b830cbfe1b41d8f289c751924 = Ida9c16ae57d17b6faee8a54838860447 + ~Iaf3a0b5ea5d9eda47fcced9260922bc6 + 1;
            Ib788a897a1d1b86b2c16caade11846ee = I2bcab411f9bec1541259751bcb9e0823(I25b70c6b830cbfe1b41d8f289c751924);
            I0b2760b437be2cb79382f8d6a7b8969e    = Ib788a897a1d1b86b2c16caade11846ee;

            I2a5d65eeffa18dd9af9fe36463dafd7c = Ida9c16ae57d17b6faee8a54838860447 + ~Ic8f0049e1298b14b4e039075dc0d5f74 + 1;
            I6a5fec9dad124f6d8c5574bcc2643ede = I2bcab411f9bec1541259751bcb9e0823(I2a5d65eeffa18dd9af9fe36463dafd7c);
            I1b0fdaeebe5fee6fbb2e13aac5e233a1    = I6a5fec9dad124f6d8c5574bcc2643ede;

            Ibafa6e10bd4edf5d224fdeb2f9adbf98 = Ida9c16ae57d17b6faee8a54838860447 + ~If63bb4681bf1116c0d1db3aa21bf52ac + 1;
            I3936f324b08bea1bc5f8bcd12437b161 = I2bcab411f9bec1541259751bcb9e0823(Ibafa6e10bd4edf5d224fdeb2f9adbf98);
            Iee872d17e4a28075be0ad7086c3acc91    = I3936f324b08bea1bc5f8bcd12437b161;

            Ifc25402bd879bc5c43b4945b60cd4540 = Ia3b9fb112f39dd0ccbf7555659369efb + ~I5c278aad08b7c4b0237d68f88fcb3f3a + 1;
            I1a59337d4da3e3ad1a738a9c3b56ef8c = I2bcab411f9bec1541259751bcb9e0823(Ifc25402bd879bc5c43b4945b60cd4540);
            I87656ddd4ef8f1ae36c7566d5e7892d8    = I1a59337d4da3e3ad1a738a9c3b56ef8c;

            Iec48da6882325d8a33e0e0e845eb18a0 = Ia3b9fb112f39dd0ccbf7555659369efb + ~I9222c4c0eb2b110fd80547d46ba17036 + 1;
            Ic3e3b4cba05d80c0ceaa6e25a906a602 = I2bcab411f9bec1541259751bcb9e0823(Iec48da6882325d8a33e0e0e845eb18a0);
            I865cd0535644db7f17db1180c85f1744    = Ic3e3b4cba05d80c0ceaa6e25a906a602;

            I0fd05e46862fdf8e614afaa3fd478602 = Ia3b9fb112f39dd0ccbf7555659369efb + ~I95ccc219b5f5038641b38dff6db0b222 + 1;
            Ife0830e12b8bbb5aa0b8c2c0e4191e59 = I2bcab411f9bec1541259751bcb9e0823(I0fd05e46862fdf8e614afaa3fd478602);
            I71d46741fa94df65e1bdf6abff53d2ba    = Ife0830e12b8bbb5aa0b8c2c0e4191e59;

            I6253a59dca81842d9ab6e58cf204abbf = Ia3b9fb112f39dd0ccbf7555659369efb + ~I566c72342c69969892480fae41232c37 + 1;
            I95eaa4ac5199ebbb06f780d1376062ec = I2bcab411f9bec1541259751bcb9e0823(I6253a59dca81842d9ab6e58cf204abbf);
            Ic223d7941250d739ce9bb0ae5013646e    = I95eaa4ac5199ebbb06f780d1376062ec;

            Ib18d64bc58b354358ee6ac16785880e2 = Ib1bfcdc0c972aafc99116ed8c0511445 + ~I21842d06e25948ef461d1fd03485f86c + 1;
            Ib40ccfdb9ea28f333a7cc67f2446c923 = I2bcab411f9bec1541259751bcb9e0823(Ib18d64bc58b354358ee6ac16785880e2);
            I1ef9b548b943a1f2012b91c7e0b445f2    = Ib40ccfdb9ea28f333a7cc67f2446c923;

            I28689b693a7a5f761a1f252aa3ef3b67 = Ib1bfcdc0c972aafc99116ed8c0511445 + ~Ib2c1636a66f6479d6123a038cbc668d5 + 1;
            I507515355429e697cd5496809aa03cfb = I2bcab411f9bec1541259751bcb9e0823(I28689b693a7a5f761a1f252aa3ef3b67);
            I88b6d7894d82ff394e89c7471c80dd5b    = I507515355429e697cd5496809aa03cfb;

            I1a4e6d12f9776d5e61094e0b5edf71d9 = Ib1bfcdc0c972aafc99116ed8c0511445 + ~I69c2b063e61e14f5d49b907095ece00f + 1;
            I6bcc3a323e67f95eb4bf28a0704d3c50 = I2bcab411f9bec1541259751bcb9e0823(I1a4e6d12f9776d5e61094e0b5edf71d9);
            Ia5fc7e1f991f30042b848888a546534b    = I6bcc3a323e67f95eb4bf28a0704d3c50;

            I8e1ad23b7ac662bb827a83d3709f0adb = Ib1bfcdc0c972aafc99116ed8c0511445 + ~Ia0f7deea6b1ce1050dcf97fa99de9178 + 1;
            I55e3a2566ef3ac257021a294376be634 = I2bcab411f9bec1541259751bcb9e0823(I8e1ad23b7ac662bb827a83d3709f0adb);
            If699df4c8261ebce5c5d1aebe062cd61    = I55e3a2566ef3ac257021a294376be634;

            I000ad2287813072cc18dad933758f2ab = I7adff505c50450a04f1717cac1adebe7 + ~I37e360420c7dd061de93a6647513676d + 1;
            I40f10dc3289ea8a59f593f62066aaff8 = I2bcab411f9bec1541259751bcb9e0823(I000ad2287813072cc18dad933758f2ab);
            I19338369553e96bb2476d80fe84dec3e    = I40f10dc3289ea8a59f593f62066aaff8;

            I7bc3698b51b89ac38ba5f4b5428a0c96 = I7adff505c50450a04f1717cac1adebe7 + ~I535b29f7177b4fc009ee998f1f4f7d7f + 1;
            Ieeabde5600d81208346ebd50d4a95d83 = I2bcab411f9bec1541259751bcb9e0823(I7bc3698b51b89ac38ba5f4b5428a0c96);
            I9844ff02042cbc04dd5f4179908bbb2d    = Ieeabde5600d81208346ebd50d4a95d83;

            I78aea1705621e2845a331c3e61a8055b = I7adff505c50450a04f1717cac1adebe7 + ~I45ef0ac486fe043f57e8a46aa91461a3 + 1;
            Ibb9220dcdd6d7fc2b6d6ca5f4cc93a8b = I2bcab411f9bec1541259751bcb9e0823(I78aea1705621e2845a331c3e61a8055b);
            I89cc6a060b714985b24f724adc782e7b    = Ibb9220dcdd6d7fc2b6d6ca5f4cc93a8b;

            I0a31314c3580f5f9e61e79c133e5d794 = I7adff505c50450a04f1717cac1adebe7 + ~I992b9876530d53c1b62d98511bf41942 + 1;
            I05a3aebc90966144a6809e460d6ceda1 = I2bcab411f9bec1541259751bcb9e0823(I0a31314c3580f5f9e61e79c133e5d794);
            I39d94ce7fbe37a74404e0043060441ed    = I05a3aebc90966144a6809e460d6ceda1;

            I0e274fd7bfc0388fef95a8ceb939ee91 = I699feb4382974a02b21cb387c13f7f3f + ~I8e470b68bf35c647af42b6e46201e570 + 1;
            I7e3150622eb318e94f99b36016ac7d2f = I2bcab411f9bec1541259751bcb9e0823(I0e274fd7bfc0388fef95a8ceb939ee91);
            I0a1c9a8d59dbcffd6847f3a65107c407    = I7e3150622eb318e94f99b36016ac7d2f;

            Id6f39ddcb73d3f4ec081a365d11d1ef4 = I699feb4382974a02b21cb387c13f7f3f + ~I8cbafa797ef136d7e50c909dc160deb1 + 1;
            Ifb146b2073d447377a1b21fe21baa4da = I2bcab411f9bec1541259751bcb9e0823(Id6f39ddcb73d3f4ec081a365d11d1ef4);
            I2328556c467a9e639f2b6ba1d0cb99b7    = Ifb146b2073d447377a1b21fe21baa4da;

            I807770bfa86d160459d6ec3c0f4d6a0b = I699feb4382974a02b21cb387c13f7f3f + ~I850c257a0412bd9bd6001817bd9d0ee1 + 1;
            Ifa5048ac43025e9cdf3f3436c37bb835 = I2bcab411f9bec1541259751bcb9e0823(I807770bfa86d160459d6ec3c0f4d6a0b);
            I5c9d75d6431d69db1abe412e591000a7    = Ifa5048ac43025e9cdf3f3436c37bb835;

            I31c89b8a11a3090bfd74b112cbc474bb = I699feb4382974a02b21cb387c13f7f3f + ~Ib8861f627f6273c0a031bf43e7812a5d + 1;
            I837ba4049e4973924e51d642f7f481ad = I2bcab411f9bec1541259751bcb9e0823(I31c89b8a11a3090bfd74b112cbc474bb);
            I8dc3dcdefc85b6ff8ecfa09cfc7e69fa    = I837ba4049e4973924e51d642f7f481ad;

            I79b82cb1bfc72bd5a9d313b9e9c9203c = Idc99c3b23e49aca3c98f0685ea34441c + ~Ia526539cc0f844b802d412b7a17cb6a6 + 1;
            I2910e5e74ca008b7e5502d787cb88a6d = I2bcab411f9bec1541259751bcb9e0823(I79b82cb1bfc72bd5a9d313b9e9c9203c);
            I69f6c909ea6b207c200b154e00e13a05    = I2910e5e74ca008b7e5502d787cb88a6d;

            Ib1046ae03c9a77fd2c0b3e9838e9af87 = Idc99c3b23e49aca3c98f0685ea34441c + ~I71bc7271cc432bb3c5d0b7a416cdfc60 + 1;
            Ia24816d601e29172628cad0c364b47e9 = I2bcab411f9bec1541259751bcb9e0823(Ib1046ae03c9a77fd2c0b3e9838e9af87);
            Id365c9f8f7f97c777bd5da0ce9490511    = Ia24816d601e29172628cad0c364b47e9;

            Ic63723fd43cbbbde51c233a3cca15d3f = Idc99c3b23e49aca3c98f0685ea34441c + ~I12e8b8cf609c2fbdc72efce9bb5dabee + 1;
            I8f99af880f329241cfc9616ff9859091 = I2bcab411f9bec1541259751bcb9e0823(Ic63723fd43cbbbde51c233a3cca15d3f);
            Idf0206d2ad2bdef7db1d30a2d715cc6a    = I8f99af880f329241cfc9616ff9859091;

            I3abbb59abada1aec6941185f95f738bd = Idc99c3b23e49aca3c98f0685ea34441c + ~Ieb5bac4ef0f5e4e0b826cdc43ae71471 + 1;
            Iea7c2970a7d80c55c1a6d6933c6c81c9 = I2bcab411f9bec1541259751bcb9e0823(I3abbb59abada1aec6941185f95f738bd);
            I07d1c54431eed887554a136f15f86d22    = Iea7c2970a7d80c55c1a6d6933c6c81c9;

            I8d5bd7039a77ce82ce0f6cbba9c2a076 = Ib67318fa6954ec8f3247927d34e74f8c + ~I26cf25e680483bf4e556d74efec35ee7 + 1;
            I75a12697a4ee6de46fc098b0f02b8349 = I2bcab411f9bec1541259751bcb9e0823(I8d5bd7039a77ce82ce0f6cbba9c2a076);
            Ic16809a3c82787ed88819fc9e9613f85    = I75a12697a4ee6de46fc098b0f02b8349;

            I527ad0b9382dd7b6e657dc1a32d8e472 = Ib67318fa6954ec8f3247927d34e74f8c + ~I9cbe73d708c561d43d05945552d32dde + 1;
            I623d1f0b6829caf5dc0f0eab0ca47f74 = I2bcab411f9bec1541259751bcb9e0823(I527ad0b9382dd7b6e657dc1a32d8e472);
            I1613ae89442495e703a52e65b8a0bf9f    = I623d1f0b6829caf5dc0f0eab0ca47f74;

            I8de02f32e14e719f4930d99743c04a20 = Ib67318fa6954ec8f3247927d34e74f8c + ~Ieb9720b6beb2363d651346ef0233cd49 + 1;
            Ieabf207f10f7df1e9059f1e953d7b399 = I2bcab411f9bec1541259751bcb9e0823(I8de02f32e14e719f4930d99743c04a20);
            I6089da825af433e847c0b1bb9ff7d373    = Ieabf207f10f7df1e9059f1e953d7b399;

            I7614dd5e9628c761dd9b2a512cb1da98 = Ib67318fa6954ec8f3247927d34e74f8c + ~I3cd0883d9f0ba7475f474f1e318ef023 + 1;
            I1399b55530e343bd85606e7c7529d453 = I2bcab411f9bec1541259751bcb9e0823(I7614dd5e9628c761dd9b2a512cb1da98);
            I6aa7fccf4e225fa70063fd24dab74e6b    = I1399b55530e343bd85606e7c7529d453;

            Icae7efa4742dd0ad943ee1f67b0c9b14 = I8774ce3f11362915c4331d1026e452dd + ~Ic989dc794ce4356856b3916ab1889589 + 1;
            I39ee898ed8a8af64552e1aa145437310 = I2bcab411f9bec1541259751bcb9e0823(Icae7efa4742dd0ad943ee1f67b0c9b14);
            Ibe2a5f680405f233256b6fd806b72ae5    = I39ee898ed8a8af64552e1aa145437310;

            Ieb1854b79e9a2bc6cf5aa1c319e8e753 = I8774ce3f11362915c4331d1026e452dd + ~I82a225237aeb1ceb31e8cd18b1e45c6f + 1;
            I0af241f9f65af3bff2bb0d69977bb0c6 = I2bcab411f9bec1541259751bcb9e0823(Ieb1854b79e9a2bc6cf5aa1c319e8e753);
            I662d408ffd8fb9f249e531a167161429    = I0af241f9f65af3bff2bb0d69977bb0c6;

            Iff50b77f300183ca59a67ccbcc9573c4 = I8774ce3f11362915c4331d1026e452dd + ~I2ea27544ba4cc14d0f7ccf7158a27a2f + 1;
            I9de68705b5430023d2eb5554370bb188 = I2bcab411f9bec1541259751bcb9e0823(Iff50b77f300183ca59a67ccbcc9573c4);
            Ie95b8a5c2da6c0877d49c646c194f5b7    = I9de68705b5430023d2eb5554370bb188;

            I4868604f8178663de759d4c63dc6c4bd = I8774ce3f11362915c4331d1026e452dd + ~I5f8a41ab83a9257e534973e981e28e9b + 1;
            Icdf7ba01c4813abe3cfa760f2d8d5c84 = I2bcab411f9bec1541259751bcb9e0823(I4868604f8178663de759d4c63dc6c4bd);
            If940f33461f5e297e158db54f6aad610    = Icdf7ba01c4813abe3cfa760f2d8d5c84;

            Ife992a151986c58df4cba79b6bc4ac0a = I2392b2d17ffed6073875fbe8e92534cf + ~Ibcb80df5bed66f8498561e3f3ffa4ec4 + 1;
            Ia6b995eb6bbaad8a638c80d587d45ab9 = I2bcab411f9bec1541259751bcb9e0823(Ife992a151986c58df4cba79b6bc4ac0a);
            I54aa9d4c6333d94970eae97aeb3603fa    = Ia6b995eb6bbaad8a638c80d587d45ab9;

            I9ab973fb74d9fac5d78eb8fc2c7ecf36 = I2392b2d17ffed6073875fbe8e92534cf + ~Ib7fde6a2ec1ff0a3af10bccf3012e63f + 1;
            I75c2987dcebc9cdca578aeebec96fccc = I2bcab411f9bec1541259751bcb9e0823(I9ab973fb74d9fac5d78eb8fc2c7ecf36);
            Ib82fc62720e6346e1c05cc33d596447e    = I75c2987dcebc9cdca578aeebec96fccc;

            I5ee7916e859b86a98538659401685016 = I2392b2d17ffed6073875fbe8e92534cf + ~I0e420136675d5f0d1aa027d589ee8741 + 1;
            I6fab90e9a0f606d7c26346c89c6f1d47 = I2bcab411f9bec1541259751bcb9e0823(I5ee7916e859b86a98538659401685016);
            I24873624848b61f313865e10e77e35c6    = I6fab90e9a0f606d7c26346c89c6f1d47;

            I48c284cefb8cfb5a938a8f23ce4d7f03 = I3a4f0d3e32596ef05477f494768d4266 + ~Iba75ff0f3b67c7e28cf627706733d528 + 1;
            Iab2f70a1d3093b3194e9047a8fe8e487 = I2bcab411f9bec1541259751bcb9e0823(I48c284cefb8cfb5a938a8f23ce4d7f03);
            Icc3915d8325c22fc172f731553798fef    = Iab2f70a1d3093b3194e9047a8fe8e487;

            I5c1fc666b77a689478654dd29519f458 = I3a4f0d3e32596ef05477f494768d4266 + ~I4854ff71aa885da3d07acaaa24740d7c + 1;
            Ic84b6224be8eb8eefc9ad9bcc2280291 = I2bcab411f9bec1541259751bcb9e0823(I5c1fc666b77a689478654dd29519f458);
            I93b9837e63103431a0fdaf319a465c90    = Ic84b6224be8eb8eefc9ad9bcc2280291;

            I38bba98b59184c75ba3b27e1dcf52182 = I3a4f0d3e32596ef05477f494768d4266 + ~I4aab6ff52e3fba90bb7417cb50766125 + 1;
            I64a0e60fdcc93d84606774196b2b7598 = I2bcab411f9bec1541259751bcb9e0823(I38bba98b59184c75ba3b27e1dcf52182);
            I91237af3aa2af551dbbc626bb701215e    = I64a0e60fdcc93d84606774196b2b7598;

            I6905b65403c16b0211643227ece536f6 = Icd08ff59cf6be3ba97698dd55703339e + ~Id65f22fa8fc9c47bfd00c796b63c9fa4 + 1;
            Iaa6a4f3826d87e43dd3213dc5083184b = I2bcab411f9bec1541259751bcb9e0823(I6905b65403c16b0211643227ece536f6);
            Ib254d9701567f642d3586641edf85128    = Iaa6a4f3826d87e43dd3213dc5083184b;

            I3ed34401bba9d5f229bc98480aedd9a5 = Icd08ff59cf6be3ba97698dd55703339e + ~If7543e2f5a158b1f3f3a4078ec54cab5 + 1;
            I94fd5b790a9dceab1b4b3f1b5e30a0d9 = I2bcab411f9bec1541259751bcb9e0823(I3ed34401bba9d5f229bc98480aedd9a5);
            I25c50067a62d2b3599d15f12f89d384e    = I94fd5b790a9dceab1b4b3f1b5e30a0d9;

            Ib4d05804277cddc7f00ac17ac14f5325 = Icd08ff59cf6be3ba97698dd55703339e + ~I1ba7f209cb735471073e8051026a148c + 1;
            I9c8c1d22021bbe798b1863ae1dfc3965 = I2bcab411f9bec1541259751bcb9e0823(Ib4d05804277cddc7f00ac17ac14f5325);
            I238be7f0e4a209a6b4201a024c8aed82    = I9c8c1d22021bbe798b1863ae1dfc3965;

            I41babdca6d3fa462849592d37b0a7998 = I985fb7ed22a8476ea322c9e3c2b3851c + ~Ia81c31ea4f4786136b539c9766987596 + 1;
            I870366e9c3b29c1683a7528f4b5d5329 = I2bcab411f9bec1541259751bcb9e0823(I41babdca6d3fa462849592d37b0a7998);
            I233f5ddadd45c0df2108ea6c1d634f3c    = I870366e9c3b29c1683a7528f4b5d5329;

            I58cfec706dc929ebfdeaca6e01b00c0a = I985fb7ed22a8476ea322c9e3c2b3851c + ~I6a3824a6598bbaa138e1e763ad85f5f7 + 1;
            I066db3b79f8b4581f96567d943a7e7db = I2bcab411f9bec1541259751bcb9e0823(I58cfec706dc929ebfdeaca6e01b00c0a);
            I87a320ddaa1478146ff6e519dc65c40a    = I066db3b79f8b4581f96567d943a7e7db;

            I7efe3c5b2fc69840a79545e0399ce749 = I985fb7ed22a8476ea322c9e3c2b3851c + ~I711c5cf9fd8c5161bac36060b3443503 + 1;
            Iabd6f58c4760c939dfd58e4f426bcab9 = I2bcab411f9bec1541259751bcb9e0823(I7efe3c5b2fc69840a79545e0399ce749);
            Ibf03d6940c0a38bef038a28b6a7b625d    = Iabd6f58c4760c939dfd58e4f426bcab9;

            I70e3eeb2b3966676d16a6aa4c85753ab = Ib985709316b1b0a9d3fa3c1eaf6c641f + ~Ie380b37a78242e6d45b659d568887457 + 1;
            Ia3505661cb9b7eacbd47774346d12f5b = I2bcab411f9bec1541259751bcb9e0823(I70e3eeb2b3966676d16a6aa4c85753ab);
            I90942470e2057e50ce4f5745ed68b81c    = Ia3505661cb9b7eacbd47774346d12f5b;

            I2a32d545d1e7beecc7531174c7e8dfbc = Ib985709316b1b0a9d3fa3c1eaf6c641f + ~I72108531a608f6d5e51a481c68d7b271 + 1;
            I4e7245fc882e3e284d8c152c8998b028 = I2bcab411f9bec1541259751bcb9e0823(I2a32d545d1e7beecc7531174c7e8dfbc);
            I77fbc3f3b65962b610e39f4b085ecb7e    = I4e7245fc882e3e284d8c152c8998b028;

            Ib8fb40e4ba0ba1f5e9f5a99d1271ed06 = Ib985709316b1b0a9d3fa3c1eaf6c641f + ~Ic9740baafb1c92e3a25f0a1e7bc46486 + 1;
            Ibe962754759204890883a6de0993a64b = I2bcab411f9bec1541259751bcb9e0823(Ib8fb40e4ba0ba1f5e9f5a99d1271ed06);
            I701845efaf1b02aefa381d4f6b45c401    = Ibe962754759204890883a6de0993a64b;

            Ica792cb9850a61fa4a8bd8a4b6c6ca05 = Ib985709316b1b0a9d3fa3c1eaf6c641f + ~Ie3591b22e0e127f04658da68d4846be9 + 1;
            Id2ef1e193163adc702763541f37fec4d = I2bcab411f9bec1541259751bcb9e0823(Ica792cb9850a61fa4a8bd8a4b6c6ca05);
            Id446ddfd713c6e1592c562cfb123ea8b    = Id2ef1e193163adc702763541f37fec4d;

            I779e5997c66649d6d54fd7f0514c47bd = I4be898887dff6e2cebe53f135ece131b + ~I484ec87270fcc959a486ebce40a9a03c + 1;
            I8a925721cf106d4e6ca1f69bbc2f53d4 = I2bcab411f9bec1541259751bcb9e0823(I779e5997c66649d6d54fd7f0514c47bd);
            If4f752779d27392e7536565d425bce25    = I8a925721cf106d4e6ca1f69bbc2f53d4;

            I5aa578b0c2831453683fa44af1878cb8 = I4be898887dff6e2cebe53f135ece131b + ~Ibdd9957b7f1a319b797c021933ff75d7 + 1;
            Ib97671e4daa1b606aa01c5e8f753a9e8 = I2bcab411f9bec1541259751bcb9e0823(I5aa578b0c2831453683fa44af1878cb8);
            If112169057d6293326a56443ac3cf517    = Ib97671e4daa1b606aa01c5e8f753a9e8;

            I735d6229ef1a4ecda0a1f1dbdfb53fc1 = I4be898887dff6e2cebe53f135ece131b + ~Ib1461f456ebc14f449eee77e386a4c69 + 1;
            Icdd0962fd06355a7dcbb491543eb9cb6 = I2bcab411f9bec1541259751bcb9e0823(I735d6229ef1a4ecda0a1f1dbdfb53fc1);
            I78f727f8d85b5d7f0ffa57f02538f939    = Icdd0962fd06355a7dcbb491543eb9cb6;

            I62affd47512c5e8f0979244115624d97 = I4be898887dff6e2cebe53f135ece131b + ~I409129c0bf5d361e9916b6dc98e69a7d + 1;
            I003f9dc1b83f386f070b0a2e8c7ce4f4 = I2bcab411f9bec1541259751bcb9e0823(I62affd47512c5e8f0979244115624d97);
            I01ec629f60c17c2251f977205234cd44    = I003f9dc1b83f386f070b0a2e8c7ce4f4;

            I14fe27afb3df5531b18dc9604e8dbe65 = I004db04f61fb57aba81e15cc015442b3 + ~I5d80b7c7d102d2c2bfa73a68c73376be + 1;
            I66e8ad34c764833f038cff700a237fcb = I2bcab411f9bec1541259751bcb9e0823(I14fe27afb3df5531b18dc9604e8dbe65);
            I23f774adb64807c0edaa9941c75651b6    = I66e8ad34c764833f038cff700a237fcb;

            Ib1b1626c84dad8ad13c058f921ffd57d = I004db04f61fb57aba81e15cc015442b3 + ~Ib2c327648cce481482eaf0467e9227d4 + 1;
            I614bddda696787a552e28cfaa81a3aa3 = I2bcab411f9bec1541259751bcb9e0823(Ib1b1626c84dad8ad13c058f921ffd57d);
            I2361ef4fd70e4c05b25289d0845564c4    = I614bddda696787a552e28cfaa81a3aa3;

            Idf4a4bdddb88c21c5afe10a02373a6eb = I004db04f61fb57aba81e15cc015442b3 + ~Iaf1d3be13e6441a7a9ab3f286a7dc21b + 1;
            I38c22e6b7c066be10ec1f8929dbf88f9 = I2bcab411f9bec1541259751bcb9e0823(Idf4a4bdddb88c21c5afe10a02373a6eb);
            Ic3067b434ca17be7bad595e1f9b822c5    = I38c22e6b7c066be10ec1f8929dbf88f9;

            Iadefc2a3d07ed4b2c3c46b2ab5dec252 = I004db04f61fb57aba81e15cc015442b3 + ~Ie4f4faa470f572da2081b63b6df6e392 + 1;
            I245816ec4a0392af2cfa4b44a4e93610 = I2bcab411f9bec1541259751bcb9e0823(Iadefc2a3d07ed4b2c3c46b2ab5dec252);
            I3546ddbae9c9db4517802db56cee35f0    = I245816ec4a0392af2cfa4b44a4e93610;

            I19315957077b037ffc6415dbb06ef789 = I8f7e3dfb2f728d4cd1e79b82b62b0406 + ~I8636f5c91b567780d3324e4b8a320fc2 + 1;
            I83253182662d56779685c9742f55789f = I2bcab411f9bec1541259751bcb9e0823(I19315957077b037ffc6415dbb06ef789);
            I35e91092ed503831ed818f36a1ce1537    = I83253182662d56779685c9742f55789f;

            I1f9be09334407fc86c83a7c127e17bbe = I8f7e3dfb2f728d4cd1e79b82b62b0406 + ~Idcc745602c4b7b34df9c3d68f9a9d76d + 1;
            I963a4391dba3d12756b89dda1e962c3f = I2bcab411f9bec1541259751bcb9e0823(I1f9be09334407fc86c83a7c127e17bbe);
            I973f185cf29e13193abf0108d4faa9d1    = I963a4391dba3d12756b89dda1e962c3f;

            I28e17a5af7a7286a2643100d6d058dc0 = I8f7e3dfb2f728d4cd1e79b82b62b0406 + ~Id5c9a9b9c34c8f9d56df0aa8d780c9d3 + 1;
            Ie959690f46f82cbb15ae0cee69f3135f = I2bcab411f9bec1541259751bcb9e0823(I28e17a5af7a7286a2643100d6d058dc0);
            Iee58b0442a6cccf0990ebb551b47fa92    = Ie959690f46f82cbb15ae0cee69f3135f;

            Icb2297c397bfe56be251ffb6b249a020 = I8f7e3dfb2f728d4cd1e79b82b62b0406 + ~I5011dfbbb0eccfebcff255e4a2c5e64c + 1;
            Ic475c578935fa69db2b1c834539750af = I2bcab411f9bec1541259751bcb9e0823(Icb2297c397bfe56be251ffb6b249a020);
            I2cb3207a5c1b25386ac7eb532955f260    = Ic475c578935fa69db2b1c834539750af;

            I64a48984527d660002f1f82c376c7a84 = I991054370345e61638ddaf81785505bd + ~I2cf5304a672431888916e08b3c15f0c7 + 1;
            I4f9bc0f2aeafb89fbaa0d0af7dbda06a = I2bcab411f9bec1541259751bcb9e0823(I64a48984527d660002f1f82c376c7a84);
            Icd4f07bc30c66f7f5b431ed97e7ac7b6    = I4f9bc0f2aeafb89fbaa0d0af7dbda06a;

            I238b5fc70ce9f05b6322a2691b3a0207 = I991054370345e61638ddaf81785505bd + ~I989091b3586964ab598f166a89279d16 + 1;
            I393fa73117dcbf1fb1b74ea1fc7e6c99 = I2bcab411f9bec1541259751bcb9e0823(I238b5fc70ce9f05b6322a2691b3a0207);
            Ifec6f3a1e10144acb320d5d502ed1ea3    = I393fa73117dcbf1fb1b74ea1fc7e6c99;

            I00c16e7ad3821981032a42d5baa767b3 = I991054370345e61638ddaf81785505bd + ~I5f7b6e6a30348ae86057f7e56f625846 + 1;
            I95836c571386b3b6de07c9195932fe22 = I2bcab411f9bec1541259751bcb9e0823(I00c16e7ad3821981032a42d5baa767b3);
            Ic87bff64a597e6d02583041b552328ee    = I95836c571386b3b6de07c9195932fe22;

            I42fd5b094da200b33036e6cb8c7d0286 = I991054370345e61638ddaf81785505bd + ~Ie32ca6b91d1c55883be8f63acca78764 + 1;
            I6dd6f9abc962974c292d22f17a21a936 = I2bcab411f9bec1541259751bcb9e0823(I42fd5b094da200b33036e6cb8c7d0286);
            I489f21ef8243ef8caa1c29f034c3e2ac    = I6dd6f9abc962974c292d22f17a21a936;

            I98b7e26a0e9ec9ad750ff87cc0641a73 = Ifa1f503965270d10e7a5c9a15576069b + ~I9164fa2a9a33da6612ea692cf3fa7d2f + 1;
            I9f9e6bc8d2cc6e41813d42ffcd5cff01 = I2bcab411f9bec1541259751bcb9e0823(I98b7e26a0e9ec9ad750ff87cc0641a73);
            I773901563077961acada85962209d68a    = I9f9e6bc8d2cc6e41813d42ffcd5cff01;

            I3ec904916870171bf837e162d1030052 = Ifa1f503965270d10e7a5c9a15576069b + ~Ie8befb003fe83e774e8d1d01d4e2f4ad + 1;
            I2ba75ccf97b5caf5aa676a9e3c42a366 = I2bcab411f9bec1541259751bcb9e0823(I3ec904916870171bf837e162d1030052);
            Ifbd176fe3e78bc2dc2e0e77ba3ccd2d0    = I2ba75ccf97b5caf5aa676a9e3c42a366;

            Iedb11b97900b7dd769d31f8a89521975 = Ifa1f503965270d10e7a5c9a15576069b + ~I1f1f2fefd3381ee48ab0ec9c9301754b + 1;
            I006699f0e016e7022b2706751965c42c = I2bcab411f9bec1541259751bcb9e0823(Iedb11b97900b7dd769d31f8a89521975);
            I53f68a4cb81c71ee7bd6f61171b7478d    = I006699f0e016e7022b2706751965c42c;

            Id0dceec6497c9f13ada07138986d4145 = Ifa1f503965270d10e7a5c9a15576069b + ~I6c7965d39dc839a9df56e628c77a5457 + 1;
            I66d5992f4f39337782cfbbb9fec3b2c8 = I2bcab411f9bec1541259751bcb9e0823(Id0dceec6497c9f13ada07138986d4145);
            I7568ec59f1359bedce86dbc6af50df71    = I66d5992f4f39337782cfbbb9fec3b2c8;

            Ibfe7d9bac29b8838f20cdcfe8ef7da0c = I24f773842a4742fb58d09cae45717b2f + ~I288ff69a7395e74f7de8da5a6a7f9062 + 1;
            Ie5f503c91ddf6eff2b9645e6e3c22b2e = I2bcab411f9bec1541259751bcb9e0823(Ibfe7d9bac29b8838f20cdcfe8ef7da0c);
            Id2bf82d6bf0a201f80a58357038a0992    = Ie5f503c91ddf6eff2b9645e6e3c22b2e;

            I4d6c95605595942a34573d6ed55eb326 = I24f773842a4742fb58d09cae45717b2f + ~I98a2aa729628adde0b6047869bd12743 + 1;
            Ieb7e6a2425e93a2b96a94f0e2c4442c3 = I2bcab411f9bec1541259751bcb9e0823(I4d6c95605595942a34573d6ed55eb326);
            I22442354ca2b77306f25839ce6124699    = Ieb7e6a2425e93a2b96a94f0e2c4442c3;

            Id6d8f32958dfa1a98958a84e7f1aed02 = I24f773842a4742fb58d09cae45717b2f + ~I1140fa91b5e22ba0c094c03295781e5a + 1;
            I4a0483f2d2585cd44fe35191d7cd88b1 = I2bcab411f9bec1541259751bcb9e0823(Id6d8f32958dfa1a98958a84e7f1aed02);
            I71a5c2876a07d8edd001ef2d108e59c1    = I4a0483f2d2585cd44fe35191d7cd88b1;

            I971cdf9ddd1bfff5664eec35f22da335 = I24f773842a4742fb58d09cae45717b2f + ~Ieac9cea5f36bd82f87105b530e8fb614 + 1;
            I00e8b3cde14889fcb0b40dc5582a58f9 = I2bcab411f9bec1541259751bcb9e0823(I971cdf9ddd1bfff5664eec35f22da335);
            Iaf333aa6b135927cf1ad1f76298ccd63    = I00e8b3cde14889fcb0b40dc5582a58f9;

            Idd8bc1412a0dc5f489ef253a6164ceea = I5bac7e0d778a547a0ae764fe259b6f7a + ~I5a4f0749acdc34fd0786e4b3d062f88b + 1;
            Ib53dbb62231f729a278d2afa3acffdbf = I2bcab411f9bec1541259751bcb9e0823(Idd8bc1412a0dc5f489ef253a6164ceea);
            Ia71cfd8cf9bea4e600ea204e41271c7d    = Ib53dbb62231f729a278d2afa3acffdbf;

            Idbeec36de0128e5924e214877c82bf11 = I5bac7e0d778a547a0ae764fe259b6f7a + ~I283107989a436e2c720123b8d9e335c2 + 1;
            I5503d6011d58dfa4e1ec524eb1875c7d = I2bcab411f9bec1541259751bcb9e0823(Idbeec36de0128e5924e214877c82bf11);
            I164b032929ac2b8cf1a6672859639a30    = I5503d6011d58dfa4e1ec524eb1875c7d;

            I50a9cd240979bc56421bf85011ae99ed = I5bac7e0d778a547a0ae764fe259b6f7a + ~Ic488e78b5c73251b673301e84c4b5b0b + 1;
            Id86fbda00d923c29c99b4a9fe52d513a = I2bcab411f9bec1541259751bcb9e0823(I50a9cd240979bc56421bf85011ae99ed);
            I2ef0447f5c64fd5c65e23c16069a62ef    = Id86fbda00d923c29c99b4a9fe52d513a;

            I6437095f6bad2d4fb2fbe0361f60bba1 = I5bac7e0d778a547a0ae764fe259b6f7a + ~I79657595561eac53237215fb4110f09d + 1;
            I3ba6e9f7d7fa98ad776299f8cd8a8363 = I2bcab411f9bec1541259751bcb9e0823(I6437095f6bad2d4fb2fbe0361f60bba1);
            Ide7008ee7f1fba156dc6145b3505e553    = I3ba6e9f7d7fa98ad776299f8cd8a8363;

            Ie9b6eb3bbac26635aa00c38110958d46 = I255577ebee6768871df0224fc1db2db3 + ~I079932780612fbce79cbe9b58bb6c2b5 + 1;
            I67b512efbaf9c063a4ac75cb97a8abdb = I2bcab411f9bec1541259751bcb9e0823(Ie9b6eb3bbac26635aa00c38110958d46);
            I129a7ced6bc6f48f20fa552e2519925c    = I67b512efbaf9c063a4ac75cb97a8abdb;

            I9f34e81e3ffb85539a6273babc2a732e = I255577ebee6768871df0224fc1db2db3 + ~I61f5ebea2bbe443b644c95ee559c2234 + 1;
            If5f5eecf512463544c8b2419c0a58779 = I2bcab411f9bec1541259751bcb9e0823(I9f34e81e3ffb85539a6273babc2a732e);
            I67123cf825352e52cf0158060ad69a13    = If5f5eecf512463544c8b2419c0a58779;

            Id0a1ab8472d704001e0eba0317b117d6 = I255577ebee6768871df0224fc1db2db3 + ~I9b46463a6c54c3668e76190d942b7b38 + 1;
            I81cdc8b54bc7f98798713985e8f4553e = I2bcab411f9bec1541259751bcb9e0823(Id0a1ab8472d704001e0eba0317b117d6);
            I09923d784a9f9625a37221f639537941    = I81cdc8b54bc7f98798713985e8f4553e;

            I9e632217cd0561d8faa28e4b8850d995 = Ia7fb4af3d3529a32f902a52cf5598474 + ~Ia92defa0ca87c7c30fbe901da40a575e + 1;
            I35bb2eb0cb589f694001ba1509cbf7f8 = I2bcab411f9bec1541259751bcb9e0823(I9e632217cd0561d8faa28e4b8850d995);
            I5947be93fdb18bf0ad341fb826c9e6d7    = I35bb2eb0cb589f694001ba1509cbf7f8;

            Iedeb5b7b2fa8acf1ea083102678710ea = Ia7fb4af3d3529a32f902a52cf5598474 + ~I21255a0ad20a9668c958faf68d53b2bc + 1;
            I3bf8f19c98c78f8e1c315e75a533bb1c = I2bcab411f9bec1541259751bcb9e0823(Iedeb5b7b2fa8acf1ea083102678710ea);
            I08621ee033cd49702ad08af4d31eb999    = I3bf8f19c98c78f8e1c315e75a533bb1c;

            I972431d1f5af0bdf4828e4f85591e358 = Ia7fb4af3d3529a32f902a52cf5598474 + ~I3ff883ad434cd5153b67186b6b21418d + 1;
            I71cbdcd6e3a873851e9084bc9dcd99bd = I2bcab411f9bec1541259751bcb9e0823(I972431d1f5af0bdf4828e4f85591e358);
            Id5eca60b22d3835119571fe4b1a03479    = I71cbdcd6e3a873851e9084bc9dcd99bd;

            I1f41024b715d8312944ccbf70e95bb40 = I2c98806141f064c9e92935b23a84ede1 + ~I914bef0326cf82d350344317eb1359be + 1;
            Iebad2e3d84bae3d4807badae823aec52 = I2bcab411f9bec1541259751bcb9e0823(I1f41024b715d8312944ccbf70e95bb40);
            I7267ba2b9cb511a48a3a7044e854f7da    = Iebad2e3d84bae3d4807badae823aec52;

            Ia6bb5ca05f5d0af452c994dd50004e1d = I2c98806141f064c9e92935b23a84ede1 + ~I6f69796a6fe6da57066319ec8210c1a3 + 1;
            I054f07cdf6a44100034c7e2fb438055f = I2bcab411f9bec1541259751bcb9e0823(Ia6bb5ca05f5d0af452c994dd50004e1d);
            I5893fa21ec8bbdcea9677cc12fc4057a    = I054f07cdf6a44100034c7e2fb438055f;

            I9a1d1d1c862808f9a769cbdb3bc634e1 = I2c98806141f064c9e92935b23a84ede1 + ~I92abaae6fb89206885616877cca1e25a + 1;
            If3b82307d1ad78e262f76ba9b711e1a6 = I2bcab411f9bec1541259751bcb9e0823(I9a1d1d1c862808f9a769cbdb3bc634e1);
            I564896fe01ec799a0fbe790473753559    = If3b82307d1ad78e262f76ba9b711e1a6;

            I9734eb86f4e73ba217739baf5cb1b13c = I5680847bc8d224fa4ed93b2fc0d841e1 + ~Ie43a7f8082f91c2955076a6373028b55 + 1;
            I0f40c8301521c136b3ede2cc9e8352a3 = I2bcab411f9bec1541259751bcb9e0823(I9734eb86f4e73ba217739baf5cb1b13c);
            If279ab7c515c4039c8272b913c2fa107    = I0f40c8301521c136b3ede2cc9e8352a3;

            Ifc0fe00f86569956df72d8a960337e8c = I5680847bc8d224fa4ed93b2fc0d841e1 + ~I8786eb767f02164cdc32f14f41b5d0e1 + 1;
            I3615a34cbf1646a7cd0f1da43d62faa5 = I2bcab411f9bec1541259751bcb9e0823(Ifc0fe00f86569956df72d8a960337e8c);
            Ib61705ff5820f531eb17c40ed05f6ec3    = I3615a34cbf1646a7cd0f1da43d62faa5;

            I223341a807a1d555f759632f67815159 = I5680847bc8d224fa4ed93b2fc0d841e1 + ~I33668b0ef7defef974b7a4c0f87689c0 + 1;
            I0bbd697ad8d3877570ab9e200e66164a = I2bcab411f9bec1541259751bcb9e0823(I223341a807a1d555f759632f67815159);
            I50149e5de41ca2998c4e8cc4b19e166b    = I0bbd697ad8d3877570ab9e200e66164a;

            I6c1f5cdf5f2917118941f4af14d67fef = I365254279ebb10dd7ba0b3482d5e34cd + ~Ibfb57f2b507c27759a3556759f23977b + 1;
            I298f7389a7fd8e927b7e3354f0d32344 = I2bcab411f9bec1541259751bcb9e0823(I6c1f5cdf5f2917118941f4af14d67fef);
            Id40cac3272643f3f91b73c6aa1740f3b    = I298f7389a7fd8e927b7e3354f0d32344;

            Ie84e88fd1aa2a0b90aa1715fcd27a329 = I365254279ebb10dd7ba0b3482d5e34cd + ~I064499f0315fbeec7b6cb50583388a07 + 1;
            I9960d39fce3c5b9945965dedac46dfed = I2bcab411f9bec1541259751bcb9e0823(Ie84e88fd1aa2a0b90aa1715fcd27a329);
            Ic63eee2d700493c41ee2d186ff7111b9    = I9960d39fce3c5b9945965dedac46dfed;

            I558f70d7039a8bb58d8ea3f72e43dac0 = I365254279ebb10dd7ba0b3482d5e34cd + ~Ica0a119af1728ae253c16cc3eb93f802 + 1;
            I02f48e93599dc91bb24a144a0ef1a933 = I2bcab411f9bec1541259751bcb9e0823(I558f70d7039a8bb58d8ea3f72e43dac0);
            I51de42598e0df4a76cf7b02c61ae9550    = I02f48e93599dc91bb24a144a0ef1a933;

            I9924269ed3de12f1f2a28893c7f95292 = I365254279ebb10dd7ba0b3482d5e34cd + ~Ib7875bf9d30d071e62a474c50d88ba06 + 1;
            I7e31af1959a0374af6c2767e4837c566 = I2bcab411f9bec1541259751bcb9e0823(I9924269ed3de12f1f2a28893c7f95292);
            Ia89a1a58f6327ee3c105cae860942171    = I7e31af1959a0374af6c2767e4837c566;

            If1153befd1396be2798cc14535ddeb8a = I365254279ebb10dd7ba0b3482d5e34cd + ~I338daeacf82ad288b14c6b5bd4099870 + 1;
            I8d18e2ecaf2bda4a0ba47d9782e9917a = I2bcab411f9bec1541259751bcb9e0823(If1153befd1396be2798cc14535ddeb8a);
            Ib149a5872e31cd5df77b66298b4aad12    = I8d18e2ecaf2bda4a0ba47d9782e9917a;

            I9bc447b20687fb3e7eff45792bd4dc3a = I57bf4ad773cc058ae1bb7b1911dc3174 + ~I7b12345fe53174cadef6811fb8869b42 + 1;
            Id0a13655f967dfd3000b8dcf4a57f555 = I2bcab411f9bec1541259751bcb9e0823(I9bc447b20687fb3e7eff45792bd4dc3a);
            Iaa16c14572ad0442eb3c58a97bef5ada    = Id0a13655f967dfd3000b8dcf4a57f555;

            If590520f01e452db9867a8d6d5dab29b = I57bf4ad773cc058ae1bb7b1911dc3174 + ~I6521c9167261db6eb37f50b66159ddb7 + 1;
            Ibf384c0b998b5a5f7808c54292c6b844 = I2bcab411f9bec1541259751bcb9e0823(If590520f01e452db9867a8d6d5dab29b);
            I88d5d48e05b1c9a6d8060f58917e3834    = Ibf384c0b998b5a5f7808c54292c6b844;

            Id93ee7d283016ab9b0aaa21237237c54 = I57bf4ad773cc058ae1bb7b1911dc3174 + ~I44e5ce0cdf812c5b73e6e638da36e414 + 1;
            I58b8202ae510e96b4f6ae334f3b282c6 = I2bcab411f9bec1541259751bcb9e0823(Id93ee7d283016ab9b0aaa21237237c54);
            I4269e18c2df4d39c683ffb7d01a08322    = I58b8202ae510e96b4f6ae334f3b282c6;

            Ic1cf03baabaed466fe532e4db3a9ea78 = I57bf4ad773cc058ae1bb7b1911dc3174 + ~I6fdccefd034e8b4b86cfa997502512ae + 1;
            Icbc75d6e4d0bcc42cdf813529b017e0e = I2bcab411f9bec1541259751bcb9e0823(Ic1cf03baabaed466fe532e4db3a9ea78);
            Ia29017fa9327fdaa7c10b2797f8aa6ec    = Icbc75d6e4d0bcc42cdf813529b017e0e;

            If3031f9aa8f6eba90eac12db7839fefd = I57bf4ad773cc058ae1bb7b1911dc3174 + ~Ibe085a39ecb07a8dca62002afa38df93 + 1;
            I6fa1835a8e7f8ea435c4515b1c059cc9 = I2bcab411f9bec1541259751bcb9e0823(If3031f9aa8f6eba90eac12db7839fefd);
            Ia142ac799256541fe33f898a6a31dd71    = I6fa1835a8e7f8ea435c4515b1c059cc9;

            I0dc2708970ca2b6c092273b6626bacd6 = I57072dfb29c4a3d2e2b40e46e62f0d95 + ~I9785922874bba479ce4a9bf1759e2933 + 1;
            Id3984a3dd1009c9c76347b9843f27b25 = I2bcab411f9bec1541259751bcb9e0823(I0dc2708970ca2b6c092273b6626bacd6);
            I4c039794243933a9bb7ad6db7eda6a87    = Id3984a3dd1009c9c76347b9843f27b25;

            Ia58944aebf0b4f0a7d76a1444fced9de = I57072dfb29c4a3d2e2b40e46e62f0d95 + ~I0e3286fca6cd040758950259ab663df7 + 1;
            Id5fd757abdc0b2e1b1d4c5dab96ee08a = I2bcab411f9bec1541259751bcb9e0823(Ia58944aebf0b4f0a7d76a1444fced9de);
            I0debb3ed4f9540c162cd525588e0ae3f    = Id5fd757abdc0b2e1b1d4c5dab96ee08a;

            Iedd8e69679d10e05f2889f1d71cf0e7b = I57072dfb29c4a3d2e2b40e46e62f0d95 + ~I9ae284c0089ae462a1bb9d168bde2fd0 + 1;
            I98ab1b82b2991b4cb3bec530711bdc43 = I2bcab411f9bec1541259751bcb9e0823(Iedd8e69679d10e05f2889f1d71cf0e7b);
            I681eed68ee814fb18fd794207d9266e1    = I98ab1b82b2991b4cb3bec530711bdc43;

            I90f0d471914a2333b9dc14d6d01cf927 = I57072dfb29c4a3d2e2b40e46e62f0d95 + ~I202aa0814e7e28a6bd21db116b652b4d + 1;
            I610d0ed6f55a4906aac1be5823358392 = I2bcab411f9bec1541259751bcb9e0823(I90f0d471914a2333b9dc14d6d01cf927);
            Ic260784b8910f5a0483afee9b68efb31    = I610d0ed6f55a4906aac1be5823358392;

            Idceeb22013af64b6bb9f0d773e9ffe9a = I57072dfb29c4a3d2e2b40e46e62f0d95 + ~I1f88dddf05f255942e2749891a7733da + 1;
            I2ed0ad73f73f9f4e1b7ec38af320ee4d = I2bcab411f9bec1541259751bcb9e0823(Idceeb22013af64b6bb9f0d773e9ffe9a);
            I22cd2d30a7684002cacca4deae4c95a0    = I2ed0ad73f73f9f4e1b7ec38af320ee4d;

            If43574342e60a625fb6bee5a495e88f3 = Id8cafb6f76321bdaba9711133be7be99 + ~Ie7e196fbb66ba6bee51ef0064ca519c2 + 1;
            I3dfc4dd447cd1f4e40506f516c106861 = I2bcab411f9bec1541259751bcb9e0823(If43574342e60a625fb6bee5a495e88f3);
            I136b4136d582f9fad21f90297cfafea3    = I3dfc4dd447cd1f4e40506f516c106861;

            Id285f055275014d9f23d35f91879afa1 = Id8cafb6f76321bdaba9711133be7be99 + ~Id7619819e1297844d92c8bf3a1d61926 + 1;
            Idfeea354b3f9ca8c671851fd90f4e1bc = I2bcab411f9bec1541259751bcb9e0823(Id285f055275014d9f23d35f91879afa1);
            Id8d6be9677d3b0ceca26b3b671757c2c    = Idfeea354b3f9ca8c671851fd90f4e1bc;

            I8c803ab08db372802117de4fa4e2a187 = Id8cafb6f76321bdaba9711133be7be99 + ~If8a259e0c4f1839e852abec6e1b904ee + 1;
            I415d8306edb869fc838eb518aad75168 = I2bcab411f9bec1541259751bcb9e0823(I8c803ab08db372802117de4fa4e2a187);
            I6a93f928c104ea211dcc8a461506327d    = I415d8306edb869fc838eb518aad75168;

            I13ba48a6b360f3cff5f37ce60cb735c6 = Id8cafb6f76321bdaba9711133be7be99 + ~Ib2f34922b0d5346500de093275bebc94 + 1;
            I1dc6b2aef1bb326c3d5c19f97a2e1d4f = I2bcab411f9bec1541259751bcb9e0823(I13ba48a6b360f3cff5f37ce60cb735c6);
            I240da147648bec33195a5f5c273fc6f4    = I1dc6b2aef1bb326c3d5c19f97a2e1d4f;

            I4547cd1dad45dfd01e335e8cf20eadd6 = Id8cafb6f76321bdaba9711133be7be99 + ~If1d0be4e9b995ec98c346e8392b9518a + 1;
            Ie2f47a06ca4b6d5823cbbe099f5de0f0 = I2bcab411f9bec1541259751bcb9e0823(I4547cd1dad45dfd01e335e8cf20eadd6);
            I55494d0e8454e3cbb4158559e0d29984    = Ie2f47a06ca4b6d5823cbbe099f5de0f0;

            I0a305655b815b0cc159ac1c5f4ce30f8 = I6344e71ca2b0fd39d36caedd889c3085 + ~Ibb157b97546cb19fa7c1c0a7c79b1d38 + 1;
            I55b7a58384e50ade254c3c8934c290f6 = I2bcab411f9bec1541259751bcb9e0823(I0a305655b815b0cc159ac1c5f4ce30f8);
            Ied3cc579b3cf126081acf8e1117007cf    = I55b7a58384e50ade254c3c8934c290f6;

            I3633737da6b74284b0ea9a06c3f5875f = I6344e71ca2b0fd39d36caedd889c3085 + ~I3fdec80112b3fc543b217d1c253406da + 1;
            I53bf5dca5911aec50866be5a720d4aa2 = I2bcab411f9bec1541259751bcb9e0823(I3633737da6b74284b0ea9a06c3f5875f);
            I76140bdc374dd6031097575fd231b468    = I53bf5dca5911aec50866be5a720d4aa2;

            Ia949c1b338d1cba07cf6bb6572c3e322 = I6344e71ca2b0fd39d36caedd889c3085 + ~I56a4443759b3d786bc9a34a0dc32abf0 + 1;
            Ie57f78d4c002e69e0e92b25bad752d3f = I2bcab411f9bec1541259751bcb9e0823(Ia949c1b338d1cba07cf6bb6572c3e322);
            I650345d21e5c2e7a9bf1810630161089    = Ie57f78d4c002e69e0e92b25bad752d3f;

            I9a0185f8400159415bc0ad6c38284041 = I0c99a68e0bed90afce18807acf7d55bb + ~I8fb1602dcdcd2912ea8aec42e2b7848f + 1;
            I2ac511a908c9973254672fd38cabccd3 = I2bcab411f9bec1541259751bcb9e0823(I9a0185f8400159415bc0ad6c38284041);
            Ie852635f073dc918e7b1075ffad46f24    = I2ac511a908c9973254672fd38cabccd3;

            I3eeffe43e7deed7ee77a7f5a3bce3cd2 = I0c99a68e0bed90afce18807acf7d55bb + ~I5aa85d9503b0e4ff46bbd63e873053ca + 1;
            I8f06d78dd2e6be736f4e4f41fadf130d = I2bcab411f9bec1541259751bcb9e0823(I3eeffe43e7deed7ee77a7f5a3bce3cd2);
            I9ec80c14eb5f0f305e1a9e6107a6001e    = I8f06d78dd2e6be736f4e4f41fadf130d;

            I85af0c31ca7002ae569d9f5ce39943f7 = I0c99a68e0bed90afce18807acf7d55bb + ~Ic826d371f2cfc503f5d9e43dc17481e1 + 1;
            I65450e396e33720967b7a6271e3a70e1 = I2bcab411f9bec1541259751bcb9e0823(I85af0c31ca7002ae569d9f5ce39943f7);
            I80ba56447ab19b33610c23105b0b1637    = I65450e396e33720967b7a6271e3a70e1;

            I3dfb8d2fad83fbd807fbfc6330c5b857 = I1c95650979c86310ae2a949961c9db11 + ~I7de222bc26e38b8b6543819701740302 + 1;
            I876c6361d2164d03cad2ffc8bf920ac0 = I2bcab411f9bec1541259751bcb9e0823(I3dfb8d2fad83fbd807fbfc6330c5b857);
            Ib9132d9fa7180c3fcbacb7c570d6b0f2    = I876c6361d2164d03cad2ffc8bf920ac0;

            Ic12be21bcba5fa49437cc44dd8a7f064 = I1c95650979c86310ae2a949961c9db11 + ~Ia7673d73f0535906a99d6cb467892104 + 1;
            Id3b8e1157a3e9eea4d210f466740f673 = I2bcab411f9bec1541259751bcb9e0823(Ic12be21bcba5fa49437cc44dd8a7f064);
            I01621f113f636a9caf9b5ca0bb20ef77    = Id3b8e1157a3e9eea4d210f466740f673;

            I713a384d022d3012e3d0019f5c4ac077 = I1c95650979c86310ae2a949961c9db11 + ~I5502f383dff392ef1be4cbbf9dbc3c2f + 1;
            I6973de59fb6014d7c4bf5b982cddc4d8 = I2bcab411f9bec1541259751bcb9e0823(I713a384d022d3012e3d0019f5c4ac077);
            I3eeddb549c6e1f07469c0e0dca68be92    = I6973de59fb6014d7c4bf5b982cddc4d8;

            I80550019479d0323d0dd7e7d0f767d83 = I04eaefa5d133e53494fc270b07be7043 + ~Iea765ae5e9c65b3186445b15c56f69e5 + 1;
            I26cb99c4cc37be5f52dfeeca60d5d102 = I2bcab411f9bec1541259751bcb9e0823(I80550019479d0323d0dd7e7d0f767d83);
            Ibe664dd203ed4162abcd36eb8d57bfa6    = I26cb99c4cc37be5f52dfeeca60d5d102;

            Ib8a866f080dd997e0b6c93b6c844d1bc = I04eaefa5d133e53494fc270b07be7043 + ~I103ec7cf279f527fc6e3648a19a12a8a + 1;
            Ie9835b1d512d9c9c4f2801956fbf13cb = I2bcab411f9bec1541259751bcb9e0823(Ib8a866f080dd997e0b6c93b6c844d1bc);
            Ia66176893fe306ecfb415d948c50486d    = Ie9835b1d512d9c9c4f2801956fbf13cb;

            Id542de206d736ee3769ea0bd037cb627 = I04eaefa5d133e53494fc270b07be7043 + ~I96e6f1dc0cd451da6ac9170d5f83976d + 1;
            I89057e4e979b903ae1f10f9dd2f196fe = I2bcab411f9bec1541259751bcb9e0823(Id542de206d736ee3769ea0bd037cb627);
            I8bd4210dcbfc1956381b460fd9ef789b    = I89057e4e979b903ae1f10f9dd2f196fe;

            I77e6cdb09c92492c3303d0213de9c291 = I4a64fa2412eb8058c2dfd9351d7b297d + ~Icf266f710358631b7119ef526acb301c + 1;
            If1299e6b34cd1f2239d64ade23f33f01 = I2bcab411f9bec1541259751bcb9e0823(I77e6cdb09c92492c3303d0213de9c291);
            I1ba6328ea9cb7cebcce47d5407d0eae7    = If1299e6b34cd1f2239d64ade23f33f01;

            I788c33a9f94b26f4ce0f515891d06f90 = I4a64fa2412eb8058c2dfd9351d7b297d + ~Ib20dec1346f227042c749ec1abfa4d39 + 1;
            I3f106ef1876021bb3cc5866d2b5698f4 = I2bcab411f9bec1541259751bcb9e0823(I788c33a9f94b26f4ce0f515891d06f90);
            I9e79c17bd782bb7981b4a3623baf96a1    = I3f106ef1876021bb3cc5866d2b5698f4;

            Iaf7074c2b570a296fe2ea8a5a7097ca0 = I4a64fa2412eb8058c2dfd9351d7b297d + ~Id6fa8ec5d1062fc3e09bdac65ff79f45 + 1;
            If6cb9fec3dc380f1c4894bccfa35b33c = I2bcab411f9bec1541259751bcb9e0823(Iaf7074c2b570a296fe2ea8a5a7097ca0);
            I7c6f64d73ff9c6e7f2ed69713e056a2b    = If6cb9fec3dc380f1c4894bccfa35b33c;

            I8964c6d3f8e02866a6ad86553ab05d99 = I4a64fa2412eb8058c2dfd9351d7b297d + ~I10cd840a369d3e25556a41beede2be27 + 1;
            I313980f8406e9f26d5eaa53270a23b9e = I2bcab411f9bec1541259751bcb9e0823(I8964c6d3f8e02866a6ad86553ab05d99);
            I00b962a9bf04b62244591051d2dfdbbd    = I313980f8406e9f26d5eaa53270a23b9e;

            I2aa25edaca90c9dae8ed63b48d333c17 = Ie8bb2fcb752c6a33254963d1ebb4130d + ~I0f3c4fb63ef1e88168b4d28175a0b68c + 1;
            I792b5aea212da69a9c18f5723e820432 = I2bcab411f9bec1541259751bcb9e0823(I2aa25edaca90c9dae8ed63b48d333c17);
            I3a660b57588325989319701026f658e6    = I792b5aea212da69a9c18f5723e820432;

            I51a440917c7ae23339bec6f8a745c103 = Ie8bb2fcb752c6a33254963d1ebb4130d + ~Iac6fcccf3a0cfe04edc0d998b60c2681 + 1;
            I98f245ec9b667dc065c9494c00ecdf88 = I2bcab411f9bec1541259751bcb9e0823(I51a440917c7ae23339bec6f8a745c103);
            Ibae27cccf3f64e8653c1e244e940e421    = I98f245ec9b667dc065c9494c00ecdf88;

            I56ce875e4619d4d8d6ca2fa0ddee91b1 = Ie8bb2fcb752c6a33254963d1ebb4130d + ~I1fbcaf2f6be01b129ebc24dee8a65396 + 1;
            I15254b39b6e136520a9497d8684f9d94 = I2bcab411f9bec1541259751bcb9e0823(I56ce875e4619d4d8d6ca2fa0ddee91b1);
            I27b89a5001312b2aa48fe385d8a52063    = I15254b39b6e136520a9497d8684f9d94;

            I80607da8f92f5a5d2e4798a62a7b1c5c = Ie8bb2fcb752c6a33254963d1ebb4130d + ~Id85c2285fcc45211f0fa6963b74a663a + 1;
            I6c8312a9d655f143a0b65d91907ce533 = I2bcab411f9bec1541259751bcb9e0823(I80607da8f92f5a5d2e4798a62a7b1c5c);
            Ic6a7476db711a812d146331c562ca7c9    = I6c8312a9d655f143a0b65d91907ce533;

            Ic4dcaa520e26bac40b3876f02074f856 = Iac05b7e3ae18f948b72c356ccfb8000f + ~I2ba94ef71f97b9ba731b306d4a5fd02c + 1;
            Ie6df2f89b05947f6be3b64e3b4f23df3 = I2bcab411f9bec1541259751bcb9e0823(Ic4dcaa520e26bac40b3876f02074f856);
            I01ca07fe91b5f1edf87300b3583e77c5    = Ie6df2f89b05947f6be3b64e3b4f23df3;

            I3b2714d34081a3b6cccc47fa1638e72e = Iac05b7e3ae18f948b72c356ccfb8000f + ~Ifbaae8b3da03911a4c96d4efdb9283c5 + 1;
            Ia71232b0b468b729fa1262957cbe9faa = I2bcab411f9bec1541259751bcb9e0823(I3b2714d34081a3b6cccc47fa1638e72e);
            I6da707fd74249175d1f68dccb66390c0    = Ia71232b0b468b729fa1262957cbe9faa;

            I2db1d1ee8f546c00e512875ce2e13cee = Iac05b7e3ae18f948b72c356ccfb8000f + ~Ifba1584d599da13b98a3b76b4db10974 + 1;
            If75d8d882c6afc3df62096486b8e5b80 = I2bcab411f9bec1541259751bcb9e0823(I2db1d1ee8f546c00e512875ce2e13cee);
            I0ae62aae426b75b06d95c46baf33f08e    = If75d8d882c6afc3df62096486b8e5b80;

            If80a6bb104ff3b2020e909103c104063 = Iac05b7e3ae18f948b72c356ccfb8000f + ~Ie0bdfac78159144aa65090028931a3bf + 1;
            I7ed551b891500784c827992eb53f9ef9 = I2bcab411f9bec1541259751bcb9e0823(If80a6bb104ff3b2020e909103c104063);
            Iec512b5870f295a50921e7e0289a7d35    = I7ed551b891500784c827992eb53f9ef9;

            Iadb72cc5444816fbd132256493930bb4 = I27da3f75cca6c49e55db90306aa68e94 + ~I5529d6db17b6184c45cc4487e5a2c24a + 1;
            I5b5a24fd7116acd8ad2161513848c6a2 = I2bcab411f9bec1541259751bcb9e0823(Iadb72cc5444816fbd132256493930bb4);
            I3aac84acd9d78070472b1cbc745c80a7    = I5b5a24fd7116acd8ad2161513848c6a2;

            I3a8ec1ad07bfada3d2c6ffca88b8b678 = I27da3f75cca6c49e55db90306aa68e94 + ~I685699f60c76b00df87c9c53e9a8e448 + 1;
            Id7055f4e578533dbd25d0505f8e47f34 = I2bcab411f9bec1541259751bcb9e0823(I3a8ec1ad07bfada3d2c6ffca88b8b678);
            Ibbb900f56de318bf6e65b49791835ef4    = Id7055f4e578533dbd25d0505f8e47f34;

            I0aa042b86d9f68d22a49b4eb480a9088 = I27da3f75cca6c49e55db90306aa68e94 + ~Idb862697f62a6c678072de760e176096 + 1;
            I9c78f3a2aa3986718caf8e70d4d939d4 = I2bcab411f9bec1541259751bcb9e0823(I0aa042b86d9f68d22a49b4eb480a9088);
            I2c2ac1e722fba72c759f1d37b88a9a10    = I9c78f3a2aa3986718caf8e70d4d939d4;

            I89a387374771b68d87d7ff2dcc810829 = I27da3f75cca6c49e55db90306aa68e94 + ~I28fa30cd1f3b476fa6a354863108cbcf + 1;
            I2def789e23f8ea0edee6f58200144096 = I2bcab411f9bec1541259751bcb9e0823(I89a387374771b68d87d7ff2dcc810829);
            Ida0a18f1b79aff4ddf0e8f7e27794674    = I2def789e23f8ea0edee6f58200144096;

            I2935b3d5c3bba4dddfc7ae03fa77b229 = Idc7fed723190098341225fe01ba65ced + ~Ie3361a270ebc41698ef4651bb3548a49 + 1;
            I319c2cb3a815a6347511f0c398876a3c = I2bcab411f9bec1541259751bcb9e0823(I2935b3d5c3bba4dddfc7ae03fa77b229);
            I9f2029db42c5a968b370587c958c8929    = I319c2cb3a815a6347511f0c398876a3c;

            I4e0c0248f4aa97d263d64dfec36e3aa2 = Idc7fed723190098341225fe01ba65ced + ~Id0842da8068ee88d99af7acea50e7b77 + 1;
            I0603434655e30a66d4e00b2bc2c878c0 = I2bcab411f9bec1541259751bcb9e0823(I4e0c0248f4aa97d263d64dfec36e3aa2);
            If5755f4f61a89d91a91188c17ff5dc5a    = I0603434655e30a66d4e00b2bc2c878c0;

            Ia2871d7493b2727d2cb2fbab596b7e6a = Idc7fed723190098341225fe01ba65ced + ~I7a927f4f266cc5253ec30f5c127bb17a + 1;
            Ia6f16190b83b661f68a7a217bb356bdc = I2bcab411f9bec1541259751bcb9e0823(Ia2871d7493b2727d2cb2fbab596b7e6a);
            I4419d97c3174ee4610eb6ee9c06cb256    = Ia6f16190b83b661f68a7a217bb356bdc;

            Ie57adae8873946d6c706074b52a49786 = Ife9065805598960919ee4f14c3cc6fd4 + ~I74b55d2f94073ba8f948e4b02386867c + 1;
            I68fc61dbee0900bd66be7c7f5aaf8825 = I2bcab411f9bec1541259751bcb9e0823(Ie57adae8873946d6c706074b52a49786);
            Ia964f83676273055e20a2f63c8fffa0d    = I68fc61dbee0900bd66be7c7f5aaf8825;

            If5ac85646e4b339a19af658f01d0a17f = Ife9065805598960919ee4f14c3cc6fd4 + ~I03a8a458ee0942c35001cbfe8e589222 + 1;
            I4ddd7ecf84b4ee4a4b6290f3d362f190 = I2bcab411f9bec1541259751bcb9e0823(If5ac85646e4b339a19af658f01d0a17f);
            Iab4fbc811e87df1d1f5821ea732b6a93    = I4ddd7ecf84b4ee4a4b6290f3d362f190;

            I1c092426f34be030b3e020f40517b0e1 = Ife9065805598960919ee4f14c3cc6fd4 + ~I7571c7c306861230de71a75fca79c5dc + 1;
            I8e60b67eb6a187737de2717ebb95cf6c = I2bcab411f9bec1541259751bcb9e0823(I1c092426f34be030b3e020f40517b0e1);
            I4fbefbb10724b0844c95e85495d4a87f    = I8e60b67eb6a187737de2717ebb95cf6c;

            Ic719b72ad271bc7c077067518e6bbb98 = I717c5c2d6a2be61593492ae5f17a112f + ~I45cb51c25c426c296f97a5d23a08c063 + 1;
            I7e17264500cb48d228c20542c40169cb = I2bcab411f9bec1541259751bcb9e0823(Ic719b72ad271bc7c077067518e6bbb98);
            I717217d0b5a526f04c7f5ab0835dd5c7    = I7e17264500cb48d228c20542c40169cb;

            Ib87362230682c88d68a0ba70e25f3c20 = I717c5c2d6a2be61593492ae5f17a112f + ~Ic1af7410a9d11c5324f3ee5b2e0e9dac + 1;
            I6bddfc7b277ff042899fb2acd5625c5e = I2bcab411f9bec1541259751bcb9e0823(Ib87362230682c88d68a0ba70e25f3c20);
            I235937b643e8f2848116dc76c43f47a7    = I6bddfc7b277ff042899fb2acd5625c5e;

            Ifcf097a102f8dc1f912022fed893d222 = I717c5c2d6a2be61593492ae5f17a112f + ~Ic79811a48840357d0b6303e7b19413dc + 1;
            I6daafbc7b14e2736b2a4e29c5f6fc5ff = I2bcab411f9bec1541259751bcb9e0823(Ifcf097a102f8dc1f912022fed893d222);
            I7481f17d659cce5b4c72a68a9f6be67f    = I6daafbc7b14e2736b2a4e29c5f6fc5ff;

            I56483ca3fa550dc59bfa347780cfef7b = I4c31fa8e6eb648439cdae1de1afe0d6f + ~I0cedca0e2c589104d6f3318505910594 + 1;
            I29df797d4c3ebd64fb088660bf89e922 = I2bcab411f9bec1541259751bcb9e0823(I56483ca3fa550dc59bfa347780cfef7b);
            I5715c21c80992a61bff8aabc3f80415b    = I29df797d4c3ebd64fb088660bf89e922;

            I4aa9f61be376458185c3235442c8fda0 = I4c31fa8e6eb648439cdae1de1afe0d6f + ~Ica02d19b129c8b1d491ea4747a55113e + 1;
            I9418cc6766916bf1afc1f8a01feaad4e = I2bcab411f9bec1541259751bcb9e0823(I4aa9f61be376458185c3235442c8fda0);
            I434e3216a615eb46be5c26ef914b9cd2    = I9418cc6766916bf1afc1f8a01feaad4e;

            Id91fde1007d47258273299de80721390 = I4c31fa8e6eb648439cdae1de1afe0d6f + ~I0f29300446f020dd23cf847d3e3d3530 + 1;
            I90e1a5b43e93c02512a76c5cab15c5ad = I2bcab411f9bec1541259751bcb9e0823(Id91fde1007d47258273299de80721390);
            I918326ac0a744d234d74e2c08cf41eb4    = I90e1a5b43e93c02512a76c5cab15c5ad;

            Id58498c34aff2e1216c189b9df88822c = Iead549a9af27f1fced7d9c36e7b5c3f5 + ~I77a54091bc2c3d9006ecb3471b94d8c8 + 1;
            I26977fe4cdb2f9714fae2f12ca4a809b = I2bcab411f9bec1541259751bcb9e0823(Id58498c34aff2e1216c189b9df88822c);
            I966706d314f4c0a7ec842dd699d34926    = I26977fe4cdb2f9714fae2f12ca4a809b;

            Ib52e0c68caadcf4dd9636a84f5460e53 = Iead549a9af27f1fced7d9c36e7b5c3f5 + ~I1c0df8c2c64b688ae417a238263f33db + 1;
            I59775b68e199902c38d62e28cff01393 = I2bcab411f9bec1541259751bcb9e0823(Ib52e0c68caadcf4dd9636a84f5460e53);
            I5a7d246d88ef12e999f4bdee40e5a585    = I59775b68e199902c38d62e28cff01393;

            Ie19679053b289bb5a0aad570cc81bd14 = Iead549a9af27f1fced7d9c36e7b5c3f5 + ~I696db0b98e27dcc4657dc7feb23a881b + 1;
            I9470ef82dad13754d8d061b5fd00a667 = I2bcab411f9bec1541259751bcb9e0823(Ie19679053b289bb5a0aad570cc81bd14);
            Ic2dfaf65c4e17a8dcd55f766c314d6ef    = I9470ef82dad13754d8d061b5fd00a667;

            I8862c5ef45b723c9abf5d0ab6854a900 = Iead549a9af27f1fced7d9c36e7b5c3f5 + ~I9de41d0b279b84366640880dbd18c502 + 1;
            I62eb7a176351be84d086ce3c463214e8 = I2bcab411f9bec1541259751bcb9e0823(I8862c5ef45b723c9abf5d0ab6854a900);
            I151831ba6bd0e162275c84815e3c0f12    = I62eb7a176351be84d086ce3c463214e8;

            I30db951a07af96a8ddf59360141b9a6a = Iead549a9af27f1fced7d9c36e7b5c3f5 + ~I802bd5b13c183c37e842f7e9278f35a9 + 1;
            I106eb0d8f9ea92cda7bec4fe4aed6409 = I2bcab411f9bec1541259751bcb9e0823(I30db951a07af96a8ddf59360141b9a6a);
            I5a8f1675234ebed14d719344b530bbd7    = I106eb0d8f9ea92cda7bec4fe4aed6409;

            I4855a0a0c6426d33014ce6a4c96965ce = I10422eb79364e7d0e21e1643d9060331 + ~Ib6c0e635e659f54724737f0cffd1b0fc + 1;
            Id0c12bc1a2139e57ea40c3254f30de7b = I2bcab411f9bec1541259751bcb9e0823(I4855a0a0c6426d33014ce6a4c96965ce);
            I95dce76a8d0e729d40fb3f573cfc06ad    = Id0c12bc1a2139e57ea40c3254f30de7b;

            I362e8db1791718290bd33a79b4fc0855 = I10422eb79364e7d0e21e1643d9060331 + ~Iad0f4602ec545dc6ef12aa34add00ed3 + 1;
            Ib809a6099992799ce0235f22ce798c9a = I2bcab411f9bec1541259751bcb9e0823(I362e8db1791718290bd33a79b4fc0855);
            I6c26c7918254426c18f2e747c91438c5    = Ib809a6099992799ce0235f22ce798c9a;

            I773f0508440fb71d73fd82a372cc0a00 = I10422eb79364e7d0e21e1643d9060331 + ~Idfa432a87877e1ce103e56891745b62a + 1;
            I1a9be3897e044e9b24ac330ef3a20419 = I2bcab411f9bec1541259751bcb9e0823(I773f0508440fb71d73fd82a372cc0a00);
            I0414ead2472e42da8a271cb0bd1debf4    = I1a9be3897e044e9b24ac330ef3a20419;

            I792891cecae468d7a87e12f2da62a718 = I10422eb79364e7d0e21e1643d9060331 + ~Iba52b84e6e215842e0ca8e72c42ebce7 + 1;
            I6e87b3400b7ddab94faf11c3910fa534 = I2bcab411f9bec1541259751bcb9e0823(I792891cecae468d7a87e12f2da62a718);
            Ic6a6f5090470a76ddb7315c022ddc104    = I6e87b3400b7ddab94faf11c3910fa534;

            I33303820ad094d7a0ab53bca722fc609 = I10422eb79364e7d0e21e1643d9060331 + ~I0297905b35f06697625420b7fc2434f7 + 1;
            I51e0ff0f52ca609663781545174b763d = I2bcab411f9bec1541259751bcb9e0823(I33303820ad094d7a0ab53bca722fc609);
            I2a00ee56a5aa639f45eb3b1bdcffe81c    = I51e0ff0f52ca609663781545174b763d;

            Iff98739de575e25104c0dc30f08912a5 = I914cb87eba8baa40cd515334e59f26b2 + ~Ifba318d4faf308168c5eac8fe92395b4 + 1;
            I5c523df1fb2161ab4efd1c9b3e6b7aef = I2bcab411f9bec1541259751bcb9e0823(Iff98739de575e25104c0dc30f08912a5);
            Ibceb2b824cd4bc10bb06ee8adc693bd1    = I5c523df1fb2161ab4efd1c9b3e6b7aef;

            I1952614b64ea451e9d0646dcce5dd1cd = I914cb87eba8baa40cd515334e59f26b2 + ~I06e05a1ed002175a75d02b8b76f52c50 + 1;
            Ia307e5901694783f7761cdf724b767d0 = I2bcab411f9bec1541259751bcb9e0823(I1952614b64ea451e9d0646dcce5dd1cd);
            Ia8b9f373fe68ac4cbca35e04376e3cca    = Ia307e5901694783f7761cdf724b767d0;

            I49c1a7d1c20a25496821ad80c7eff790 = I914cb87eba8baa40cd515334e59f26b2 + ~I894ef04bfa1b7b39ef51b7c82f7686eb + 1;
            Ia47164e8ba831b85e696e30ff59ceab1 = I2bcab411f9bec1541259751bcb9e0823(I49c1a7d1c20a25496821ad80c7eff790);
            I5d1a89e85f6609b469e73e15aeffcbc4    = Ia47164e8ba831b85e696e30ff59ceab1;

            Ie2be17a55e79ca76350e033f227800de = I914cb87eba8baa40cd515334e59f26b2 + ~Id2989aaee3930698cd374e6c9feedf82 + 1;
            Ic217af0cb9728801034fdcb273a577fc = I2bcab411f9bec1541259751bcb9e0823(Ie2be17a55e79ca76350e033f227800de);
            I677fe06bad241bc8dd6a65a97f6db520    = Ic217af0cb9728801034fdcb273a577fc;

            I737a5b06f848cacf0c8da4985c73c66b = I914cb87eba8baa40cd515334e59f26b2 + ~I8487a819dcb61016798cde56f9662fcf + 1;
            Id5c8ea61025914f6e5a9b5eab9269261 = I2bcab411f9bec1541259751bcb9e0823(I737a5b06f848cacf0c8da4985c73c66b);
            If3c0f892fd71eb0ed8d1f70b4b33450b    = Id5c8ea61025914f6e5a9b5eab9269261;

            Iab160609bb21501aa55b662d2010357b = I32ed679af4ab759901aee43c9d93eb67 + ~Ic9678deca4bf44a7b99f853334f6a05c + 1;
            I924ef8499a83579e3449bbac0994775e = I2bcab411f9bec1541259751bcb9e0823(Iab160609bb21501aa55b662d2010357b);
            Ic65f0f75f56bf85122a89cdf07e98152    = I924ef8499a83579e3449bbac0994775e;

            Ief74f1a9d4a43ee5c9def7b83369bb21 = I32ed679af4ab759901aee43c9d93eb67 + ~I83b77ad1a40dc102f28153f692516eb4 + 1;
            Ia8da4833c93e9ef6188709e7082092de = I2bcab411f9bec1541259751bcb9e0823(Ief74f1a9d4a43ee5c9def7b83369bb21);
            I41d22bafaf58e4a6de04640864653a16    = Ia8da4833c93e9ef6188709e7082092de;

            Id144423f50751e661db3860a8487d004 = I32ed679af4ab759901aee43c9d93eb67 + ~I920f95bb52cdc9b07f93afc3a6b5c009 + 1;
            Icd8516e6bf231bce29ebefbc7c97bff7 = I2bcab411f9bec1541259751bcb9e0823(Id144423f50751e661db3860a8487d004);
            I06a46b86f6edede0f5f72658a19910b7    = Icd8516e6bf231bce29ebefbc7c97bff7;

            I623352a4f6705b21d461d6b32e85c12b = I32ed679af4ab759901aee43c9d93eb67 + ~I8d07beccef519ab4ce4024d911ac2346 + 1;
            I76c6762c515d0c9de1d777c0868b20af = I2bcab411f9bec1541259751bcb9e0823(I623352a4f6705b21d461d6b32e85c12b);
            I8591d0399594adacfeb006c5195c2c71    = I76c6762c515d0c9de1d777c0868b20af;

            I28d1dc8dc594977b5058b5bb9f6bfc66 = I32ed679af4ab759901aee43c9d93eb67 + ~Ia2904a5d5db43a209bd4b358ace68c6a + 1;
            If5da296bcf91d370f8341fc402eed6df = I2bcab411f9bec1541259751bcb9e0823(I28d1dc8dc594977b5058b5bb9f6bfc66);
            Id90588b5f82cd32e801fbea04d24e4a5    = If5da296bcf91d370f8341fc402eed6df;

            I5371a83bf9d6f334cf8d1c5b082527e9 = Id376dfa5141402f4d41a8858180ed87e + ~Ia209e5b03deaf4fcb8ae12b731a49e0a + 1;
            I64673b4b013682f9ce54925853c06ca4 = I2bcab411f9bec1541259751bcb9e0823(I5371a83bf9d6f334cf8d1c5b082527e9);
            Ib642d757fae818cd6d713ffb6ce18fc1    = I64673b4b013682f9ce54925853c06ca4;

            If1605d6646fd267e701668a7245b3b44 = Id376dfa5141402f4d41a8858180ed87e + ~Id2e223005a932987b6f60663773187f8 + 1;
            Iabfccf7b60f9be4e3714ad753cd8922a = I2bcab411f9bec1541259751bcb9e0823(If1605d6646fd267e701668a7245b3b44);
            Id76bff2a12cf792e52ccc463647334c0    = Iabfccf7b60f9be4e3714ad753cd8922a;

            Idf5eb1ac2c5bd92fa08ed935ae298255 = Id376dfa5141402f4d41a8858180ed87e + ~Ia8b29ca047a643f47bd3a0ffb50bf8cb + 1;
            I73ab1f85232818929b1b2e9d343584a3 = I2bcab411f9bec1541259751bcb9e0823(Idf5eb1ac2c5bd92fa08ed935ae298255);
            I92ffa890ed6d83d4fc543504e4d421c1    = I73ab1f85232818929b1b2e9d343584a3;

            I44ce30330c4d2d6033a0a970dd2bdd68 = I98a384bc62ee03f5ad7df20ef2d9af95 + ~I99d236d41be79090ca7ba1fb6faaec4c + 1;
            I06f989f65e614903ffba3594e8112235 = I2bcab411f9bec1541259751bcb9e0823(I44ce30330c4d2d6033a0a970dd2bdd68);
            Ifc4a65edeaf630b3d29437bcd6c20121    = I06f989f65e614903ffba3594e8112235;

            Ic101b8f56ea1e25c6b752583a1b01242 = I98a384bc62ee03f5ad7df20ef2d9af95 + ~Ia92b76ee5b7d82a992a1b58147c0c0be + 1;
            I0391247480cb6bd6bda2c59dcf8f7607 = I2bcab411f9bec1541259751bcb9e0823(Ic101b8f56ea1e25c6b752583a1b01242);
            Id57a11f56fc223501a9b68b8b05ebd3e    = I0391247480cb6bd6bda2c59dcf8f7607;

            Ib7cf44e681881e55d2d353280a6319d6 = I98a384bc62ee03f5ad7df20ef2d9af95 + ~Ic45d0537b94bc30713c0a0ee07b1ec40 + 1;
            Iee114a92d2238e4b8fcdfa79c4c99d6a = I2bcab411f9bec1541259751bcb9e0823(Ib7cf44e681881e55d2d353280a6319d6);
            I522ba8bfc1949337e8befe82cc1e86e6    = Iee114a92d2238e4b8fcdfa79c4c99d6a;

            I35690f724e964248dbb1e80fb1ea49f8 = Icfed259ca2bb2732d8e0c26ef67cd4cf + ~I26ae9e570a101c6f8237d7941285b924 + 1;
            Ida429b8e252b80b45435af1c6522f783 = I2bcab411f9bec1541259751bcb9e0823(I35690f724e964248dbb1e80fb1ea49f8);
            I7153e27c44ebbc2f04e9ba03cf09b5e1    = Ida429b8e252b80b45435af1c6522f783;

            I5affa2759148a6baf5b9f0cd3122348c = Icfed259ca2bb2732d8e0c26ef67cd4cf + ~Idcd5283cf7b42d403ee0e4404b5b311b + 1;
            Id3849d43e39d78fd2428109bf9677e0d = I2bcab411f9bec1541259751bcb9e0823(I5affa2759148a6baf5b9f0cd3122348c);
            Id15e4b4f186ec863f12a54acd8ef8963    = Id3849d43e39d78fd2428109bf9677e0d;

            Iaeea1f06ff0c6e9cfa43ba14420c3adc = Icfed259ca2bb2732d8e0c26ef67cd4cf + ~I337231f0dc7eb85f7d950262e0adb724 + 1;
            I5e51799e585f3dbef5e64908bcfc3e7a = I2bcab411f9bec1541259751bcb9e0823(Iaeea1f06ff0c6e9cfa43ba14420c3adc);
            I95c77eec7575cd7aa93a36f31ea635a2    = I5e51799e585f3dbef5e64908bcfc3e7a;

            Iac5a23266c3b038b4b54a916dccdf3a8 = I20861535c450d6e6bf11c45dac120454 + ~Iabe5aea929c668c9b9728d073ffb00c8 + 1;
            I6d12e4545b8befb8d09545ea00c8ea96 = I2bcab411f9bec1541259751bcb9e0823(Iac5a23266c3b038b4b54a916dccdf3a8);
            I3c8114dbe0658cc2889c787f1366abfa    = I6d12e4545b8befb8d09545ea00c8ea96;

            Icdfb7f52cc27b1cfcde90a100d29af13 = I20861535c450d6e6bf11c45dac120454 + ~Id201f81bbd80a70006a10866b8efeeff + 1;
            I98d04e6bae91796784a864c5bed637cb = I2bcab411f9bec1541259751bcb9e0823(Icdfb7f52cc27b1cfcde90a100d29af13);
            Ieacf971e9e10fb73c7df9f1da8372f30    = I98d04e6bae91796784a864c5bed637cb;

            I71484d7e00efa02a08b54a1405f2902c = I20861535c450d6e6bf11c45dac120454 + ~I530cf1f747d1df44b913f49eee90c079 + 1;
            I83b3247bed67d1e2ed488d5b7812851d = I2bcab411f9bec1541259751bcb9e0823(I71484d7e00efa02a08b54a1405f2902c);
            I35de1b03ea865f2c6381ce73e03dc220    = I83b3247bed67d1e2ed488d5b7812851d;

            I68a9b0607e69e8b3dae64689eb288a33 = I013929385ad819ddfcfcc59c22902ee3 + ~I1240c9410b897a4d0504affca5ba139e + 1;
            I868021f44830a9d81c4ba3dad804f889 = I2bcab411f9bec1541259751bcb9e0823(I68a9b0607e69e8b3dae64689eb288a33);
            Idec12e02904ea98c7580919584f2dba1    = I868021f44830a9d81c4ba3dad804f889;

            I2598c48aad48072a7f216b2ab56ee532 = I013929385ad819ddfcfcc59c22902ee3 + ~I4f169c2c8c0768f2725ed655a03acfc2 + 1;
            I685e59e3865058f29978a8cc2f1b6c7c = I2bcab411f9bec1541259751bcb9e0823(I2598c48aad48072a7f216b2ab56ee532);
            Ia370c83631a2c1bbf39c7264deafafb5    = I685e59e3865058f29978a8cc2f1b6c7c;

            I796e3a193b1b66fa9a04ca60aee11ea1 = I013929385ad819ddfcfcc59c22902ee3 + ~I342a563de39175fe4a6eb7e3e1ccac9a + 1;
            I5a76dd9f4a2078dee81102a9f205ca53 = I2bcab411f9bec1541259751bcb9e0823(I796e3a193b1b66fa9a04ca60aee11ea1);
            I05b4a07dfc0d2695eae34bea4c1c6565    = I5a76dd9f4a2078dee81102a9f205ca53;

            Ic96be7e69faf0f43b92618131cf0c98a = I013929385ad819ddfcfcc59c22902ee3 + ~Ief52461e4a5ddb128be5e439edf34862 + 1;
            Ice3bd7a4bbf0705a3dc1f89c5ceca084 = I2bcab411f9bec1541259751bcb9e0823(Ic96be7e69faf0f43b92618131cf0c98a);
            If1ecdc27e3419dd1434e403f237c2b58    = Ice3bd7a4bbf0705a3dc1f89c5ceca084;

            I648afe4114ce435bf1d13e0ad54425cf = I34fffcb07fe82f11fe142f7c37f39155 + ~I015630502f5cb4eb27b2a673e810f1dc + 1;
            I5f741a3213cecdf58440120c2ea78e87 = I2bcab411f9bec1541259751bcb9e0823(I648afe4114ce435bf1d13e0ad54425cf);
            I039c552777d0fb40bebcdd2d4a3394c2    = I5f741a3213cecdf58440120c2ea78e87;

            If05d7e30b4717e0a1bfd20b90d0539bd = I34fffcb07fe82f11fe142f7c37f39155 + ~I8bb46c3eb9f54c5d1b28dc6aa0154358 + 1;
            Idad89ade7f96091abfea876b3af0d5b4 = I2bcab411f9bec1541259751bcb9e0823(If05d7e30b4717e0a1bfd20b90d0539bd);
            Iaa52fb63184514b6d754bcc896235150    = Idad89ade7f96091abfea876b3af0d5b4;

            I5fc356af8a62a1d739cb375fb851e90f = I34fffcb07fe82f11fe142f7c37f39155 + ~I938dd59e4cdf3434086f60d000113430 + 1;
            Ie0ab4b7c79196195db0971e7c7a85adb = I2bcab411f9bec1541259751bcb9e0823(I5fc356af8a62a1d739cb375fb851e90f);
            Ied9781e625c1fa8741853dd6b8b3a9e7    = Ie0ab4b7c79196195db0971e7c7a85adb;

            I22f4c5403fbe33d18f97cf21786cdd80 = I34fffcb07fe82f11fe142f7c37f39155 + ~I46d86bfa6de26f3cfef9d802549ef2ad + 1;
            I0093585d710940feaa8ebdc5fb000806 = I2bcab411f9bec1541259751bcb9e0823(I22f4c5403fbe33d18f97cf21786cdd80);
            I767272262e9d2e85dba1aa93f578f25c    = I0093585d710940feaa8ebdc5fb000806;

            I9a1b2b9f924099f1e57fa501ba2e33ba = I61ca60fde05ed88cce714dcd8c13b827 + ~Iff1d4b06901796098f91e87a3c30f7a5 + 1;
            I76a0b74bb633743ac56cf4a0d52f80c0 = I2bcab411f9bec1541259751bcb9e0823(I9a1b2b9f924099f1e57fa501ba2e33ba);
            Ib3b4cd6d8ab17869a2278552c02635c8    = I76a0b74bb633743ac56cf4a0d52f80c0;

            If6253af4ebc430e4937269a5f4989b29 = I61ca60fde05ed88cce714dcd8c13b827 + ~I1e110e27162231650875dd1152d96e64 + 1;
            I11931fd13219c1ae615d164a8f4130f9 = I2bcab411f9bec1541259751bcb9e0823(If6253af4ebc430e4937269a5f4989b29);
            Ie7a5cb2ecb3fce35825785b9bca6b3bd    = I11931fd13219c1ae615d164a8f4130f9;

            I0427d17423548dbb33cf792883b4be8c = I61ca60fde05ed88cce714dcd8c13b827 + ~Ie7274a7ffa053ced4f12a67986d3c81b + 1;
            I6de7a344ae1574e551c7c10a1773d880 = I2bcab411f9bec1541259751bcb9e0823(I0427d17423548dbb33cf792883b4be8c);
            Ib9a0f8efd3dad427f247ce90fdfb94a4    = I6de7a344ae1574e551c7c10a1773d880;

            Ie539faf01ae85253e399308fef98afd6 = I61ca60fde05ed88cce714dcd8c13b827 + ~If6a3bd6f002d91e0773c4ab9caaaa01e + 1;
            I4920b0740cb56988ba4fc10b86195cdd = I2bcab411f9bec1541259751bcb9e0823(Ie539faf01ae85253e399308fef98afd6);
            I69a221a1bd95a588aa74b9bed0357762    = I4920b0740cb56988ba4fc10b86195cdd;

            Iae6e7c42f250cd9223f18f8830fb177d = I4907dd45c158dc7e0041c64f1fb388f6 + ~I54c260db5c1b2c76527c8fc1cee229fe + 1;
            I37d27fda03770ad37a1fbad835c076c3 = I2bcab411f9bec1541259751bcb9e0823(Iae6e7c42f250cd9223f18f8830fb177d);
            I64f125cf2ca6a6da8a9cdae9e246c24a    = I37d27fda03770ad37a1fbad835c076c3;

            Iff47ec1743b59d7f90e9042af7ce44cb = I4907dd45c158dc7e0041c64f1fb388f6 + ~I55e54359961ef6e5a63f1c2eb0ad4aa1 + 1;
            Ib868fcb71300c09a49719e0b0459ca06 = I2bcab411f9bec1541259751bcb9e0823(Iff47ec1743b59d7f90e9042af7ce44cb);
            Ifac9dd60dd6c543aa94b39c599f0819a    = Ib868fcb71300c09a49719e0b0459ca06;

            I1cf4a55ebab332defa32d2922b885285 = I4907dd45c158dc7e0041c64f1fb388f6 + ~I4f38c3d620b72f21cf6d54c7df4ba816 + 1;
            I2c67e89b58d7f998c43c68d857fa2381 = I2bcab411f9bec1541259751bcb9e0823(I1cf4a55ebab332defa32d2922b885285);
            Icf062382a1e462571569ccee75b0a3ee    = I2c67e89b58d7f998c43c68d857fa2381;

            I284913858691ad5724073b73a820047a = I4907dd45c158dc7e0041c64f1fb388f6 + ~Ib33e1c6d57e5e6fc465dc9c9a7cf29fa + 1;
            Idb770d9fc630f77beca27c3182279001 = I2bcab411f9bec1541259751bcb9e0823(I284913858691ad5724073b73a820047a);
            Ieed8b94295bed265961c4f52c3379914    = Idb770d9fc630f77beca27c3182279001;

            I35626ca53adbbf0a3a71cc6fcf43bcb1 = I2c8f6a9b9f655b317bb0af4d60fdbc4b + ~I3a8bcfdab631a268d21c87b98e9d1c49 + 1;
            I6ab74c183d97a5df7a336c6c66c66e2e = I2bcab411f9bec1541259751bcb9e0823(I35626ca53adbbf0a3a71cc6fcf43bcb1);
            I165eabcdde76821fdc308ff7a8c6d2ea    = I6ab74c183d97a5df7a336c6c66c66e2e;

            I0d74ef22d31abcec73c7c582310b1e6d = I2c8f6a9b9f655b317bb0af4d60fdbc4b + ~Iad0ecc5208263d239e4a62c5563f52ab + 1;
            Ic4fc6d6a69dccb796d208aba87ec002c = I2bcab411f9bec1541259751bcb9e0823(I0d74ef22d31abcec73c7c582310b1e6d);
            I8b3542a6d64d6a7ebba4124bc6702f3e    = Ic4fc6d6a69dccb796d208aba87ec002c;

            I15f4cf1aa0ad5ce2bda52df338e677e3 = I2c8f6a9b9f655b317bb0af4d60fdbc4b + ~Ic0b2f9717b8aacb34325fd5aaf03a366 + 1;
            I450cd05f0109ad62ae4ca7f540ac7505 = I2bcab411f9bec1541259751bcb9e0823(I15f4cf1aa0ad5ce2bda52df338e677e3);
            I7b68afec199be705d766c169f1ece981    = I450cd05f0109ad62ae4ca7f540ac7505;

            I6c5ca5e68c8844bb1617a2288b5bbc37 = I2c8f6a9b9f655b317bb0af4d60fdbc4b + ~Id92a319da408be46970faf524513fdd8 + 1;
            Ia6f1bdee90a01ee3f3e59eec00689d50 = I2bcab411f9bec1541259751bcb9e0823(I6c5ca5e68c8844bb1617a2288b5bbc37);
            I4b6c8226ef2bc20dbd31d242bdb98b8c    = Ia6f1bdee90a01ee3f3e59eec00689d50;

            I44343a9491069c3c8ea4fbd6255a5a6c = Ic7dff631559304ec59f0696c66436d62 + ~I95b923444062b4a98918c685c65996d0 + 1;
            I33193403a8d72dcd02e87ae03b668e09 = I2bcab411f9bec1541259751bcb9e0823(I44343a9491069c3c8ea4fbd6255a5a6c);
            Ic3b4a86f22caf5b6103d52b6c9d2a991    = I33193403a8d72dcd02e87ae03b668e09;

            I1d8318b94d86e1fd28323a5e5684a37b = Ic7dff631559304ec59f0696c66436d62 + ~I06c0921675f464807a63c7965796f0d0 + 1;
            I5208f3202b32a30c4abaca4c617d3b3b = I2bcab411f9bec1541259751bcb9e0823(I1d8318b94d86e1fd28323a5e5684a37b);
            Ia37592b207086f63e2d94e3d7d26c740    = I5208f3202b32a30c4abaca4c617d3b3b;

            I825e83bd88575868f4fcc9a8b8729663 = Ic7dff631559304ec59f0696c66436d62 + ~I59adad4fd84c1fc233dc58f70a12779d + 1;
            Ib607167c806dd831aaed4a42b9cf4349 = I2bcab411f9bec1541259751bcb9e0823(I825e83bd88575868f4fcc9a8b8729663);
            Id0d786026e3ab0ddbffbc20e4d409857    = Ib607167c806dd831aaed4a42b9cf4349;

            I3184a16c71cff80c8c90b40e45f114b8 = Ic7dff631559304ec59f0696c66436d62 + ~Iae182ffae6cea89363f0ccc8b5679561 + 1;
            I42b87e52c168abb775c1e1e5ddfc1958 = I2bcab411f9bec1541259751bcb9e0823(I3184a16c71cff80c8c90b40e45f114b8);
            I333837f976cfc7f90ab0a6dcd8c1ce79    = I42b87e52c168abb775c1e1e5ddfc1958;

            Iae133550f8bad8357a73e7de1372faa3 = I6a239d3e55b4a9a3be9989a85bbec545 + ~Ie40c90fdb38b3e4046ba89295ed77d7c + 1;
            Ifc4e50801a1606717efd57bd5ac6f41f = I2bcab411f9bec1541259751bcb9e0823(Iae133550f8bad8357a73e7de1372faa3);
            Id115b4708a49dcfd167e79ef6993e371    = Ifc4e50801a1606717efd57bd5ac6f41f;

            Ibccb4a43c410f698e0fff68553326a77 = I6a239d3e55b4a9a3be9989a85bbec545 + ~I13b9e098622d90a1074f636d8f351aca + 1;
            I5e7282e9a35cead2f4d1d9860d45852c = I2bcab411f9bec1541259751bcb9e0823(Ibccb4a43c410f698e0fff68553326a77);
            I666da645400344644e848ee6f7592d3c    = I5e7282e9a35cead2f4d1d9860d45852c;

            I72dc7aa294a3af89101ea62a4223170e = I6a239d3e55b4a9a3be9989a85bbec545 + ~I1972375d51767f0cffa5395a354b3493 + 1;
            I8503b90594f3d4b492cca9cf154fc3d3 = I2bcab411f9bec1541259751bcb9e0823(I72dc7aa294a3af89101ea62a4223170e);
            Ibafeadd691eee03f855ed657c01022c9    = I8503b90594f3d4b492cca9cf154fc3d3;

            I91eb3e70921e0b141a344bc57dfbc934 = I6a239d3e55b4a9a3be9989a85bbec545 + ~Idfe6aecb694385ce8c3c1544a4992a20 + 1;
            I95010cdf08c373916ab02e3794afa77a = I2bcab411f9bec1541259751bcb9e0823(I91eb3e70921e0b141a344bc57dfbc934);
            I10ec5c43a3fb65273053063001307280    = I95010cdf08c373916ab02e3794afa77a;

            I1986f22f2269cc135c6ed28d35fb0bd1 = I630f905e55f08e7d1569a08e937ad216 + ~I9859b94cda465ceaaa5674eb19e94824 + 1;
            I832fdc71e665ad2acac2576188e0d65b = I2bcab411f9bec1541259751bcb9e0823(I1986f22f2269cc135c6ed28d35fb0bd1);
            I05c778eb3588bdaccf714ba456f534c2    = I832fdc71e665ad2acac2576188e0d65b;

            Ibef24017bc71de9c002aafa7ce9a784c = I630f905e55f08e7d1569a08e937ad216 + ~I8d6927b0bcbbb318cf52987c121a07b5 + 1;
            Ic21a6f1abcecf14acaf2aa23b7dcdb6b = I2bcab411f9bec1541259751bcb9e0823(Ibef24017bc71de9c002aafa7ce9a784c);
            Icd11e8d97a6ac6c0a73e8adee1f98c4e    = Ic21a6f1abcecf14acaf2aa23b7dcdb6b;

            Ieae3ed78fa2c45507066f4e20d96e956 = I630f905e55f08e7d1569a08e937ad216 + ~Ide40b1bf9c0b642c49a5685a62af1c93 + 1;
            I49847c8c979d9ed82be80f62552e97bf = I2bcab411f9bec1541259751bcb9e0823(Ieae3ed78fa2c45507066f4e20d96e956);
            If07c2223d4262e22cca9b77c3ed5ee01    = I49847c8c979d9ed82be80f62552e97bf;

            I730fd25ffc7778fd4bb02d33cb3870d6 = I630f905e55f08e7d1569a08e937ad216 + ~Idfbc5726963cfa31bb4324143ffd08c7 + 1;
            I7a2bfe5efbe1d0dc222bff675c621485 = I2bcab411f9bec1541259751bcb9e0823(I730fd25ffc7778fd4bb02d33cb3870d6);
            If0c8ce0ff66fe2806448f1c819d58ec8    = I7a2bfe5efbe1d0dc222bff675c621485;

            I9a32313f2911b797fb0848f7d97e62b9 = I8d13eb3669785c4279c685763d4f3fad + ~I5085f161323433d8d38be2e4511b0c46 + 1;
            Ie0d874ce4b0713de7d087396a1879c54 = I2bcab411f9bec1541259751bcb9e0823(I9a32313f2911b797fb0848f7d97e62b9);
            Iccdc2371dfd9fda3e506adc2b1681ba3    = Ie0d874ce4b0713de7d087396a1879c54;

            I6373e2d64fdb5dd77733b3e4bb405121 = I8d13eb3669785c4279c685763d4f3fad + ~Ib66b897398ea0702b74bdd03774f3ae4 + 1;
            Iaf4c12394552f42e476b70f6c75003d7 = I2bcab411f9bec1541259751bcb9e0823(I6373e2d64fdb5dd77733b3e4bb405121);
            I26e61dca9d045c4661b97afe346152c8    = Iaf4c12394552f42e476b70f6c75003d7;

            Ib437aa67ab7c13b45d7a4d56ce9e79b8 = I8d13eb3669785c4279c685763d4f3fad + ~Ic227f42a20219c6638ee3343ca445acf + 1;
            I64d7f4a0df87ce07ce49350610122f79 = I2bcab411f9bec1541259751bcb9e0823(Ib437aa67ab7c13b45d7a4d56ce9e79b8);
            Id488d650b86f5def0668f4a1ef841b6a    = I64d7f4a0df87ce07ce49350610122f79;

            I0cb5c7a759f4c75d4a675f9777f15c5f = I8d13eb3669785c4279c685763d4f3fad + ~I205d5fdeae55fae7be2f06f11c949244 + 1;
            If51795ea140bec96fdefbc52291801b5 = I2bcab411f9bec1541259751bcb9e0823(I0cb5c7a759f4c75d4a675f9777f15c5f);
            I479365266255d2228ecd86c350e8d38b    = If51795ea140bec96fdefbc52291801b5;

            I0ca91c1426ba14a7b47a081cb3becd19 = I25a6f3de9a9a01cbbdd32ed848561aa4 + ~I16db9cab1981451a02dab21e2ca221b4 + 1;
            Ib0a0f80cb818018b2fe0fd4597325bb4 = I2bcab411f9bec1541259751bcb9e0823(I0ca91c1426ba14a7b47a081cb3becd19);
            I08d9c488fd85db45344e649699196263    = Ib0a0f80cb818018b2fe0fd4597325bb4;

            I0737e0cc7453e328efab2277bb712ea8 = I25a6f3de9a9a01cbbdd32ed848561aa4 + ~Idc758f8e6fabb6b31b0a7d9c0c590310 + 1;
            If01a65e097f026a816133c34d73ccff1 = I2bcab411f9bec1541259751bcb9e0823(I0737e0cc7453e328efab2277bb712ea8);
            Icde86d0ead44385b07e9a29057417417    = If01a65e097f026a816133c34d73ccff1;

            I456af863661122cc303fccb235f3c7a1 = I25a6f3de9a9a01cbbdd32ed848561aa4 + ~I3188d354c2ba494ffe210dcd89c00620 + 1;
            Ida9ed61c543afde2257053443d133119 = I2bcab411f9bec1541259751bcb9e0823(I456af863661122cc303fccb235f3c7a1);
            I21feecd24d912ef3d0aec0e375958f3f    = Ida9ed61c543afde2257053443d133119;

            Idc5916c4800e9f647d51c52444ab6fff = I25a6f3de9a9a01cbbdd32ed848561aa4 + ~Ie667e1755ae1561a2eefae9b63845dec + 1;
            I983a5656d68192a7a3d5a78f17f12ff0 = I2bcab411f9bec1541259751bcb9e0823(Idc5916c4800e9f647d51c52444ab6fff);
            I59f419b3bc183a5fe743be3878fac587    = I983a5656d68192a7a3d5a78f17f12ff0;

            I57aca70e2b8d126c120736b2606ed333 = Iba3dd4b2c2c85c4cfe770d9b52ef4634 + ~I3d700e050cb7f22b0e381f3c72a20124 + 1;
            I315445ad2d762b66f94a75d76fbfb839 = I2bcab411f9bec1541259751bcb9e0823(I57aca70e2b8d126c120736b2606ed333);
            Ib0804d8bdda49ecd0024300eed52be53    = I315445ad2d762b66f94a75d76fbfb839;

            Ic6650a6d092b749b4498c08d69cf815e = Iba3dd4b2c2c85c4cfe770d9b52ef4634 + ~Idc198bd5732ca5760d1a700a25273ce3 + 1;
            I7a97a8fe65e56b0a80c242e13e70db09 = I2bcab411f9bec1541259751bcb9e0823(Ic6650a6d092b749b4498c08d69cf815e);
            I37b0efdee34647a5111d698a5a80f367    = I7a97a8fe65e56b0a80c242e13e70db09;

            Ic2e3b8f91eb218650c7b9c515c7efe97 = Iba3dd4b2c2c85c4cfe770d9b52ef4634 + ~I2253b32e46200a23dba243819fce02f0 + 1;
            I2243095f420e4d996f1c69c965932778 = I2bcab411f9bec1541259751bcb9e0823(Ic2e3b8f91eb218650c7b9c515c7efe97);
            Id382a04e94d0749d0858041bdc5861be    = I2243095f420e4d996f1c69c965932778;

            I93a084aa1e6881ab8dc905dcdcdfd7ee = Iba3dd4b2c2c85c4cfe770d9b52ef4634 + ~If7348fdbe0400aab92e8fd6a7cf6c267 + 1;
            I0154a19f9adb43089080304978256c09 = I2bcab411f9bec1541259751bcb9e0823(I93a084aa1e6881ab8dc905dcdcdfd7ee);
            I368be992a21201268c41506396dcdcf6    = I0154a19f9adb43089080304978256c09;

            I8cba172573be52c5a90bd40e6f40a508 = Ie1b744387b5200a504e4874e14d2f282 + ~If17b4f86674bc5fb212a1f7751fb043a + 1;
            Ib8bdc3b41b3cc7132c43833802115880 = I2bcab411f9bec1541259751bcb9e0823(I8cba172573be52c5a90bd40e6f40a508);
            I603a008893b5196d9f273b47a9d63144    = Ib8bdc3b41b3cc7132c43833802115880;

            I1cccfd1516af59265731121dde878116 = Ie1b744387b5200a504e4874e14d2f282 + ~Ife7985db888089ea618413810611bfca + 1;
            I167586906b601ffc473a5b856b213f2b = I2bcab411f9bec1541259751bcb9e0823(I1cccfd1516af59265731121dde878116);
            Ie70d3a768bc09ddff6ac68aaba7d9f2c    = I167586906b601ffc473a5b856b213f2b;

            Ia171bbefe2d20b4c058126c33ef28eb8 = Ie1b744387b5200a504e4874e14d2f282 + ~Ia020344403aad35e050765a4b0cc42b7 + 1;
            I094a6ac91aacfdd2f8de8a0d776f732b = I2bcab411f9bec1541259751bcb9e0823(Ia171bbefe2d20b4c058126c33ef28eb8);
            Ifb8bd837ada3d8ed5116db29da82d2a9    = I094a6ac91aacfdd2f8de8a0d776f732b;

            I84bc44a5d53a8f66b985b70c7ec1ae7c = Ie1b744387b5200a504e4874e14d2f282 + ~I143b91852fddcdcc30bf1041332c4ed7 + 1;
            I9d4437c250c28653bbccdea6af8b6280 = I2bcab411f9bec1541259751bcb9e0823(I84bc44a5d53a8f66b985b70c7ec1ae7c);
            I978b93d46e20cb3eda70e5a976d62348    = I9d4437c250c28653bbccdea6af8b6280;

            I321b104ca3c818018d4b03adfe1110b9 = Icf76cb69aedf4db01cd3444f4c4ba471 + ~I4fb3fe065daa2708e55c812e57c19fb6 + 1;
            I4afab82ea1a6ad0a36fea0692de1d106 = I2bcab411f9bec1541259751bcb9e0823(I321b104ca3c818018d4b03adfe1110b9);
            Ib404040d4fb58f47f245184c3be01789    = I4afab82ea1a6ad0a36fea0692de1d106;

            Ia79b8994da536c86634bf6f54a21145d = Icf76cb69aedf4db01cd3444f4c4ba471 + ~I96f65790e2cacf7b529ce5b88598da00 + 1;
            I864d41b77a51fda97ea7017ed18b5fea = I2bcab411f9bec1541259751bcb9e0823(Ia79b8994da536c86634bf6f54a21145d);
            I9c664265c53ebffaad097b70ff3cbbce    = I864d41b77a51fda97ea7017ed18b5fea;

            I4df55ce80eec5fee295b5a0ae92bd6c8 = Icf76cb69aedf4db01cd3444f4c4ba471 + ~If077c67a062095cfe69f2260cee82833 + 1;
            I758ee12b430cda151b452699eb2039dc = I2bcab411f9bec1541259751bcb9e0823(I4df55ce80eec5fee295b5a0ae92bd6c8);
            I781306c6b1ce0741d9c2fa06865f7a19    = I758ee12b430cda151b452699eb2039dc;

            I46593a7956590d870fe680228081a6d2 = Icf76cb69aedf4db01cd3444f4c4ba471 + ~Iee5e74945ba15220f0f707c9c1927ba1 + 1;
            I134cd61326b70030c027a3821d98a994 = I2bcab411f9bec1541259751bcb9e0823(I46593a7956590d870fe680228081a6d2);
            I16fa2e3dc0b3eddbc72811b51d6ac8ed    = I134cd61326b70030c027a3821d98a994;

            I906e9da31de73ae45579607a014e8b54 = I4857b5b50556c8e7fff4b2d3e08e4b28 + ~Iffb7fe9c74dfc01a43e99a099c4e7e04 + 1;
            I99951d295b9065614c103b3e43fa255c = I2bcab411f9bec1541259751bcb9e0823(I906e9da31de73ae45579607a014e8b54);
            Ia6f232495726806d01b702b0e248b2f2    = I99951d295b9065614c103b3e43fa255c;

            If5dd1a1b9e3fc0e67a85da3183480aed = I4857b5b50556c8e7fff4b2d3e08e4b28 + ~Ic09b4671e867144fe9f54a09e74c5519 + 1;
            I31a4e4f3eac271c84b36c84d7de338fd = I2bcab411f9bec1541259751bcb9e0823(If5dd1a1b9e3fc0e67a85da3183480aed);
            I66b3734060600caa45d699508c5083d2    = I31a4e4f3eac271c84b36c84d7de338fd;

            Iadfb1571c78c3f0c05e4ef498267df24 = I4857b5b50556c8e7fff4b2d3e08e4b28 + ~Ic0ae1191869e636f9e4391efe93309ae + 1;
            Id36c36d2b2dd9a79f9887c9950b385c3 = I2bcab411f9bec1541259751bcb9e0823(Iadfb1571c78c3f0c05e4ef498267df24);
            I85fae6b23d086235a94a0162e2fb5310    = Id36c36d2b2dd9a79f9887c9950b385c3;

            Icebb43b184c2745cc9da9d01b06bc62f = I4857b5b50556c8e7fff4b2d3e08e4b28 + ~I4d1c47569b0bc8c651c897ac8e88bd1f + 1;
            I59455b0e53bac4fe6b1cbf609cb03da5 = I2bcab411f9bec1541259751bcb9e0823(Icebb43b184c2745cc9da9d01b06bc62f);
            I8d6443d1be42203cb834345ae7e5aff5    = I59455b0e53bac4fe6b1cbf609cb03da5;

            I6e4b0489ec7333abf2245a1b72a8923d = I0a1e9cf99f1d4725327615f50fcc3ad0 + ~I487b9b236d118786e475ccc5e4e56a6d + 1;
            Ifd633f2ea91cb88aaa2a0bf5579ed1e0 = I2bcab411f9bec1541259751bcb9e0823(I6e4b0489ec7333abf2245a1b72a8923d);
            I717332b7f76e9caf9351f1aa69b72a12    = Ifd633f2ea91cb88aaa2a0bf5579ed1e0;

            I24ac5dd30526c1d3bc7b941103a66804 = I0a1e9cf99f1d4725327615f50fcc3ad0 + ~Ic46357bb77f6183329946f7e28294365 + 1;
            I87218b174c1db735ac153604b5ff3e15 = I2bcab411f9bec1541259751bcb9e0823(I24ac5dd30526c1d3bc7b941103a66804);
            Ieebd34db071409288f489129b70ab599    = I87218b174c1db735ac153604b5ff3e15;

            I33681b2292c086fe536dae2aec70903a = I0a1e9cf99f1d4725327615f50fcc3ad0 + ~I382153cec6f7d6258574e7c532186473 + 1;
            I4608c92d52306432c114f31b9ba6dd69 = I2bcab411f9bec1541259751bcb9e0823(I33681b2292c086fe536dae2aec70903a);
            I917c874137d64a9a495335c8f8ef5374    = I4608c92d52306432c114f31b9ba6dd69;

            Ia373ca76c3b15a4148532b3822f82ba5 = I0a1e9cf99f1d4725327615f50fcc3ad0 + ~Ib9d6c5be487a434fbafcda25ca9351dc + 1;
            Iba3f6cde40827d82bc32078344b9bd81 = I2bcab411f9bec1541259751bcb9e0823(Ia373ca76c3b15a4148532b3822f82ba5);
            I15fb4fb838d4a614c468f7d49261bda3    = Iba3f6cde40827d82bc32078344b9bd81;

            I7d08adbaf66cea04be4891db610bca3f = Ie844f4c446983ce381b0bc4c0e8ef7d7 + ~Icb92c7c10f0bfc5d287228f98d8a235c + 1;
            Ib987bde3ee5a0256d0b8b3aa7357cdb2 = I2bcab411f9bec1541259751bcb9e0823(I7d08adbaf66cea04be4891db610bca3f);
            I2eb093d2a38ba8cf4be47d1d7f54ecc4    = Ib987bde3ee5a0256d0b8b3aa7357cdb2;

            Ic09ed51b20f411683a801eaad61657a3 = Ie844f4c446983ce381b0bc4c0e8ef7d7 + ~I90001da8c360ccff128f637cd672ad42 + 1;
            I3c33a2bfaa82172457b15f4f621eefee = I2bcab411f9bec1541259751bcb9e0823(Ic09ed51b20f411683a801eaad61657a3);
            I8f9affdc5cda0fecc35dd15fc5aeb244    = I3c33a2bfaa82172457b15f4f621eefee;

            I6a9af8c9009b5de47ebe9ee8b79d3831 = Ie844f4c446983ce381b0bc4c0e8ef7d7 + ~I5001118df37d08bd19d322aca8ff3996 + 1;
            I7ce33eb337b6cacaea13f748061e338a = I2bcab411f9bec1541259751bcb9e0823(I6a9af8c9009b5de47ebe9ee8b79d3831);
            I615a443d49d1479338d033d2a2cab51f    = I7ce33eb337b6cacaea13f748061e338a;

            Ife18e8a16d4437161b75a93e3dff1b5b = Ie844f4c446983ce381b0bc4c0e8ef7d7 + ~Ib0d033ba28e8c606ed92207049c76884 + 1;
            I7a8c5be75d87552ca717a87d1a832d21 = I2bcab411f9bec1541259751bcb9e0823(Ife18e8a16d4437161b75a93e3dff1b5b);
            I0635a3270a9653ca0f23c116fd5b2f97    = I7a8c5be75d87552ca717a87d1a832d21;

            I0cde86532c8db1a32d9fbe38a40b91b8 = I6067f47cccceea96ac46ff0d457b25f2 + ~I72756ea6a4997bc4afd4bfde1dfb2d26 + 1;
            Id9c9cebf44647040da33567d815c261f = I2bcab411f9bec1541259751bcb9e0823(I0cde86532c8db1a32d9fbe38a40b91b8);
            I93a7c75ebce8fbf4c613b4d11dc98b72    = Id9c9cebf44647040da33567d815c261f;

            I49c8ec4cd33e6caed8ed7dab779e7ebb = I6067f47cccceea96ac46ff0d457b25f2 + ~Iea4a7766d3b9d5d030ade1739859ef0d + 1;
            I6c522c28a0dc265facb1f21ebe51c564 = I2bcab411f9bec1541259751bcb9e0823(I49c8ec4cd33e6caed8ed7dab779e7ebb);
            I39334aa9d55bcc001ece37ce2a6c329c    = I6c522c28a0dc265facb1f21ebe51c564;

            Idb86f95570587a0711d796aac7004c25 = I6067f47cccceea96ac46ff0d457b25f2 + ~I78e1205de9119fac3ae8f43c72ac71f4 + 1;
            I86c367b0fd4548d5edfb8863f454653e = I2bcab411f9bec1541259751bcb9e0823(Idb86f95570587a0711d796aac7004c25);
            I07e328d23da9383a296ecb03679ec74b    = I86c367b0fd4548d5edfb8863f454653e;

            I2d1373d0b18992fa46a9607a86d21520 = I6067f47cccceea96ac46ff0d457b25f2 + ~I300d9f403e33d860ff5dde9f91bae11b + 1;
            I800271efe85fcbaee8fe733190e90f6d = I2bcab411f9bec1541259751bcb9e0823(I2d1373d0b18992fa46a9607a86d21520);
            I8a6e1eace6152af5c98c415804cb60fa    = I800271efe85fcbaee8fe733190e90f6d;

            I30f26e090ab14551cbac41883ad8a152 = Ifd6fd1f3cbf8884ca7f64bc42278e4fa + ~I63c0c8bef1dea4e499a16ce01e781951 + 1;
            Ia5172996abb4a6bc50046d36ec033c7f = I2bcab411f9bec1541259751bcb9e0823(I30f26e090ab14551cbac41883ad8a152);
            I6ed4d6c350e8691b3a12ab51419cfa65    = Ia5172996abb4a6bc50046d36ec033c7f;

            Ib1b4e41ab25733d1d6dd54e1fe81a419 = Ifd6fd1f3cbf8884ca7f64bc42278e4fa + ~I5a7746e9fbb8c009f83ae57423296cdf + 1;
            Ibe20363746d437eef2c85360425739d1 = I2bcab411f9bec1541259751bcb9e0823(Ib1b4e41ab25733d1d6dd54e1fe81a419);
            Ie2b9ed680dac51ac866cb830ca17ef84    = Ibe20363746d437eef2c85360425739d1;

            I146c0d5154a6de44c0536de873904ccf = Ifd6fd1f3cbf8884ca7f64bc42278e4fa + ~Ie0ce2826fd13b0e0b23c91e97787691f + 1;
            Iee695b22e8a55479dfcbaa68f5c8b6c9 = I2bcab411f9bec1541259751bcb9e0823(I146c0d5154a6de44c0536de873904ccf);
            Ie439b520bbb0c8b29a5ecea167acb1c9    = Iee695b22e8a55479dfcbaa68f5c8b6c9;

            I8eb9d4839a478a4e28b45a549b5682a4 = Ifd6fd1f3cbf8884ca7f64bc42278e4fa + ~Iebfe0fa45e4b34e142e82ddaa15243cf + 1;
            I7cdb0bf6c7195df38d701768e655af70 = I2bcab411f9bec1541259751bcb9e0823(I8eb9d4839a478a4e28b45a549b5682a4);
            I9f8ef3295578acf5b0a42d074a15a70b    = I7cdb0bf6c7195df38d701768e655af70;

            I2501ef991a59512c43693ba9d7db8571 = Iaec9fd9e79371676bfa8ff14b4feae52 + ~I275f6334127640b2de3f0f87f54fd74c + 1;
            I1057373671fd4cfba6696f8e88a2d740 = I2bcab411f9bec1541259751bcb9e0823(I2501ef991a59512c43693ba9d7db8571);
            Ief01b06341d489e36ee344fd52084ccf    = I1057373671fd4cfba6696f8e88a2d740;

            I38213f78fd4dc52f9d2c9b7b22136c1c = Iaec9fd9e79371676bfa8ff14b4feae52 + ~I3faeba79f7af7a006ab5cd256352e2db + 1;
            I7dd9da64c1516e6ae1b703defc4cdc55 = I2bcab411f9bec1541259751bcb9e0823(I38213f78fd4dc52f9d2c9b7b22136c1c);
            I3b72a085b104e17dca3d8b2824f84e97    = I7dd9da64c1516e6ae1b703defc4cdc55;

            I49ce91ac152279af421bbc6c4d9b8087 = Iaec9fd9e79371676bfa8ff14b4feae52 + ~I0c0be3347a7df9cc39997208b013f17b + 1;
            I58bf5f51208a98b2448e2b4fad3f63ac = I2bcab411f9bec1541259751bcb9e0823(I49ce91ac152279af421bbc6c4d9b8087);
            I5e1f41e23887493db1d723e1e2cbd996    = I58bf5f51208a98b2448e2b4fad3f63ac;

            I6a2b7bb2cb3ca2ab932c211a68dded55 = Iaec9fd9e79371676bfa8ff14b4feae52 + ~Ieb778442bc855e93e11c9b13f1a7ae06 + 1;
            Icb8281c05ea7168d39d6012a1d622e15 = I2bcab411f9bec1541259751bcb9e0823(I6a2b7bb2cb3ca2ab932c211a68dded55);
            I0e6f4c7bdc39bd22833f3d9fcfa55f1d    = Icb8281c05ea7168d39d6012a1d622e15;

            Idaae6ba9da8754615a2c34ef859492db = I500757c4eda5d3d899aee47b87da585b + ~Ie9fd8f7dc0c3849c0437a2a3d8607b4c + 1;
            I5b16ad2952938bc64f6c9f5ff1ab5a0b = I2bcab411f9bec1541259751bcb9e0823(Idaae6ba9da8754615a2c34ef859492db);
            Ie346802a8898b4b075be289e062b462c    = I5b16ad2952938bc64f6c9f5ff1ab5a0b;

            Icaca9fc70a3ec6c48c0e41f8168e2bb9 = I500757c4eda5d3d899aee47b87da585b + ~I45a6ef43e6e42594444adcbda26700ab + 1;
            I5d5790b480d08bf6c957f26e24467b9a = I2bcab411f9bec1541259751bcb9e0823(Icaca9fc70a3ec6c48c0e41f8168e2bb9);
            I82ea6f21706a97166ef11af548e80392    = I5d5790b480d08bf6c957f26e24467b9a;

            I4f69b8ff834c7ab3194bc9390ce0f5f6 = I500757c4eda5d3d899aee47b87da585b + ~If36016df78d833c80e1355151c038225 + 1;
            Ieb32ca618265eed3419f01907f48527d = I2bcab411f9bec1541259751bcb9e0823(I4f69b8ff834c7ab3194bc9390ce0f5f6);
            I5f38764f6ecc2dcd1fdd5316102f1f82    = Ieb32ca618265eed3419f01907f48527d;

            I037cb596cd48c5533ed22bc32518d992 = I500757c4eda5d3d899aee47b87da585b + ~I57a393cc9cc9e1abc7962aa2cc840a7c + 1;
            Ief90415b272ce5707ba28a8470132f5e = I2bcab411f9bec1541259751bcb9e0823(I037cb596cd48c5533ed22bc32518d992);
            Id4034bf7a0e92a6c92d0187e00d3df99    = Ief90415b272ce5707ba28a8470132f5e;

            I94a89577951de90edc4f73b281ad7364 = I47bf091b0fa74ad511a760bad9d2506c + ~I002869e450d79649d27441ce00bfb575 + 1;
            I386c79f4301dea9a37c9ce283e8050e4 = I2bcab411f9bec1541259751bcb9e0823(I94a89577951de90edc4f73b281ad7364);
            I44692fd63388c57268ea9035a7e4c3ef    = I386c79f4301dea9a37c9ce283e8050e4;

            Ib7493a1a384aebaa7999ff1fb867fc6b = I47bf091b0fa74ad511a760bad9d2506c + ~Id11fd3a31b70da0e64138e71840cfb83 + 1;
            I0d113fab9d7095f8d1693fec58b7c5a6 = I2bcab411f9bec1541259751bcb9e0823(Ib7493a1a384aebaa7999ff1fb867fc6b);
            I0c2892a34e5236f1366959eadfd83825    = I0d113fab9d7095f8d1693fec58b7c5a6;

            I2ceb9e423696539135c5bae5cc2d8d98 = I47bf091b0fa74ad511a760bad9d2506c + ~I0ffb8b65525af38861280645ac310e3d + 1;
            I2bbbe9e5d322d9cee76903fa813765ae = I2bcab411f9bec1541259751bcb9e0823(I2ceb9e423696539135c5bae5cc2d8d98);
            Iccef2754044e7066e191bc5e1a3805f1    = I2bbbe9e5d322d9cee76903fa813765ae;

            Ia6bbf236436b2ed22bbaae3b8849de6d = Ia4c3d0cd9957f678880de5775de76e0d + ~I8e01532a1ab9534b8de0474549d41a2e + 1;
            If5317506b6ab92c946af745a65b9e86a = I2bcab411f9bec1541259751bcb9e0823(Ia6bbf236436b2ed22bbaae3b8849de6d);
            I8ace46f1c56cfb3f4773324e0f8cae58    = If5317506b6ab92c946af745a65b9e86a;

            I33cdaee4676d546dd5507df4704ea1f8 = Ia4c3d0cd9957f678880de5775de76e0d + ~I507e9bd0265d9ca6cd21a46fa21ba084 + 1;
            Ib61ddb3ef6c7239bfc720b1761cc0221 = I2bcab411f9bec1541259751bcb9e0823(I33cdaee4676d546dd5507df4704ea1f8);
            I94ec0139bd827ef5dce2c5ee9eb9aded    = Ib61ddb3ef6c7239bfc720b1761cc0221;

            Ia44daa9ddc3e4d377267333813d4675f = Ia4c3d0cd9957f678880de5775de76e0d + ~I30fb41a57460a0b1f21065b4b97ddd42 + 1;
            I70d669976b271b2319d60114c468cae5 = I2bcab411f9bec1541259751bcb9e0823(Ia44daa9ddc3e4d377267333813d4675f);
            Ied62b116607c549ff5918d5b95e2118f    = I70d669976b271b2319d60114c468cae5;

            Ie1f8fff3f43426d6bc39e45322a532ca = If5f957fa2f055b1c2c28e8d7cfe3e9ad + ~Ifb19d75cfa0051107b5fba57bfc002b5 + 1;
            I96cb81892e2d1737d6cb25522ea2d9e4 = I2bcab411f9bec1541259751bcb9e0823(Ie1f8fff3f43426d6bc39e45322a532ca);
            I9efa5796297bc922bc5fe17f8319a515    = I96cb81892e2d1737d6cb25522ea2d9e4;

            I4ee181895efc22862b6e85802a944095 = If5f957fa2f055b1c2c28e8d7cfe3e9ad + ~I09faa07bf38acd96c4e29afd8a5167e8 + 1;
            I6c87926b040d4006c2294c516a3c46fd = I2bcab411f9bec1541259751bcb9e0823(I4ee181895efc22862b6e85802a944095);
            Ifa6908d8fda29713d7c1bbaa69b72b53    = I6c87926b040d4006c2294c516a3c46fd;

            I5c24ea83cabbb6be089ac084732cb9d6 = If5f957fa2f055b1c2c28e8d7cfe3e9ad + ~Ie8298c5c8ff538a3e37af46798f6d753 + 1;
            I549670efc854cdc29bad1d9bc03e9f5e = I2bcab411f9bec1541259751bcb9e0823(I5c24ea83cabbb6be089ac084732cb9d6);
            Ieb46857229186ce0391cddb2d30f434e    = I549670efc854cdc29bad1d9bc03e9f5e;

            Ifee2342449a3b3d0036ce2ecbc9ae189 = I3608378a5da8c66bef58528d56192530 + ~I79280400a4c9bed015106e5d006de757 + 1;
            If54c0c169048bb3e8a1423a58aed0e70 = I2bcab411f9bec1541259751bcb9e0823(Ifee2342449a3b3d0036ce2ecbc9ae189);
            I67fa03f808026b38ca5b4e71e21588bf    = If54c0c169048bb3e8a1423a58aed0e70;

            I70a9a9b8f25066612a50e411ad68e6c4 = I3608378a5da8c66bef58528d56192530 + ~I1b01cadaac7d3d15007f0afe5c0ab0f2 + 1;
            I5c956f39031611db595fbc34e6edad65 = I2bcab411f9bec1541259751bcb9e0823(I70a9a9b8f25066612a50e411ad68e6c4);
            I70938dfe09b0da9d87dafed6af3fa05c    = I5c956f39031611db595fbc34e6edad65;

            I1870059af857c79d444bef948bb536ef = I3608378a5da8c66bef58528d56192530 + ~Ie7dc322fee8ca0b6b9659e5183e0d6d6 + 1;
            I86851725f5d424c4636f9f41e5a7c7e9 = I2bcab411f9bec1541259751bcb9e0823(I1870059af857c79d444bef948bb536ef);
            Iff30a4e14b6282e9ef92e7f58230b516    = I86851725f5d424c4636f9f41e5a7c7e9;

            Iafe61ab12e232a1090123a0f16eefaca = Ie6dead855e00ea0a8e6a9b7503aaebb8 + ~I6cb09ac924c3b3b44443263e08c3315c + 1;
            Ibec300322cef05615c818b163f8a1fef = I2bcab411f9bec1541259751bcb9e0823(Iafe61ab12e232a1090123a0f16eefaca);
            I43e0faf8070869ab0528a7a4a5cdc103    = Ibec300322cef05615c818b163f8a1fef;

            I10ca809fe9a04eaf5d7784ba69314178 = Ie6dead855e00ea0a8e6a9b7503aaebb8 + ~I8741c5cc763512d16cb1186fa3323f45 + 1;
            I09cc443ecf3811a8a672c4aec1f7d6d4 = I2bcab411f9bec1541259751bcb9e0823(I10ca809fe9a04eaf5d7784ba69314178);
            Ib2f0333fac7701ae4a5589d54005b8f3    = I09cc443ecf3811a8a672c4aec1f7d6d4;

            I7a1bd0a115b3a1f85cb9c54840f5bf9b = Ie6dead855e00ea0a8e6a9b7503aaebb8 + ~I22c15857572603cc24d8a87cb47c33b0 + 1;
            Iaaf5b9288b4eb557d56908bf072cc642 = I2bcab411f9bec1541259751bcb9e0823(I7a1bd0a115b3a1f85cb9c54840f5bf9b);
            Ie4e1491da700923e81b2c1a246e528b1    = Iaaf5b9288b4eb557d56908bf072cc642;

            I986a564393d944d7d202414431c6d165 = Ie6dead855e00ea0a8e6a9b7503aaebb8 + ~I91bbec0523f77fc52a88ebcc49267e9c + 1;
            Ib224ff2bea17f6e694b10bc7cfdb898d = I2bcab411f9bec1541259751bcb9e0823(I986a564393d944d7d202414431c6d165);
            Ie8602467de2ece2013878a6b8d3129a1    = Ib224ff2bea17f6e694b10bc7cfdb898d;

            I464042aaa60a41c7e1faf3d16eeb121d = I3bae5e6862e003a8b9a476f72cc6858b + ~Iba4972a3b71a3101ab23190ed905dc17 + 1;
            Ide7d6472bf33f8dcf5c6397c7d7fb733 = I2bcab411f9bec1541259751bcb9e0823(I464042aaa60a41c7e1faf3d16eeb121d);
            I85c93c62f79b1703cb6928f96737cf27    = Ide7d6472bf33f8dcf5c6397c7d7fb733;

            I34b9a0bf2b6b562fb36291022ddf5179 = I3bae5e6862e003a8b9a476f72cc6858b + ~Ib38a46dc131d635b81fb7c196110fc4b + 1;
            Ie6193636ea1cba8b71e1d0d5f2e3c1b2 = I2bcab411f9bec1541259751bcb9e0823(I34b9a0bf2b6b562fb36291022ddf5179);
            I3dc816ee6c2a818b32f6d4e1228704bf    = Ie6193636ea1cba8b71e1d0d5f2e3c1b2;

            I17dd8612b5c7f9dcc90f17e584aab2d3 = I3bae5e6862e003a8b9a476f72cc6858b + ~Ibc03a9b6115d0941ce9233df7ef2fa57 + 1;
            Id631b0a4de889a3c3eff4df79367d3d4 = I2bcab411f9bec1541259751bcb9e0823(I17dd8612b5c7f9dcc90f17e584aab2d3);
            Id34d83701e815c01359bc5cd1b9c993c    = Id631b0a4de889a3c3eff4df79367d3d4;

            Id77cf7c05844d83e808a694971145261 = I3bae5e6862e003a8b9a476f72cc6858b + ~I38ae79956762380fadc94f8126dc1c90 + 1;
            I93d80b8bfb77e7af4d9ac734f26c4e62 = I2bcab411f9bec1541259751bcb9e0823(Id77cf7c05844d83e808a694971145261);
            I0a20e3e26261ba558d681346649cf0b3    = I93d80b8bfb77e7af4d9ac734f26c4e62;

            I276c1155d766437253f12b25066b84e4 = I4431adecba8be9e5f21bc6b3e1f8cb10 + ~I4bd98e902e805426fdd4606fcb5a5214 + 1;
            I7fba5fee37c5912e7f635feb8c111b3a = I2bcab411f9bec1541259751bcb9e0823(I276c1155d766437253f12b25066b84e4);
            I331c6e8dbe2ea1e2232f82766926d0e6    = I7fba5fee37c5912e7f635feb8c111b3a;

            Id75b386d8076893cb73baca69c3eff59 = I4431adecba8be9e5f21bc6b3e1f8cb10 + ~I6b5720d71a0b4cd10ea34affa6631a25 + 1;
            I22c14ad43399d8a1aee258826a71f50e = I2bcab411f9bec1541259751bcb9e0823(Id75b386d8076893cb73baca69c3eff59);
            Ie27046fd2751357e4a81dc62086f00be    = I22c14ad43399d8a1aee258826a71f50e;

            If62ddbe87274965cfd83189c6666401e = I4431adecba8be9e5f21bc6b3e1f8cb10 + ~Id92d779518ae724b5fef5221372f8f26 + 1;
            I3bdc4806c5c09de9a7de8d3601c57bfe = I2bcab411f9bec1541259751bcb9e0823(If62ddbe87274965cfd83189c6666401e);
            I0897ceba8201bc14a49ab30318183875    = I3bdc4806c5c09de9a7de8d3601c57bfe;

            I4f73a07452638a610b31e3ee52cb5639 = I4431adecba8be9e5f21bc6b3e1f8cb10 + ~Id55a1ab9d158ea509e5f57286a3d1b67 + 1;
            Id451569510e0d1bbba9002c2b27bb3d4 = I2bcab411f9bec1541259751bcb9e0823(I4f73a07452638a610b31e3ee52cb5639);
            Ie7b15aa8ce2492bfb433894efeb967f3    = Id451569510e0d1bbba9002c2b27bb3d4;

            I2a4faf3344d9bf4ee71da0be8994788a = I21c7a2885126d532d00484376588a469 + ~I43f52bcba1bd2e8ee5fac03320e4f19f + 1;
            I16753a377bced0688797a464157d847b = I2bcab411f9bec1541259751bcb9e0823(I2a4faf3344d9bf4ee71da0be8994788a);
            I255add08e982f701508a98db221e617d    = I16753a377bced0688797a464157d847b;

            I7d7ad0cbb962a47e229fe9d8406e6fe1 = I21c7a2885126d532d00484376588a469 + ~I391a2f354262558ff17d7d80b8c39e8c + 1;
            I76fd17f22401b66bfc0a6239a0518157 = I2bcab411f9bec1541259751bcb9e0823(I7d7ad0cbb962a47e229fe9d8406e6fe1);
            If7ca4919fa1449f38777f742ee1fb875    = I76fd17f22401b66bfc0a6239a0518157;

            I82988dc2dc83ac61380d2a5cb6551768 = I21c7a2885126d532d00484376588a469 + ~I351dc309e916f282cc1e19303eee4112 + 1;
            Ie56f8b245ab7833b6939cfea43a99874 = I2bcab411f9bec1541259751bcb9e0823(I82988dc2dc83ac61380d2a5cb6551768);
            I24cafcb5b9825321c54e84827a662fdc    = Ie56f8b245ab7833b6939cfea43a99874;

            I058c3a9848fd30010e4742d8682081ac = I21c7a2885126d532d00484376588a469 + ~Ice615e7e18356ae4c3f615dd997be943 + 1;
            I668f8103700f044c7764f2281a5b457e = I2bcab411f9bec1541259751bcb9e0823(I058c3a9848fd30010e4742d8682081ac);
            I3ede71cb7cb39774aedb9889240a2462    = I668f8103700f044c7764f2281a5b457e;

            I368121c2534820a7147858c06e58b3fc = I2c4d7339ff2fe68d060dd8d961dcab8c + ~I9306d9ef7934ffe5902306b9783c351e + 1;
            Ib75c0ca4f8b59afc2fdd7793bff7ad16 = I2bcab411f9bec1541259751bcb9e0823(I368121c2534820a7147858c06e58b3fc);
            I24da9598a6840d3ba7b12fe4f638219b    = Ib75c0ca4f8b59afc2fdd7793bff7ad16;

            I03d4541eeb1440aa72ee490c49977e32 = I2c4d7339ff2fe68d060dd8d961dcab8c + ~I70dc03a46e1ac0da826388abd3bdc503 + 1;
            I3d39fa04d24aa69d19a2db8da00eb0d3 = I2bcab411f9bec1541259751bcb9e0823(I03d4541eeb1440aa72ee490c49977e32);
            I0358ca8833007cec4ce5047db32ab7a3    = I3d39fa04d24aa69d19a2db8da00eb0d3;

            I75fdf5a355949a87b768b1e67db674e4 = I2c4d7339ff2fe68d060dd8d961dcab8c + ~I72b4ef48363856af7faacc85eafbaf2f + 1;
            I284b4ccbcb23293efe64fa45b2e0ad98 = I2bcab411f9bec1541259751bcb9e0823(I75fdf5a355949a87b768b1e67db674e4);
            I85b5354463c1c15f91ed67292da912c1    = I284b4ccbcb23293efe64fa45b2e0ad98;

            I088f4a0af0239602d422324549cb9799 = I2c4d7339ff2fe68d060dd8d961dcab8c + ~I57b40c72004f2c3072cbdefbeef72b7c + 1;
            I689ac029a268fe244a8793367c900602 = I2bcab411f9bec1541259751bcb9e0823(I088f4a0af0239602d422324549cb9799);
            Ie93731739ace44811198d0fd95b04a6a    = I689ac029a268fe244a8793367c900602;

            I787fe66b38237caf805ec14970d154c7 = Iee518b15b067eec58cccfa37f7432ea5 + ~I2882ae2eb6d79a5b96d1ed937dcfd8bf + 1;
            If53dace3e8a7be2524d711de84855015 = I2bcab411f9bec1541259751bcb9e0823(I787fe66b38237caf805ec14970d154c7);
            I464926faf4e005ad491b0bf93a365e07    = If53dace3e8a7be2524d711de84855015;

            Icef176cff3ae503dbbe2af9ecfc4c859 = Iee518b15b067eec58cccfa37f7432ea5 + ~I0dbf900b4f430b4c1106aa86b640bb37 + 1;
            Ie3fe635b63e13732c17ae2076b807b4d = I2bcab411f9bec1541259751bcb9e0823(Icef176cff3ae503dbbe2af9ecfc4c859);
            Icdaaccfead6f2d5ac2ce19caf1104d57    = Ie3fe635b63e13732c17ae2076b807b4d;

            Ie0a66e4871bfe94f6716279ecc9ef21c = Iee518b15b067eec58cccfa37f7432ea5 + ~I9dfdffbfdb83572cc3205f674e5db753 + 1;
            I1e196a61113d4db7b51f3d6b18c33da3 = I2bcab411f9bec1541259751bcb9e0823(Ie0a66e4871bfe94f6716279ecc9ef21c);
            I916d6f9429f2b0cc1bd6fb900484cde5    = I1e196a61113d4db7b51f3d6b18c33da3;

            I474adf7a975b405c288058139a08be38 = Iee518b15b067eec58cccfa37f7432ea5 + ~Ie38351e19bdc4f2ce9caf75fc3937dd4 + 1;
            Ic80e494400a5d7dcfdbf96424391e596 = I2bcab411f9bec1541259751bcb9e0823(I474adf7a975b405c288058139a08be38);
            I0142f9b3d361a0d88522f1c5f54aca84    = Ic80e494400a5d7dcfdbf96424391e596;

            Iebeadb39658f41dcf8719ed413e46144 = I42145be9c2a80288ba4a2edd91f661a3 + ~Ia8abcb8cf8d9ecc17c27ff015aa0b71f + 1;
            I69d20a7aaf2c66ed9b41fdeff0d5c6ec = I2bcab411f9bec1541259751bcb9e0823(Iebeadb39658f41dcf8719ed413e46144);
            Ie6871983b4f81b5321519647e628bd0e    = I69d20a7aaf2c66ed9b41fdeff0d5c6ec;

            Ie018b0d9f05a86207ae09ca2efac54e2 = I42145be9c2a80288ba4a2edd91f661a3 + ~I5bbbc4eedb7c61516769f429a8498ea7 + 1;
            I19b667bdb053ebd555aaa540d3a76f95 = I2bcab411f9bec1541259751bcb9e0823(Ie018b0d9f05a86207ae09ca2efac54e2);
            I17d7be125df22153fc1ed051d4e0770a    = I19b667bdb053ebd555aaa540d3a76f95;

            I51ee69807609fca0f332c8bc31afd632 = I42145be9c2a80288ba4a2edd91f661a3 + ~If49068db99aa9d09302eda27ab51fcb7 + 1;
            Ifc3d9cc420aa1274fed24b38c4d9fd8a = I2bcab411f9bec1541259751bcb9e0823(I51ee69807609fca0f332c8bc31afd632);
            I50b13959e06243e54fad2088eaf65aa7    = Ifc3d9cc420aa1274fed24b38c4d9fd8a;

            Iee1cb471704b2a8718a68ef93fd2e356 = I42145be9c2a80288ba4a2edd91f661a3 + ~Ibba6269b560db9d4913e1e515ed8270d + 1;
            Ie8a6ed15370edd38bfc92290bf7bb55a = I2bcab411f9bec1541259751bcb9e0823(Iee1cb471704b2a8718a68ef93fd2e356);
            I7a423d609b492f73d5a322849b4b1cce    = Ie8a6ed15370edd38bfc92290bf7bb55a;

            I1731c0e3be86eec142c3732ee836e4d5 = I9dc297ad41fafcda77f5347f331cfc25 + ~Iec844d10736440b96f9d6c651e604efd + 1;
            Ife5a1b49d4b0342f06ef83750ab914d4 = I2bcab411f9bec1541259751bcb9e0823(I1731c0e3be86eec142c3732ee836e4d5);
            Iefec67e214d1868670a34a7297d4a1c8    = Ife5a1b49d4b0342f06ef83750ab914d4;

            Id3b8c0ca32331f94fd98c8dae72bb15d = I9dc297ad41fafcda77f5347f331cfc25 + ~I7dbd1aeba00bb8b257990b7bb294211f + 1;
            I9906c49536062867b98ed290e49bbe50 = I2bcab411f9bec1541259751bcb9e0823(Id3b8c0ca32331f94fd98c8dae72bb15d);
            Iae7da7fdc002b635ce4285d6916d8156    = I9906c49536062867b98ed290e49bbe50;

            I6a86b0a82441c6c14436a3e0af6b0fb7 = I9dc297ad41fafcda77f5347f331cfc25 + ~I0b3a936c3f7e0391111e696b2445803b + 1;
            I41be66295070bec696e91d0f9efdc233 = I2bcab411f9bec1541259751bcb9e0823(I6a86b0a82441c6c14436a3e0af6b0fb7);
            Ic561e44b2caeae84df6720f1afa3e8f6    = I41be66295070bec696e91d0f9efdc233;

            I8c92ff598084da7a50f7c68da96620b3 = I9dc297ad41fafcda77f5347f331cfc25 + ~Ie392719059587a201c0148138ba2a2d4 + 1;
            I4838b956d8a597e78bef9a0fce82542e = I2bcab411f9bec1541259751bcb9e0823(I8c92ff598084da7a50f7c68da96620b3);
            I5be062f5b52e104ca67e615ce75a7c80    = I4838b956d8a597e78bef9a0fce82542e;

            I8bd1862e7bc2e83e9863389d532e6623 = I846700c79f30ca954cc2933fc94d355b + ~I02e672436ade3ee620c72c0d9ceee664 + 1;
            Ia06cb40e9a3341f34625c5804e02c07f = I2bcab411f9bec1541259751bcb9e0823(I8bd1862e7bc2e83e9863389d532e6623);
            Iecdde23e34c34ee0055be41f44959a19    = Ia06cb40e9a3341f34625c5804e02c07f;

            I8053269f8bd78a931878c8350693e1d6 = I846700c79f30ca954cc2933fc94d355b + ~Ie4d20df6b1e7a42f0df9a3cc26b12ac1 + 1;
            I4eaad70758412eab097822b2feda7a57 = I2bcab411f9bec1541259751bcb9e0823(I8053269f8bd78a931878c8350693e1d6);
            Ibe09be9cad0e56d5403868d072d7d628    = I4eaad70758412eab097822b2feda7a57;

            I2ff66cdd7314276232715ef2361ad184 = I846700c79f30ca954cc2933fc94d355b + ~Ie04e44d8e0756cdf34cf9ad53da76e47 + 1;
            If89e1da3daa6fd3090781723173b140b = I2bcab411f9bec1541259751bcb9e0823(I2ff66cdd7314276232715ef2361ad184);
            I464e1f3c13acaf466afb354a9b35ba0a    = If89e1da3daa6fd3090781723173b140b;

            Icf541c76bfaf37fe6111de037d205f15 = I846700c79f30ca954cc2933fc94d355b + ~I4852d6bacfd82fef6fab4502d61e9a37 + 1;
            I9ac67c519fd5a55d0ffb727389781492 = I2bcab411f9bec1541259751bcb9e0823(Icf541c76bfaf37fe6111de037d205f15);
            I160a465c22073a53510e8a4c489c3321    = I9ac67c519fd5a55d0ffb727389781492;

            I68319c8b9febef9f564832429c91b85a = I8af96a91457316e49e3f7dd5e57c82da + ~I508cea40d87bec2672f980d145c89b55 + 1;
            I73799799e5469ae887dec9b46c9c965d = I2bcab411f9bec1541259751bcb9e0823(I68319c8b9febef9f564832429c91b85a);
            I9e86d3e49827861b24f4fbeb308ad3a4    = I73799799e5469ae887dec9b46c9c965d;

            I127772614218dd7c50d3136b4f174d7a = I8af96a91457316e49e3f7dd5e57c82da + ~I80af3dcb716f3474a7257700aef89b81 + 1;
            I7ebd7c3f0617cf500deeb8c152c09af2 = I2bcab411f9bec1541259751bcb9e0823(I127772614218dd7c50d3136b4f174d7a);
            Ib96b7d796e20967e89a47e01bf424e59    = I7ebd7c3f0617cf500deeb8c152c09af2;

            Ib8d1aea4ad24c6ceb44f2cc672e1ff90 = I8af96a91457316e49e3f7dd5e57c82da + ~I6d4867d03d9187e95e27e99f7aecddec + 1;
            I2ee7d4f522ba17ca941c67079309c398 = I2bcab411f9bec1541259751bcb9e0823(Ib8d1aea4ad24c6ceb44f2cc672e1ff90);
            I565e666f6ba14b4c25e0dd402a3266e1    = I2ee7d4f522ba17ca941c67079309c398;

            I9ca26c8104bf15f48b19dc3256914544 = I8af96a91457316e49e3f7dd5e57c82da + ~I9200526d94c38e638370e9a2d7fed75c + 1;
            I62d13683ba05cfc27d9ae9a82fb04689 = I2bcab411f9bec1541259751bcb9e0823(I9ca26c8104bf15f48b19dc3256914544);
            I97e8bac5becd5128bc70f3bb48f73e6c    = I62d13683ba05cfc27d9ae9a82fb04689;

            Icc76d9ffc3f3d7b410205eeb8232a33b = I7d1c247500d7d32e406b2a5f7e2b745b + ~I844b9a89ffb7a5e48979fdea546e244a + 1;
            Ic06032eaed49f01d3d5513b2d145eaaf = I2bcab411f9bec1541259751bcb9e0823(Icc76d9ffc3f3d7b410205eeb8232a33b);
            Iced39475c6e5e3d8f36d2a5c5a80f146    = Ic06032eaed49f01d3d5513b2d145eaaf;

            I7fc4551d8a0445f79b87b4ba5f2ffeaa = I7d1c247500d7d32e406b2a5f7e2b745b + ~I9d05dc0e39e85c23b62f343a8de12e64 + 1;
            Idba6350812d3c90bee79636db48257e2 = I2bcab411f9bec1541259751bcb9e0823(I7fc4551d8a0445f79b87b4ba5f2ffeaa);
            Idcbd423c2b963c1f693dea2ddf428195    = Idba6350812d3c90bee79636db48257e2;

            I6b3c66c4e3fa0ef0cf0b52eaa4dac7a8 = I7d1c247500d7d32e406b2a5f7e2b745b + ~Ie96877deef8b1676138f814c4a720800 + 1;
            I6e7ed391604c7e0ff7cca99d5aeddc9f = I2bcab411f9bec1541259751bcb9e0823(I6b3c66c4e3fa0ef0cf0b52eaa4dac7a8);
            If1640e294bdcc51ee12fca5b3a33be6d    = I6e7ed391604c7e0ff7cca99d5aeddc9f;

            Ie34c07af9f6adb9e4b636dce3d0682c0 = I7d1c247500d7d32e406b2a5f7e2b745b + ~I15b8aa7d973edcf3b2365040f5570d82 + 1;
            Ib78d45cc282f110ed3ddaeb706a0fc12 = I2bcab411f9bec1541259751bcb9e0823(Ie34c07af9f6adb9e4b636dce3d0682c0);
            I4754c6c355e632d2ed1336b5a88c3b46    = Ib78d45cc282f110ed3ddaeb706a0fc12;

            Ib869a349250a765d2f8660e0dbdcf312 = I66d85c030a8864505298919046056305 + ~Ibddcc2e26fba20dfe2a2d399be2bc45b + 1;
            I0f5d081f9846ad888eac13d4916f5b8c = I2bcab411f9bec1541259751bcb9e0823(Ib869a349250a765d2f8660e0dbdcf312);
            I1634d703ad5d6e58a97b13ef957bdbec    = I0f5d081f9846ad888eac13d4916f5b8c;

            I1a4fb631fdc7b5454c266589962ff5f0 = I66d85c030a8864505298919046056305 + ~Ic6e3847f035738243f4c5f71f296da57 + 1;
            I607bdd63c3ee70e2721de3f994d2923e = I2bcab411f9bec1541259751bcb9e0823(I1a4fb631fdc7b5454c266589962ff5f0);
            I804e1e6a01edeb780b0159ecae707b71    = I607bdd63c3ee70e2721de3f994d2923e;

            I9de4e0e86e9edcf948d9eddf0401b94a = I66d85c030a8864505298919046056305 + ~Ie9c5e7c98281cd1deb6acc51590c9d9a + 1;
            I5453775d628c6c01c088278b6e090ddf = I2bcab411f9bec1541259751bcb9e0823(I9de4e0e86e9edcf948d9eddf0401b94a);
            Iea3c0f3c3c3017fe87a3b01647189fe0    = I5453775d628c6c01c088278b6e090ddf;

            Iee7b4838986c962969c00a0bbe53ce0b = I66d85c030a8864505298919046056305 + ~Ic3f8e77259ee3eb5be80e11b607818bd + 1;
            Iff51257cd95c2f3a38c64ae872317410 = I2bcab411f9bec1541259751bcb9e0823(Iee7b4838986c962969c00a0bbe53ce0b);
            I756b7d7e6bd3e71afa472e7e4727264a    = Iff51257cd95c2f3a38c64ae872317410;

            Id81b11a8ca1dd8989e36cef637ae6aab = I4841257ae596d9d3e4eb1e6f886956b0 + ~Ia5e26c2417aba1005971749f4ab2f367 + 1;
            Ie5faf4f522c8d24bc2d3725be57453e3 = I2bcab411f9bec1541259751bcb9e0823(Id81b11a8ca1dd8989e36cef637ae6aab);
            Ifbeae0a2acf80eda6ffd050d3bb07eb3    = Ie5faf4f522c8d24bc2d3725be57453e3;

            Ibe96deab015b799fe7f69bae8432952c = I4841257ae596d9d3e4eb1e6f886956b0 + ~If6b40a030cb120fe017bf9d39e1a35d1 + 1;
            I7952b4b62af35c930dcffe35b1629100 = I2bcab411f9bec1541259751bcb9e0823(Ibe96deab015b799fe7f69bae8432952c);
            I990ab4dcb70ee860c2c40f306ef314d3    = I7952b4b62af35c930dcffe35b1629100;

            I986b52155cc1470299321a4933241ed7 = I4841257ae596d9d3e4eb1e6f886956b0 + ~Ifdcd91f925b63e0817798aa6e9200e50 + 1;
            I47337a0b371f749c3f7f5118362c2301 = I2bcab411f9bec1541259751bcb9e0823(I986b52155cc1470299321a4933241ed7);
            Ib131087ea9ccc4bd161c3f9ac2c72303    = I47337a0b371f749c3f7f5118362c2301;

            I04be63a04f3942ce749cc9bd7540e055 = I4841257ae596d9d3e4eb1e6f886956b0 + ~Iabf228f57ac154c417389f6711af1950 + 1;
            I21ea597751b3243936aea7c07cc90f70 = I2bcab411f9bec1541259751bcb9e0823(I04be63a04f3942ce749cc9bd7540e055);
            I9a967ac9d11583faaa783984229aeb2c    = I21ea597751b3243936aea7c07cc90f70;

            Ia7adea5b0ec86e9fcd427a5468d72b64 = Icd6f7ec117f9ab4eda8c5eba41386ffa + ~I9fdfe73e77c384d33196c0f2d2a2fde2 + 1;
            Ibdce05e98adef0314000dba3c482ace6 = I2bcab411f9bec1541259751bcb9e0823(Ia7adea5b0ec86e9fcd427a5468d72b64);
            Ib9921dfcf121e5f4ac4d8be83a868210    = Ibdce05e98adef0314000dba3c482ace6;

            Ie8990d8abd23f8f9f79d7fe38c57fa8c = Icd6f7ec117f9ab4eda8c5eba41386ffa + ~I30b5c7aadb5312ce96e833704bb3a320 + 1;
            If0dbc84f59311eeabfb57b5fd0c3b632 = I2bcab411f9bec1541259751bcb9e0823(Ie8990d8abd23f8f9f79d7fe38c57fa8c);
            If22d8fd45caed08b2c7cee8b7349700f    = If0dbc84f59311eeabfb57b5fd0c3b632;

            I9d2f90ddddbdbb525d5f070f32546b64 = Icd6f7ec117f9ab4eda8c5eba41386ffa + ~Ia18bdb8d2f02b50281f0acd4a45ac973 + 1;
            I74f2e7798a8383b78a5e7b816c2370af = I2bcab411f9bec1541259751bcb9e0823(I9d2f90ddddbdbb525d5f070f32546b64);
            Iabf029e67c7f827faf17b6518cd1bfa3    = I74f2e7798a8383b78a5e7b816c2370af;

            I905256d73bdb63bf860e15687350795f = Icd6f7ec117f9ab4eda8c5eba41386ffa + ~If37de611ce4fa330c4fc9dcb87d4d95c + 1;
            I58ee302a3a1faa2b44d9052bffbc2a03 = I2bcab411f9bec1541259751bcb9e0823(I905256d73bdb63bf860e15687350795f);
            Iaeab83001c6285630e3404ae67227f46    = I58ee302a3a1faa2b44d9052bffbc2a03;

            I9adcfc18e4471209edbe9a379e996067 = Ibc0498839d1d9b6dc853b8e5d7a88fa3 + ~Id924dafd31fd0af0b28c7e6b7e95ec37 + 1;
            I979a71fc0942bf62c06405bb63a717c5 = I2bcab411f9bec1541259751bcb9e0823(I9adcfc18e4471209edbe9a379e996067);
            I53ac6d02d2bfc9aca9469148753070a7    = I979a71fc0942bf62c06405bb63a717c5;

            I3d7d048348bf833f744a9f73889b7802 = Ibc0498839d1d9b6dc853b8e5d7a88fa3 + ~I926c049036f53f0a0a6ad369de116c57 + 1;
            I30be0ac758b5a0fbacb1c51a36ca8a73 = I2bcab411f9bec1541259751bcb9e0823(I3d7d048348bf833f744a9f73889b7802);
            I61992979f60b26d313efd1dc23bb54ab    = I30be0ac758b5a0fbacb1c51a36ca8a73;

            Id619e8d4040014d0e415ff71c5e0591f = Ibc0498839d1d9b6dc853b8e5d7a88fa3 + ~Id0762ac7710c93249bc11c6ce4ae51a0 + 1;
            I9c50e0a8a01aaed98ae54530d5c76ba1 = I2bcab411f9bec1541259751bcb9e0823(Id619e8d4040014d0e415ff71c5e0591f);
            I8b46b3f0835310114208963de7ac8e97    = I9c50e0a8a01aaed98ae54530d5c76ba1;

            Iaf3de2ef283e03dd72002026e1299224 = Ibc0498839d1d9b6dc853b8e5d7a88fa3 + ~If3c44eb85217da3b6bddb5aed97a9bb7 + 1;
            I0daac80ebeec26e428328344a398ce57 = I2bcab411f9bec1541259751bcb9e0823(Iaf3de2ef283e03dd72002026e1299224);
            Icda26ba6f5c7f77a80776b2c1bbc975d    = I0daac80ebeec26e428328344a398ce57;

            I64551529c0028ec145407be7f5dfef71 = I142ebca7f155e287e38ddf45423ab0fd + ~I33703f538ec70268e6c00ad6eef6c4e0 + 1;
            I6739f13ea431943bb5bacb4a05140063 = I2bcab411f9bec1541259751bcb9e0823(I64551529c0028ec145407be7f5dfef71);
            I0863565b3ae88137a2384750436f9e19    = I6739f13ea431943bb5bacb4a05140063;

            I5ebe580a943b65fb16ea722ba101fd05 = I142ebca7f155e287e38ddf45423ab0fd + ~Ifc7eec6765af08463751db128f8818b3 + 1;
            Ifa0e560fe6445b006ab74096a807b90f = I2bcab411f9bec1541259751bcb9e0823(I5ebe580a943b65fb16ea722ba101fd05);
            Id646110f8d09cd47dc7695e05f73efc6    = Ifa0e560fe6445b006ab74096a807b90f;

            I0921901599c43b27e701758026dd3ee1 = I142ebca7f155e287e38ddf45423ab0fd + ~I9de5e90485b3f22e9003dc8a7b22a79b + 1;
            I9595c0fd77d6a0610eb859dcd2b67d1d = I2bcab411f9bec1541259751bcb9e0823(I0921901599c43b27e701758026dd3ee1);
            I5999eef2304e579a3d47e4f15ba336e1    = I9595c0fd77d6a0610eb859dcd2b67d1d;

            I6033532f27c26b2d42bb3ea128f80dfa = I142ebca7f155e287e38ddf45423ab0fd + ~I8c36318c45dabe6bf540381373f09fe5 + 1;
            I6f3e685e70fa700b52bec62d0aed942c = I2bcab411f9bec1541259751bcb9e0823(I6033532f27c26b2d42bb3ea128f80dfa);
            Idd302bdc6ff8368a6b73d53bbc8f8425    = I6f3e685e70fa700b52bec62d0aed942c;
end

   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
              Ifc045af19c3f10d92d2b0dfb4fbbde38 <= {(SUM_LEN){1'b0}};
       end else begin
           if (I86a86d41a29fd0d7596d668e79aca825) begin
              if (Ib325dab091dfc3a1a269adb3ea9c75cd <= HamDist_sum_mm) begin
                  Ifc045af19c3f10d92d2b0dfb4fbbde38 <= Ifc045af19c3f10d92d2b0dfb4fbbde38 + 1;
              end
           end
           else if (start_dec) begin
                  Ifc045af19c3f10d92d2b0dfb4fbbde38 <= {(SUM_LEN){1'b0}};
           end
       end
   end

   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
                 Ieb085b219090cde5da2190093ce43730 <= 'h0;
       end else begin
          if (Ibd047e2643dc68affb5b4f25b82ded31) begin
             if (HamDist_loop == 0)
                 Ieb085b219090cde5da2190093ce43730 <= HamDist_sum_mm;
             else
                 Ieb085b219090cde5da2190093ce43730 <= Ib79e305e6f44a4a6ebef1db5c70246ea;
          end
       end
   end

   always_comb Ib79e305e6f44a4a6ebef1db5c70246ea = ((Ieb085b219090cde5da2190093ce43730 * HamDist_iir1 + HamDist_sum_mm *HamDist_iir2 + HamDist_iir3));



   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
                 Ib325dab091dfc3a1a269adb3ea9c75cd <= {(SUM_LEN){1'b0}};
       end else begin
          if (Ibd047e2643dc68affb5b4f25b82ded31) begin
             if (HamDist_loop == 0)
                 Ib325dab091dfc3a1a269adb3ea9c75cd <= {(SUM_LEN){1'b0}};
             else
                 Ib325dab091dfc3a1a269adb3ea9c75cd <= HamDist_sum_mm;
          end
       end
   end





   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
          converged_loops_ended <= 1'b0;
          converged_pass_fail <= 1'b0;
       end else begin
          if (start_dec) begin
               converged_loops_ended <= 1'b0;
               converged_pass_fail <= 1'b0;
          end else begin
               if (I65e382d77592c7d1af308d171b27ff3c) begin
                       if (
                         (HamDist_sum_mm*100 > Ieb085b219090cde5da2190093ce43730 * HamDist_loop_percentage) ||
                         (Ifc045af19c3f10d92d2b0dfb4fbbde38 > HamDist_loop_max)
                         ) begin
                         converged_loops_ended <= 1'b1;
                         converged_pass_fail <= 1'b0;
                       end else if (HamDist_sum_mm == 0) begin
                         converged_loops_ended <= 1'b1;
                         converged_pass_fail <= 1'b1;
                       end

               end  //I65e382d77592c7d1af308d171b27ff3c
               else begin // else I8bf8854bebe108183caeb845c7676ae4 I65e382d77592c7d1af308d171b27ff3c
                    //wait for I8fc42c6ddf9966db3b09e84365034357 start_dec to I01bc6f8efa4202821e95f4fdf6298b30 I0d149b90e7394297301c90191ae775f0 I3262d48df5d75e3452f0f16b313b7808
                    //converged_loops_ended <= 1'b0;
                    //converged_pass_fail <= 1'b0;
               end


          end  //start_dec
       end  //rstn
   end

//tmp_bit valid Ied2b5c0139cec8ad2873829dc1117d50 I6d3acefe6d7dfb94a5d66dcaa1bbbb76
// I7fa3b767c460b54a2be4d49030b349c7 I9a4c07402cc2f3740fb5849a16920e13 I7243f8be75253afbadf7477867021f8b I13b5bfe96f3e2fe411c9f66f4a582adf I724a00e315992b82d662231ea0dcbe50 or I190ebdd6b6c2b422296a6ee2cce59699 I0aa6f4210bf373c95eda00232e93cd98
always_comb HamDist_cntr_inc_converged_valid = I6d3acefe6d7dfb94a5d66dcaa1bbbb76;

//I3e47b75000b0924b6c9ba5759a7cf15d I6b2ded51d81a4403d8a4bd25fa1e57ee Ied2b5c0139cec8ad2873829dc1117d50 valid ??

always_comb I86a86d41a29fd0d7596d668e79aca825 = I6d3acefe6d7dfb94a5d66dcaa1bbbb76;
always_comb hamming_code_calc_out             = I86a86d41a29fd0d7596d668e79aca825;


`ifdef ENCRYPT
`endif

endmodule

//C Ia642a85aab89544a289fb1f29eab689d: Ib6f6b4efd9391d1fa207d325ff1bbd60 I83878c91171338902e0fe0fb97a8c47a:0.100000 I7290d6b1f1458098d2f225877e609ba6:2.197225 percent_probability_int:'d4500

 //Ic07b0b4d7660314f711a68fc47c4ab38 I48d8d6f5a3efbf52837d6b788a22859a valid Ic13367945d5d4c91047b3b50234aa7ab Ic47d187067c6cf953245f128b5fde62a
//y_int:
 //462d03cd366ba17b39e149628fe20b0640ff49b27104e774ce83
//Iebc6097498b06421e2759a773c992ed3:
 //612c501115962aad76ce8207211dbe3416e483efed
//C Ia642a85aab89544a289fb1f29eab689d: Ib6f6b4efd9391d1fa207d325ff1bbd60 I83878c91171338902e0fe0fb97a8c47a:0.225962 I7290d6b1f1458098d2f225877e609ba6:1.231257 percent_probability_int:'d2522
