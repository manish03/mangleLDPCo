 reg  ['h7fff:0] [$clog2('h7000+1)-1:0] I8a0037ad2845a3fbba9da380a8b8a576 ;
