//`include "GF2_LDPC_fgallag_0x00006_assign_inc.sv"
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00000] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00000] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00001] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00001] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00002] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00003] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00002] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00004] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00005] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00003] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00006] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00007] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00004] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00008] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00009] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00005] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0000a] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0000b] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00006] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0000c] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0000d] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00007] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0000e] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0000f] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00008] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00010] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00011] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00009] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00012] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00013] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0000a] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00014] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00015] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0000b] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00016] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00017] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0000c] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00018] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00019] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0000d] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0001a] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0001b] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0000e] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0001c] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0001d] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0000f] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0001e] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0001f] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00010] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00020] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00021] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00011] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00022] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00023] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00012] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00024] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00025] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00013] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00026] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00027] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00014] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00028] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00029] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00015] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0002a] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0002b] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00016] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0002c] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0002d] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00017] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0002e] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0002f] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00018] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00030] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00031] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00019] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00032] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00033] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0001a] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00034] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00035] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0001b] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00036] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00037] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0001c] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00038] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00039] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0001d] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0003a] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0003b] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0001e] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0003c] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0003d] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0001f] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0003e] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0003f] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00020] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00040] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00041] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00021] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00042] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00043] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00022] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00044] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00045] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00023] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00046] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00047] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00024] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00048] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00049] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00025] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0004a] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0004b] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00026] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0004c] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0004d] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00027] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0004e] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0004f] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00028] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00050] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00051] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00029] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00052] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00053] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0002a] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00054] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00055] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0002b] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00056] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00057] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0002c] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00058] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00059] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0002d] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0005a] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0005b] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0002e] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0005c] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0005d] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0002f] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0005e] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0005f] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00030] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00060] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00061] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00031] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00062] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00063] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00032] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00064] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00065] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00033] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00066] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00067] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00034] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00068] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00069] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00035] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0006a] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0006b] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00036] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0006c] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0006d] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00037] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0006e] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0006f] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00038] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00070] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00071] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00039] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00072] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00073] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0003a] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00074] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00075] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0003b] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00076] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00077] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0003c] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00078] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00079] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0003d] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0007a] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0007b] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0003e] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0007c] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0007d] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0003f] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0007e] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0007f] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00040] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00080] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00081] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00041] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00082] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00083] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00042] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00084] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00085] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00043] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00086] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00087] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00044] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00088] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00089] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00045] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0008a] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0008b] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00046] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0008c] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0008d] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00047] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0008e] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0008f] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00048] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00090] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00091] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00049] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00092] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00093] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0004a] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00094] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00095] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0004b] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00096] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00097] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0004c] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00098] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00099] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0004d] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0009a] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0009b] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0004e] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0009c] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0009d] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0004f] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0009e] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0009f] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00050] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000a0] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000a1] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00051] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000a2] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000a3] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00052] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000a4] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000a5] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00053] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000a6] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000a7] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00054] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000a8] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000a9] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00055] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000aa] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000ab] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00056] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000ac] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000ad] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00057] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000ae] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000af] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00058] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000b0] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000b1] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00059] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000b2] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000b3] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0005a] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000b4] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000b5] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0005b] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000b6] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000b7] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0005c] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000b8] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000b9] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0005d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000ba] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0005e] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000bc] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000bd] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0005f] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000be] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000bf] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00060] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000c0] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00061] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000c2] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000c3] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00062] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000c4] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000c5] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00063] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000c6] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00064] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000c8] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000c9] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00065] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000ca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00066] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000cc] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00067] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000ce] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000cf] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00068] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000d0] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00069] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000d2] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000d3] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0006a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000d4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0006b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000d6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0006c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000d8] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0006d] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000da] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000db] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0006e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000dc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0006f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000de] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00070] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000e0] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00071] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000e2] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000e3] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00072] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000e4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00073] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000e6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00074] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000e8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00075] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000ea] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00076] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000ec] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000ed] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00077] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000ee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00078] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000f0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00079] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000f2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0007a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000f4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0007b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000f6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0007c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000f8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0007d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000fa] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0007e] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000fc] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000fd] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0007f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h000fe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00080] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00100] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00081] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00102] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00082] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00104] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00083] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00106] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00084] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00108] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00085] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0010a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00086] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0010c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00087] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0010e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00088] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00110] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00089] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00112] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0008a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00114] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0008b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00116] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0008c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00118] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0008d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0011a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0008e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0011c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0008f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0011e] ;
//end
//always_comb begin
              I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00090] = 
          (!fgallag_sel['h00006]) ? 
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00120] : //%
                       Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00121] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00091] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00122] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00092] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00124] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00093] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00126] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00094] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00128] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00095] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0012a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00096] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0012c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00097] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0012e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00098] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00130] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00099] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00132] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0009a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00134] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0009b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00136] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0009c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00138] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0009d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0013a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0009e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0013c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0009f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0013e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000a0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00140] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000a1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00142] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000a2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00144] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000a3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00146] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000a4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00148] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000a5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0014a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000a6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0014c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000a7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0014e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000a8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00150] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000a9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00152] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000aa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00154] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000ab] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00156] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000ac] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00158] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000ad] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0015a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000ae] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0015c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000af] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0015e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000b0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00160] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000b1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00162] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000b2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00164] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000b3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00166] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000b4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00168] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000b5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0016a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000b6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0016c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000b7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0016e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000b8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00170] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000b9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00172] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000ba] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00174] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000bb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00176] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000bc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00178] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000bd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0017a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000be] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0017c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000bf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0017e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000c0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00180] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000c1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00182] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000c2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00184] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000c3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00186] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000c4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00188] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000c5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0018a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000c6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0018c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000c7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0018e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000c8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00190] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000c9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00192] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000ca] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00194] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000cb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00196] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000cc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00198] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000cd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0019a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000ce] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0019c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000cf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0019e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000d0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001a0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000d1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001a2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000d2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001a4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000d3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001a6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000d4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001a8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000d5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001aa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000d6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001ac] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000d7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001ae] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000d8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001b0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000d9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001b2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000da] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001b4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000db] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001b6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000dc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001b8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000dd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001ba] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000de] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001bc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000df] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001be] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000e0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001c0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000e1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001c2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000e2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001c4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000e3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001c6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000e4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001c8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000e5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001ca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000e6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001cc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000e7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001ce] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000e8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001d0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000e9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001d2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000ea] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001d4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000eb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001d6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000ec] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001d8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000ed] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001da] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000ee] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001dc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000ef] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001de] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000f0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001e0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000f1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001e2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000f2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001e4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000f3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001e6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000f4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001e8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000f5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001ea] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000f6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001ec] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000f7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001ee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000f8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001f0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000f9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001f2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000fa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001f4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000fb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001f6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000fc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001f8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000fd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001fa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000fe] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001fc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000ff] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h001fe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00100] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00200] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00101] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00202] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00102] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00204] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00103] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00206] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00104] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00208] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00105] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0020a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00106] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0020c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00107] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0020e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00108] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00210] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00109] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00212] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0010a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00214] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0010b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00216] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0010c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00218] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0010d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0021a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0010e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0021c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0010f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0021e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00110] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00220] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00111] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00222] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00112] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00224] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00113] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00226] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00114] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00228] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00115] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0022a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00116] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0022c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00117] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0022e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00118] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00230] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00119] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00232] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0011a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00234] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0011b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00236] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0011c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00238] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0011d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0023a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0011e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0023c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0011f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0023e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00120] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00240] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00121] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00242] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00122] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00244] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00123] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00246] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00124] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00248] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00125] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0024a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00126] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0024c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00127] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0024e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00128] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00250] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00129] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00252] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0012a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00254] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0012b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00256] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0012c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00258] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0012d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0025a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0012e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0025c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0012f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0025e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00130] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00260] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00131] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00262] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00132] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00264] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00133] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00266] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00134] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00268] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00135] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0026a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00136] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0026c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00137] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0026e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00138] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00270] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00139] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00272] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0013a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00274] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0013b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00276] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0013c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00278] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0013d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0027a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0013e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0027c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0013f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0027e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00140] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00280] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00141] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00282] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00142] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00284] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00143] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00286] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00144] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00288] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00145] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0028a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00146] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0028c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00147] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0028e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00148] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00290] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00149] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00292] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0014a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00294] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0014b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00296] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0014c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00298] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0014d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0029a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0014e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0029c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0014f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0029e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00150] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002a0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00151] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002a2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00152] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002a4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00153] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002a6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00154] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002a8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00155] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002aa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00156] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002ac] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00157] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002ae] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00158] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002b0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00159] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002b2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0015a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002b4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0015b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002b6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0015c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002b8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0015d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002ba] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0015e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002bc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0015f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002be] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00160] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002c0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00161] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002c2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00162] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002c4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00163] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002c6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00164] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002c8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00165] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002ca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00166] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002cc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00167] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002ce] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00168] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002d0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00169] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002d2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0016a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002d4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0016b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002d6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0016c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002d8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0016d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002da] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0016e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002dc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0016f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002de] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00170] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002e0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00171] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002e2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00172] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002e4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00173] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002e6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00174] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002e8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00175] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002ea] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00176] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002ec] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00177] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002ee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00178] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002f0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00179] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002f2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0017a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002f4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0017b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002f6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0017c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002f8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0017d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002fa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0017e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002fc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0017f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h002fe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00180] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00300] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00181] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00302] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00182] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00304] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00183] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00306] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00184] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00308] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00185] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0030a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00186] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0030c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00187] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0030e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00188] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00310] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00189] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00312] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0018a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00314] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0018b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00316] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0018c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00318] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0018d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0031a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0018e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0031c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0018f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0031e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00190] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00320] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00191] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00322] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00192] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00324] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00193] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00326] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00194] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00328] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00195] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0032a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00196] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0032c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00197] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0032e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00198] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00330] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00199] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00332] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0019a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00334] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0019b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00336] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0019c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00338] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0019d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0033a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0019e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0033c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0019f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0033e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001a0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00340] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001a1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00342] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001a2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00344] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001a3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00346] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001a4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00348] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001a5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0034a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001a6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0034c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001a7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0034e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001a8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00350] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001a9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00352] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001aa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00354] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001ab] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00356] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001ac] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00358] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001ad] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0035a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001ae] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0035c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001af] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0035e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001b0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00360] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001b1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00362] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001b2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00364] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001b3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00366] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001b4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00368] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001b5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0036a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001b6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0036c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001b7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0036e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001b8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00370] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001b9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00372] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001ba] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00374] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001bb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00376] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001bc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00378] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001bd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0037a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001be] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0037c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001bf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0037e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001c0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00380] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001c1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00382] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001c2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00384] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001c3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00386] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001c4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00388] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001c5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0038a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001c6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0038c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001c7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0038e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001c8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00390] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001c9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00392] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001ca] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00394] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001cb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00396] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001cc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00398] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001cd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0039a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001ce] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0039c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001cf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0039e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001d0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003a0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001d1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003a2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001d2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003a4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001d3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003a6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001d4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003a8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001d5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003aa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001d6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003ac] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001d7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003ae] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001d8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003b0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001d9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003b2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001da] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003b4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001db] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003b6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001dc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003b8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001dd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003ba] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001de] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003bc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001df] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003be] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001e0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003c0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001e1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003c2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001e2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003c4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001e3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003c6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001e4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003c8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001e5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003ca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001e6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003cc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001e7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003ce] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001e8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003d0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001e9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003d2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001ea] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003d4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001eb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003d6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001ec] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003d8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001ed] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003da] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001ee] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003dc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001ef] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003de] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001f0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003e0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001f1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003e2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001f2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003e4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001f3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003e6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001f4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003e8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001f5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003ea] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001f6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003ec] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001f7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003ee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001f8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003f0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001f9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003f2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001fa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003f4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001fb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003f6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001fc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003f8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001fd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003fa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001fe] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003fc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001ff] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h003fe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00200] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00400] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00201] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00402] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00202] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00404] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00203] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00406] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00204] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00408] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00205] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0040a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00206] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0040c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00207] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0040e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00208] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00410] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00209] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00412] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0020a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00414] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0020b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00416] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0020c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00418] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0020d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0041a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0020e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0041c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0020f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0041e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00210] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00420] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00211] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00422] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00212] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00424] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00213] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00426] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00214] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00428] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00215] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0042a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00216] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0042c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00217] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0042e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00218] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00430] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00219] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00432] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0021a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00434] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0021b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00436] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0021c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00438] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0021d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0043a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0021e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0043c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0021f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0043e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00220] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00440] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00221] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00442] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00222] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00444] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00223] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00446] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00224] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00448] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00225] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0044a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00226] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0044c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00227] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0044e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00228] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00450] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00229] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00452] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0022a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00454] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0022b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00456] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0022c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00458] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0022d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0045a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0022e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0045c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0022f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0045e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00230] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00460] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00231] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00462] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00232] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00464] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00233] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00466] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00234] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00468] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00235] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0046a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00236] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0046c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00237] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0046e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00238] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00470] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00239] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00472] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0023a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00474] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0023b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00476] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0023c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00478] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0023d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0047a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0023e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0047c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0023f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0047e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00240] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00480] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00241] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00482] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00242] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00484] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00243] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00486] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00244] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00488] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00245] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0048a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00246] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0048c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00247] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0048e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00248] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00490] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00249] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00492] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0024a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00494] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0024b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00496] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0024c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00498] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0024d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0049a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0024e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0049c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0024f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0049e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00250] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004a0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00251] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004a2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00252] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004a4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00253] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004a6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00254] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004a8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00255] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004aa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00256] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004ac] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00257] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004ae] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00258] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004b0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00259] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004b2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0025a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004b4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0025b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004b6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0025c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004b8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0025d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004ba] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0025e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004bc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0025f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004be] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00260] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004c0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00261] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004c2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00262] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004c4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00263] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004c6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00264] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004c8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00265] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004ca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00266] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004cc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00267] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004ce] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00268] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004d0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00269] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004d2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0026a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004d4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0026b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004d6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0026c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004d8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0026d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004da] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0026e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004dc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0026f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004de] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00270] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004e0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00271] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004e2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00272] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004e4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00273] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004e6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00274] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004e8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00275] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004ea] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00276] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004ec] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00277] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004ee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00278] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004f0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00279] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004f2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0027a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004f4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0027b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004f6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0027c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004f8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0027d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004fa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0027e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004fc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0027f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h004fe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00280] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00500] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00281] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00502] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00282] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00504] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00283] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00506] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00284] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00508] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00285] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0050a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00286] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0050c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00287] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0050e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00288] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00510] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00289] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00512] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0028a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00514] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0028b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00516] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0028c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00518] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0028d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0051a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0028e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0051c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0028f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0051e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00290] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00520] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00291] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00522] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00292] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00524] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00293] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00526] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00294] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00528] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00295] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0052a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00296] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0052c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00297] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0052e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00298] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00530] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00299] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00532] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0029a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00534] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0029b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00536] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0029c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00538] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0029d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0053a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0029e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0053c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0029f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0053e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002a0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00540] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002a1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00542] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002a2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00544] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002a3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00546] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002a4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00548] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002a5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0054a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002a6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0054c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002a7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0054e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002a8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00550] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002a9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00552] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002aa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00554] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002ab] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00556] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002ac] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00558] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002ad] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0055a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002ae] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0055c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002af] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0055e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002b0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00560] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002b1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00562] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002b2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00564] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002b3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00566] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002b4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00568] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002b5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0056a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002b6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0056c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002b7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0056e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002b8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00570] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002b9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00572] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002ba] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00574] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002bb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00576] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002bc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00578] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002bd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0057a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002be] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0057c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002bf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0057e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002c0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00580] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002c1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00582] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002c2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00584] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002c3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00586] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002c4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00588] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002c5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0058a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002c6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0058c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002c7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0058e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002c8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00590] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002c9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00592] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002ca] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00594] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002cb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00596] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002cc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00598] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002cd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0059a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002ce] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0059c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002cf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0059e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002d0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005a0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002d1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005a2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002d2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005a4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002d3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005a6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002d4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005a8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002d5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005aa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002d6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005ac] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002d7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005ae] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002d8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005b0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002d9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005b2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002da] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005b4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002db] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005b6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002dc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005b8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002dd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005ba] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002de] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005bc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002df] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005be] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002e0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005c0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002e1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005c2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002e2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005c4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002e3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005c6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002e4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005c8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002e5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005ca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002e6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005cc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002e7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005ce] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002e8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005d0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002e9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005d2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002ea] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005d4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002eb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005d6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002ec] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005d8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002ed] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005da] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002ee] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005dc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002ef] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005de] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002f0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005e0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002f1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005e2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002f2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005e4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002f3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005e6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002f4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005e8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002f5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005ea] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002f6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005ec] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002f7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005ee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002f8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005f0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002f9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005f2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002fa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005f4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002fb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005f6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002fc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005f8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002fd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005fa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002fe] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005fc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002ff] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h005fe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00300] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00600] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00301] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00602] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00302] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00604] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00303] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00606] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00304] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00608] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00305] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0060a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00306] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0060c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00307] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0060e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00308] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00610] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00309] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00612] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0030a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00614] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0030b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00616] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0030c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00618] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0030d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0061a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0030e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0061c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0030f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0061e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00310] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00620] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00311] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00622] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00312] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00624] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00313] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00626] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00314] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00628] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00315] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0062a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00316] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0062c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00317] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0062e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00318] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00630] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00319] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00632] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0031a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00634] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0031b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00636] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0031c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00638] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0031d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0063a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0031e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0063c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0031f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0063e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00320] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00640] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00321] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00642] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00322] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00644] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00323] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00646] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00324] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00648] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00325] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0064a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00326] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0064c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00327] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0064e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00328] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00650] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00329] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00652] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0032a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00654] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0032b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00656] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0032c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00658] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0032d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0065a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0032e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0065c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0032f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0065e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00330] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00660] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00331] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00662] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00332] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00664] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00333] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00666] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00334] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00668] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00335] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0066a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00336] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0066c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00337] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0066e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00338] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00670] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00339] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00672] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0033a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00674] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0033b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00676] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0033c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00678] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0033d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0067a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0033e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0067c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0033f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0067e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00340] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00680] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00341] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00682] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00342] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00684] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00343] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00686] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00344] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00688] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00345] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0068a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00346] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0068c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00347] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0068e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00348] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00690] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00349] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00692] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0034a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00694] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0034b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00696] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0034c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00698] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0034d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0069a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0034e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0069c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0034f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0069e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00350] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006a0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00351] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006a2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00352] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006a4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00353] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006a6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00354] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006a8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00355] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006aa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00356] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006ac] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00357] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006ae] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00358] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006b0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00359] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006b2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0035a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006b4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0035b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006b6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0035c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006b8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0035d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006ba] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0035e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006bc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0035f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006be] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00360] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006c0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00361] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006c2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00362] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006c4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00363] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006c6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00364] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006c8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00365] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006ca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00366] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006cc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00367] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006ce] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00368] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006d0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00369] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006d2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0036a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006d4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0036b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006d6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0036c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006d8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0036d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006da] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0036e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006dc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0036f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006de] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00370] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006e0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00371] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006e2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00372] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006e4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00373] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006e6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00374] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006e8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00375] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006ea] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00376] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006ec] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00377] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006ee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00378] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006f0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00379] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006f2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0037a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006f4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0037b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006f6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0037c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006f8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0037d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006fa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0037e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006fc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0037f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h006fe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00380] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00700] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00381] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00702] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00382] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00704] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00383] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00706] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00384] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00708] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00385] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0070a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00386] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0070c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00387] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0070e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00388] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00710] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00389] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00712] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0038a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00714] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0038b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00716] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0038c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00718] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0038d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0071a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0038e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0071c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0038f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0071e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00390] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00720] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00391] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00722] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00392] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00724] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00393] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00726] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00394] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00728] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00395] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0072a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00396] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0072c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00397] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0072e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00398] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00730] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00399] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00732] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0039a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00734] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0039b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00736] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0039c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00738] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0039d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0073a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0039e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0073c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0039f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0073e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003a0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00740] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003a1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00742] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003a2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00744] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003a3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00746] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003a4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00748] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003a5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0074a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003a6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0074c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003a7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0074e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003a8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00750] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003a9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00752] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003aa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00754] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003ab] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00756] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003ac] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00758] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003ad] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0075a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003ae] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0075c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003af] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0075e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003b0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00760] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003b1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00762] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003b2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00764] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003b3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00766] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003b4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00768] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003b5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0076a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003b6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0076c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003b7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0076e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003b8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00770] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003b9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00772] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003ba] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00774] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003bb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00776] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003bc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00778] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003bd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0077a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003be] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0077c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003bf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0077e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003c0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00780] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003c1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00782] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003c2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00784] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003c3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00786] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003c4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00788] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003c5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0078a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003c6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0078c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003c7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0078e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003c8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00790] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003c9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00792] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003ca] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00794] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003cb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00796] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003cc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00798] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003cd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0079a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003ce] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0079c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003cf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0079e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003d0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007a0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003d1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007a2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003d2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007a4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003d3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007a6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003d4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007a8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003d5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007aa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003d6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007ac] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003d7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007ae] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003d8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007b0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003d9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007b2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003da] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007b4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003db] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007b6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003dc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007b8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003dd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007ba] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003de] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007bc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003df] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007be] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003e0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007c0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003e1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007c2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003e2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007c4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003e3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007c6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003e4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007c8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003e5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007ca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003e6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007cc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003e7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007ce] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003e8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007d0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003e9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007d2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003ea] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007d4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003eb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007d6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003ec] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007d8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003ed] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007da] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003ee] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007dc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003ef] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007de] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003f0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007e0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003f1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007e2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003f2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007e4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003f3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007e6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003f4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007e8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003f5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007ea] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003f6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007ec] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003f7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007ee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003f8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007f0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003f9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007f2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003fa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007f4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003fb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007f6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003fc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007f8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003fd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007fa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003fe] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007fc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003ff] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h007fe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00400] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00800] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00401] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00802] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00402] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00804] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00403] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00806] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00404] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00808] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00405] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0080a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00406] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0080c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00407] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0080e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00408] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00810] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00409] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00812] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0040a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00814] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0040b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00816] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0040c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00818] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0040d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0081a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0040e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0081c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0040f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0081e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00410] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00820] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00411] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00822] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00412] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00824] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00413] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00826] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00414] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00828] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00415] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0082a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00416] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0082c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00417] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0082e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00418] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00830] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00419] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00832] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0041a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00834] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0041b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00836] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0041c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00838] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0041d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0083a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0041e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0083c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0041f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0083e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00420] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00840] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00421] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00842] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00422] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00844] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00423] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00846] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00424] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00848] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00425] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0084a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00426] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0084c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00427] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0084e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00428] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00850] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00429] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00852] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0042a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00854] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0042b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00856] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0042c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00858] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0042d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0085a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0042e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0085c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0042f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0085e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00430] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00860] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00431] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00862] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00432] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00864] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00433] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00866] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00434] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00868] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00435] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0086a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00436] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0086c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00437] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0086e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00438] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00870] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00439] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00872] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0043a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00874] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0043b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00876] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0043c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00878] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0043d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0087a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0043e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0087c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0043f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0087e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00440] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00880] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00441] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00882] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00442] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00884] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00443] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00886] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00444] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00888] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00445] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0088a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00446] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0088c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00447] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0088e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00448] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00890] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00449] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00892] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0044a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00894] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0044b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00896] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0044c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00898] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0044d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0089a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0044e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0089c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0044f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0089e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00450] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008a0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00451] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008a2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00452] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008a4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00453] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008a6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00454] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008a8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00455] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008aa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00456] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008ac] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00457] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008ae] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00458] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008b0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00459] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008b2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0045a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008b4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0045b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008b6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0045c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008b8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0045d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008ba] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0045e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008bc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0045f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008be] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00460] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008c0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00461] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008c2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00462] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008c4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00463] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008c6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00464] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008c8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00465] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008ca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00466] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008cc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00467] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008ce] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00468] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008d0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00469] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008d2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0046a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008d4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0046b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008d6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0046c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008d8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0046d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008da] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0046e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008dc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0046f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008de] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00470] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008e0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00471] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008e2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00472] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008e4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00473] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008e6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00474] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008e8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00475] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008ea] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00476] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008ec] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00477] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008ee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00478] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008f0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00479] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008f2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0047a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008f4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0047b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008f6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0047c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008f8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0047d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008fa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0047e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008fc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0047f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h008fe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00480] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00900] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00481] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00902] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00482] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00904] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00483] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00906] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00484] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00908] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00485] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0090a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00486] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0090c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00487] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0090e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00488] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00910] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00489] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00912] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0048a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00914] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0048b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00916] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0048c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00918] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0048d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0091a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0048e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0091c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0048f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0091e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00490] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00920] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00491] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00922] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00492] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00924] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00493] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00926] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00494] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00928] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00495] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0092a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00496] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0092c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00497] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0092e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00498] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00930] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00499] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00932] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0049a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00934] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0049b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00936] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0049c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00938] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0049d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0093a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0049e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0093c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0049f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0093e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004a0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00940] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004a1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00942] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004a2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00944] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004a3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00946] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004a4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00948] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004a5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0094a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004a6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0094c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004a7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0094e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004a8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00950] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004a9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00952] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004aa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00954] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004ab] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00956] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004ac] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00958] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004ad] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0095a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004ae] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0095c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004af] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0095e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004b0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00960] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004b1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00962] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004b2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00964] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004b3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00966] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004b4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00968] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004b5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0096a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004b6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0096c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004b7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0096e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004b8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00970] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004b9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00972] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004ba] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00974] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004bb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00976] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004bc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00978] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004bd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0097a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004be] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0097c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004bf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0097e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004c0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00980] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004c1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00982] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004c2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00984] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004c3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00986] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004c4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00988] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004c5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0098a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004c6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0098c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004c7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0098e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004c8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00990] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004c9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00992] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004ca] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00994] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004cb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00996] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004cc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00998] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004cd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0099a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004ce] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0099c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004cf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0099e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004d0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009a0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004d1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009a2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004d2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009a4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004d3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009a6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004d4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009a8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004d5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009aa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004d6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009ac] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004d7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009ae] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004d8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009b0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004d9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009b2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004da] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009b4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004db] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009b6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004dc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009b8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004dd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009ba] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004de] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009bc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004df] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009be] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004e0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009c0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004e1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009c2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004e2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009c4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004e3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009c6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004e4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009c8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004e5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009ca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004e6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009cc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004e7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009ce] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004e8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009d0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004e9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009d2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004ea] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009d4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004eb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009d6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004ec] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009d8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004ed] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009da] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004ee] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009dc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004ef] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009de] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004f0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009e0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004f1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009e2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004f2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009e4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004f3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009e6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004f4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009e8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004f5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009ea] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004f6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009ec] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004f7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009ee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004f8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009f0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004f9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009f2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004fa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009f4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004fb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009f6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004fc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009f8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004fd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009fa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004fe] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009fc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004ff] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h009fe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00500] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a00] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00501] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a02] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00502] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a04] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00503] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a06] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00504] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a08] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00505] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a0a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00506] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a0c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00507] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a0e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00508] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a10] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00509] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a12] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0050a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a14] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0050b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a16] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0050c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a18] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0050d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a1a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0050e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a1c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0050f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a1e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00510] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a20] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00511] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a22] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00512] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a24] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00513] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a26] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00514] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a28] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00515] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a2a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00516] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a2c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00517] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a2e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00518] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a30] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00519] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a32] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0051a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a34] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0051b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a36] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0051c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a38] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0051d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a3a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0051e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a3c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0051f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a3e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00520] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a40] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00521] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a42] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00522] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a44] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00523] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a46] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00524] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a48] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00525] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a4a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00526] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a4c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00527] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a4e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00528] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a50] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00529] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a52] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0052a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a54] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0052b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a56] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0052c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a58] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0052d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a5a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0052e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a5c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0052f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a5e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00530] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a60] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00531] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a62] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00532] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a64] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00533] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a66] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00534] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a68] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00535] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a6a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00536] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a6c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00537] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a6e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00538] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a70] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00539] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a72] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0053a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a74] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0053b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a76] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0053c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a78] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0053d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a7a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0053e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a7c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0053f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a7e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00540] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a80] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00541] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a82] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00542] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a84] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00543] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a86] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00544] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a88] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00545] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a8a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00546] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a8c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00547] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a8e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00548] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a90] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00549] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a92] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0054a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a94] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0054b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a96] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0054c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a98] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0054d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a9a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0054e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a9c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0054f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00a9e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00550] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aa0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00551] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aa2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00552] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aa4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00553] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aa6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00554] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aa8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00555] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aaa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00556] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aac] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00557] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aae] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00558] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ab0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00559] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ab2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0055a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ab4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0055b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ab6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0055c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ab8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0055d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aba] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0055e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00abc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0055f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00abe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00560] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ac0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00561] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ac2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00562] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ac4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00563] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ac6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00564] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ac8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00565] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00566] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00acc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00567] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ace] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00568] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ad0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00569] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ad2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0056a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ad4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0056b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ad6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0056c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ad8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0056d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ada] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0056e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00adc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0056f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ade] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00570] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ae0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00571] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ae2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00572] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ae4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00573] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ae6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00574] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ae8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00575] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aea] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00576] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aec] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00577] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00aee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00578] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00af0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00579] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00af2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0057a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00af4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0057b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00af6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0057c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00af8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0057d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00afa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0057e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00afc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0057f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00afe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00580] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b00] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00581] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b02] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00582] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b04] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00583] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b06] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00584] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b08] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00585] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b0a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00586] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b0c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00587] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b0e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00588] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b10] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00589] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b12] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0058a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b14] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0058b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b16] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0058c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b18] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0058d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b1a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0058e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b1c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0058f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b1e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00590] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b20] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00591] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b22] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00592] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b24] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00593] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b26] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00594] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b28] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00595] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b2a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00596] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b2c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00597] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b2e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00598] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b30] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00599] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b32] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0059a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b34] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0059b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b36] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0059c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b38] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0059d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b3a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0059e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b3c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0059f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b3e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005a0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b40] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005a1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b42] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005a2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b44] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005a3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b46] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005a4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b48] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005a5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b4a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005a6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b4c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005a7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b4e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005a8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b50] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005a9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b52] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005aa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b54] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005ab] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b56] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005ac] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b58] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005ad] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b5a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005ae] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b5c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005af] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b5e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005b0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b60] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005b1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b62] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005b2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b64] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005b3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b66] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005b4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b68] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005b5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b6a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005b6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b6c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005b7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b6e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005b8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b70] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005b9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b72] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005ba] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b74] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005bb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b76] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005bc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b78] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005bd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b7a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005be] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b7c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005bf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b7e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005c0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b80] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005c1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b82] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005c2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b84] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005c3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b86] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005c4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b88] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005c5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b8a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005c6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b8c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005c7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b8e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005c8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b90] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005c9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b92] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005ca] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b94] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005cb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b96] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005cc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b98] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005cd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b9a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005ce] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b9c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005cf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00b9e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005d0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ba0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005d1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ba2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005d2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ba4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005d3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ba6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005d4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ba8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005d5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00baa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005d6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bac] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005d7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bae] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005d8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bb0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005d9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bb2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005da] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bb4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005db] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bb6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005dc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bb8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005dd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bba] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005de] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bbc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005df] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bbe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005e0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bc0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005e1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bc2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005e2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bc4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005e3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bc6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005e4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bc8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005e5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005e6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bcc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005e7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bce] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005e8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bd0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005e9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bd2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005ea] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bd4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005eb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bd6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005ec] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bd8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005ed] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bda] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005ee] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bdc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005ef] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bde] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005f0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00be0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005f1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00be2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005f2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00be4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005f3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00be6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005f4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00be8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005f5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bea] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005f6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bec] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005f7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005f8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bf0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005f9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bf2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005fa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bf4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005fb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bf6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005fc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bf8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005fd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bfa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005fe] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bfc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005ff] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00bfe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00600] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c00] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00601] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c02] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00602] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c04] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00603] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c06] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00604] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c08] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00605] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c0a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00606] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c0c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00607] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c0e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00608] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c10] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00609] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c12] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0060a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c14] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0060b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c16] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0060c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c18] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0060d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c1a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0060e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c1c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0060f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c1e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00610] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c20] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00611] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c22] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00612] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c24] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00613] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c26] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00614] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c28] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00615] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c2a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00616] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c2c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00617] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c2e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00618] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c30] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00619] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c32] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0061a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c34] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0061b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c36] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0061c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c38] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0061d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c3a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0061e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c3c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0061f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c3e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00620] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c40] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00621] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c42] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00622] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c44] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00623] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c46] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00624] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c48] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00625] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c4a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00626] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c4c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00627] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c4e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00628] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c50] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00629] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c52] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0062a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c54] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0062b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c56] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0062c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c58] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0062d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c5a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0062e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c5c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0062f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c5e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00630] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c60] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00631] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c62] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00632] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c64] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00633] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c66] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00634] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c68] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00635] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c6a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00636] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c6c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00637] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c6e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00638] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c70] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00639] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c72] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0063a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c74] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0063b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c76] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0063c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c78] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0063d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c7a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0063e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c7c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0063f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c7e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00640] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c80] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00641] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c82] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00642] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c84] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00643] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c86] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00644] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c88] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00645] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c8a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00646] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c8c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00647] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c8e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00648] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c90] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00649] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c92] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0064a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c94] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0064b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c96] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0064c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c98] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0064d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c9a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0064e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c9c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0064f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00c9e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00650] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ca0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00651] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ca2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00652] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ca4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00653] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ca6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00654] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ca8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00655] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00caa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00656] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cac] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00657] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cae] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00658] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cb0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00659] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cb2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0065a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cb4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0065b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cb6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0065c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cb8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0065d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cba] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0065e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cbc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0065f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cbe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00660] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cc0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00661] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cc2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00662] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cc4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00663] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cc6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00664] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cc8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00665] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00666] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ccc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00667] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cce] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00668] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cd0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00669] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cd2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0066a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cd4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0066b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cd6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0066c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cd8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0066d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cda] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0066e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cdc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0066f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cde] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00670] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ce0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00671] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ce2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00672] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ce4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00673] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ce6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00674] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ce8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00675] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cea] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00676] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cec] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00677] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00678] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cf0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00679] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cf2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0067a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cf4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0067b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cf6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0067c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cf8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0067d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cfa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0067e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cfc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0067f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00cfe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00680] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d00] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00681] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d02] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00682] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d04] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00683] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d06] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00684] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d08] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00685] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d0a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00686] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d0c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00687] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d0e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00688] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d10] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00689] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d12] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0068a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d14] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0068b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d16] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0068c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d18] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0068d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d1a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0068e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d1c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0068f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d1e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00690] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d20] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00691] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d22] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00692] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d24] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00693] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d26] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00694] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d28] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00695] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d2a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00696] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d2c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00697] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d2e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00698] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d30] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00699] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d32] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0069a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d34] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0069b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d36] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0069c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d38] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0069d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d3a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0069e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d3c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0069f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d3e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006a0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d40] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006a1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d42] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006a2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d44] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006a3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d46] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006a4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d48] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006a5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d4a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006a6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d4c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006a7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d4e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006a8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d50] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006a9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d52] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006aa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d54] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006ab] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d56] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006ac] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d58] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006ad] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d5a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006ae] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d5c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006af] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d5e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006b0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d60] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006b1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d62] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006b2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d64] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006b3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d66] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006b4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d68] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006b5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d6a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006b6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d6c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006b7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d6e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006b8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d70] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006b9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d72] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006ba] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d74] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006bb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d76] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006bc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d78] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006bd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d7a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006be] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d7c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006bf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d7e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006c0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d80] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006c1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d82] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006c2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d84] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006c3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d86] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006c4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d88] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006c5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d8a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006c6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d8c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006c7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d8e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006c8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d90] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006c9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d92] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006ca] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d94] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006cb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d96] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006cc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d98] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006cd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d9a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006ce] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d9c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006cf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00d9e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006d0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00da0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006d1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00da2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006d2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00da4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006d3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00da6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006d4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00da8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006d5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00daa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006d6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dac] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006d7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dae] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006d8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00db0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006d9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00db2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006da] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00db4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006db] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00db6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006dc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00db8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006dd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dba] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006de] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dbc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006df] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dbe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006e0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dc0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006e1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dc2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006e2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dc4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006e3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dc6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006e4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dc8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006e5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006e6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dcc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006e7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dce] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006e8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dd0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006e9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dd2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006ea] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dd4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006eb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dd6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006ec] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dd8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006ed] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dda] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006ee] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ddc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006ef] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dde] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006f0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00de0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006f1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00de2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006f2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00de4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006f3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00de6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006f4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00de8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006f5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dea] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006f6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dec] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006f7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006f8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00df0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006f9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00df2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006fa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00df4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006fb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00df6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006fc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00df8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006fd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dfa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006fe] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dfc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006ff] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00dfe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00700] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e00] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00701] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e02] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00702] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e04] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00703] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e06] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00704] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e08] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00705] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e0a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00706] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e0c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00707] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e0e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00708] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e10] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00709] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e12] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0070a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e14] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0070b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e16] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0070c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e18] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0070d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e1a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0070e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e1c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0070f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e1e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00710] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e20] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00711] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e22] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00712] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e24] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00713] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e26] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00714] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e28] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00715] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e2a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00716] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e2c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00717] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e2e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00718] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e30] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00719] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e32] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0071a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e34] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0071b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e36] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0071c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e38] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0071d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e3a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0071e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e3c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0071f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e3e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00720] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e40] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00721] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e42] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00722] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e44] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00723] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e46] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00724] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e48] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00725] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e4a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00726] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e4c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00727] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e4e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00728] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e50] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00729] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e52] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0072a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e54] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0072b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e56] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0072c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e58] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0072d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e5a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0072e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e5c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0072f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e5e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00730] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e60] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00731] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e62] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00732] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e64] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00733] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e66] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00734] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e68] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00735] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e6a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00736] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e6c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00737] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e6e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00738] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e70] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00739] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e72] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0073a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e74] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0073b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e76] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0073c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e78] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0073d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e7a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0073e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e7c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0073f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e7e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00740] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e80] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00741] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e82] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00742] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e84] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00743] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e86] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00744] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e88] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00745] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e8a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00746] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e8c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00747] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e8e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00748] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e90] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00749] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e92] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0074a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e94] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0074b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e96] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0074c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e98] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0074d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e9a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0074e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e9c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0074f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00e9e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00750] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ea0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00751] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ea2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00752] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ea4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00753] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ea6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00754] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ea8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00755] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eaa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00756] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eac] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00757] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eae] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00758] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eb0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00759] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eb2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0075a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eb4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0075b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eb6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0075c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eb8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0075d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eba] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0075e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ebc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0075f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ebe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00760] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ec0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00761] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ec2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00762] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ec4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00763] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ec6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00764] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ec8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00765] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00766] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ecc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00767] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ece] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00768] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ed0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00769] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ed2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0076a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ed4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0076b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ed6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0076c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ed8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0076d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eda] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0076e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00edc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0076f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ede] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00770] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ee0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00771] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ee2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00772] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ee4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00773] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ee6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00774] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ee8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00775] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eea] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00776] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eec] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00777] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00eee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00778] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ef0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00779] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ef2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0077a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ef4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0077b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ef6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0077c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ef8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0077d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00efa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0077e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00efc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0077f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00efe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00780] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f00] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00781] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f02] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00782] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f04] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00783] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f06] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00784] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f08] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00785] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f0a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00786] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f0c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00787] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f0e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00788] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f10] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00789] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f12] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0078a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f14] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0078b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f16] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0078c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f18] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0078d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f1a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0078e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f1c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0078f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f1e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00790] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f20] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00791] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f22] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00792] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f24] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00793] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f26] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00794] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f28] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00795] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f2a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00796] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f2c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00797] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f2e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00798] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f30] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00799] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f32] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0079a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f34] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0079b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f36] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0079c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f38] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0079d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f3a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0079e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f3c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0079f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f3e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007a0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f40] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007a1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f42] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007a2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f44] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007a3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f46] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007a4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f48] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007a5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f4a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007a6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f4c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007a7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f4e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007a8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f50] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007a9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f52] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007aa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f54] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007ab] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f56] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007ac] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f58] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007ad] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f5a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007ae] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f5c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007af] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f5e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007b0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f60] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007b1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f62] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007b2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f64] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007b3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f66] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007b4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f68] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007b5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f6a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007b6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f6c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007b7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f6e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007b8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f70] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007b9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f72] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007ba] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f74] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007bb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f76] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007bc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f78] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007bd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f7a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007be] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f7c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007bf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f7e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007c0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f80] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007c1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f82] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007c2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f84] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007c3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f86] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007c4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f88] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007c5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f8a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007c6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f8c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007c7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f8e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007c8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f90] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007c9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f92] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007ca] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f94] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007cb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f96] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007cc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f98] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007cd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f9a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007ce] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f9c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007cf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00f9e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007d0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fa0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007d1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fa2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007d2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fa4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007d3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fa6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007d4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fa8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007d5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00faa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007d6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fac] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007d7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fae] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007d8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fb0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007d9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fb2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007da] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fb4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007db] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fb6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007dc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fb8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007dd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fba] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007de] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fbc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007df] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fbe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007e0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fc0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007e1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fc2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007e2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fc4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007e3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fc6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007e4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fc8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007e5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007e6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fcc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007e7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fce] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007e8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fd0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007e9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fd2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007ea] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fd4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007eb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fd6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007ec] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fd8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007ed] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fda] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007ee] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fdc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007ef] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fde] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007f0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fe0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007f1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fe2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007f2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fe4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007f3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fe6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007f4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fe8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007f5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fea] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007f6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fec] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007f7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00fee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007f8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ff0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007f9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ff2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007fa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ff4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007fb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ff6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007fc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ff8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007fd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ffa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007fe] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ffc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007ff] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h00ffe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00800] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01000] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00801] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01002] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00802] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01004] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00803] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01006] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00804] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01008] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00805] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0100a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00806] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0100c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00807] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0100e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00808] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01010] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00809] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01012] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0080a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01014] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0080b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01016] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0080c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01018] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0080d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0101a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0080e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0101c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0080f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0101e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00810] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01020] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00811] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01022] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00812] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01024] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00813] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01026] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00814] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01028] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00815] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0102a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00816] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0102c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00817] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0102e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00818] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01030] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00819] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01032] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0081a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01034] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0081b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01036] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0081c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01038] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0081d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0103a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0081e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0103c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0081f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0103e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00820] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01040] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00821] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01042] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00822] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01044] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00823] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01046] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00824] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01048] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00825] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0104a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00826] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0104c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00827] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0104e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00828] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01050] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00829] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01052] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0082a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01054] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0082b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01056] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0082c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01058] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0082d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0105a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0082e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0105c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0082f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0105e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00830] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01060] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00831] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01062] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00832] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01064] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00833] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01066] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00834] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01068] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00835] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0106a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00836] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0106c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00837] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0106e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00838] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01070] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00839] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01072] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0083a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01074] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0083b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01076] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0083c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01078] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0083d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0107a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0083e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0107c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0083f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0107e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00840] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01080] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00841] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01082] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00842] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01084] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00843] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01086] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00844] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01088] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00845] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0108a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00846] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0108c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00847] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0108e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00848] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01090] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00849] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01092] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0084a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01094] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0084b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01096] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0084c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01098] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0084d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0109a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0084e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0109c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0084f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0109e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00850] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010a0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00851] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010a2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00852] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010a4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00853] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010a6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00854] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010a8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00855] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010aa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00856] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010ac] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00857] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010ae] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00858] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010b0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00859] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010b2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0085a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010b4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0085b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010b6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0085c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010b8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0085d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010ba] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0085e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010bc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0085f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010be] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00860] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010c0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00861] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010c2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00862] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010c4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00863] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010c6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00864] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010c8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00865] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010ca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00866] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010cc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00867] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010ce] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00868] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010d0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00869] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010d2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0086a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010d4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0086b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010d6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0086c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010d8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0086d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010da] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0086e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010dc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0086f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010de] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00870] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010e0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00871] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010e2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00872] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010e4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00873] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010e6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00874] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010e8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00875] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010ea] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00876] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010ec] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00877] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010ee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00878] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010f0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00879] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010f2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0087a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010f4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0087b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010f6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0087c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010f8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0087d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010fa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0087e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010fc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0087f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h010fe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00880] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01100] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00881] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01102] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00882] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01104] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00883] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01106] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00884] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01108] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00885] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0110a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00886] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0110c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00887] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0110e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00888] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01110] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00889] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01112] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0088a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01114] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0088b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01116] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0088c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01118] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0088d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0111a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0088e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0111c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0088f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0111e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00890] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01120] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00891] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01122] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00892] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01124] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00893] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01126] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00894] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01128] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00895] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0112a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00896] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0112c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00897] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0112e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00898] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01130] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00899] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01132] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0089a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01134] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0089b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01136] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0089c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01138] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0089d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0113a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0089e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0113c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0089f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0113e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008a0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01140] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008a1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01142] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008a2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01144] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008a3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01146] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008a4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01148] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008a5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0114a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008a6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0114c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008a7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0114e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008a8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01150] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008a9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01152] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008aa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01154] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008ab] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01156] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008ac] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01158] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008ad] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0115a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008ae] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0115c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008af] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0115e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008b0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01160] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008b1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01162] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008b2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01164] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008b3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01166] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008b4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01168] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008b5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0116a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008b6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0116c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008b7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0116e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008b8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01170] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008b9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01172] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008ba] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01174] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008bb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01176] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008bc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01178] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008bd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0117a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008be] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0117c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008bf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0117e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008c0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01180] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008c1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01182] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008c2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01184] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008c3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01186] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008c4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01188] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008c5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0118a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008c6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0118c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008c7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0118e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008c8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01190] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008c9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01192] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008ca] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01194] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008cb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01196] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008cc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01198] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008cd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0119a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008ce] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0119c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008cf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0119e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008d0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011a0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008d1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011a2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008d2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011a4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008d3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011a6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008d4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011a8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008d5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011aa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008d6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011ac] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008d7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011ae] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008d8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011b0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008d9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011b2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008da] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011b4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008db] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011b6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008dc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011b8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008dd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011ba] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008de] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011bc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008df] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011be] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008e0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011c0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008e1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011c2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008e2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011c4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008e3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011c6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008e4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011c8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008e5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011ca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008e6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011cc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008e7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011ce] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008e8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011d0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008e9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011d2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008ea] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011d4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008eb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011d6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008ec] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011d8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008ed] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011da] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008ee] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011dc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008ef] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011de] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008f0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011e0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008f1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011e2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008f2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011e4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008f3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011e6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008f4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011e8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008f5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011ea] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008f6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011ec] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008f7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011ee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008f8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011f0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008f9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011f2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008fa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011f4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008fb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011f6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008fc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011f8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008fd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011fa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008fe] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011fc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008ff] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h011fe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00900] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01200] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00901] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01202] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00902] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01204] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00903] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01206] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00904] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01208] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00905] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0120a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00906] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0120c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00907] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0120e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00908] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01210] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00909] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01212] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0090a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01214] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0090b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01216] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0090c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01218] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0090d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0121a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0090e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0121c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0090f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0121e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00910] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01220] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00911] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01222] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00912] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01224] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00913] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01226] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00914] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01228] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00915] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0122a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00916] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0122c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00917] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0122e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00918] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01230] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00919] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01232] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0091a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01234] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0091b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01236] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0091c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01238] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0091d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0123a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0091e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0123c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0091f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0123e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00920] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01240] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00921] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01242] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00922] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01244] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00923] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01246] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00924] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01248] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00925] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0124a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00926] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0124c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00927] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0124e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00928] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01250] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00929] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01252] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0092a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01254] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0092b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01256] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0092c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01258] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0092d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0125a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0092e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0125c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0092f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0125e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00930] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01260] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00931] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01262] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00932] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01264] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00933] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01266] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00934] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01268] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00935] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0126a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00936] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0126c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00937] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0126e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00938] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01270] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00939] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01272] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0093a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01274] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0093b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01276] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0093c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01278] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0093d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0127a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0093e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0127c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0093f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0127e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00940] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01280] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00941] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01282] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00942] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01284] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00943] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01286] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00944] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01288] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00945] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0128a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00946] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0128c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00947] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0128e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00948] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01290] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00949] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01292] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0094a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01294] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0094b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01296] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0094c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01298] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0094d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0129a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0094e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0129c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0094f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0129e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00950] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012a0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00951] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012a2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00952] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012a4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00953] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012a6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00954] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012a8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00955] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012aa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00956] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012ac] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00957] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012ae] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00958] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012b0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00959] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012b2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0095a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012b4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0095b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012b6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0095c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012b8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0095d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012ba] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0095e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012bc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0095f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012be] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00960] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012c0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00961] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012c2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00962] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012c4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00963] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012c6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00964] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012c8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00965] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012ca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00966] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012cc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00967] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012ce] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00968] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012d0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00969] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012d2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0096a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012d4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0096b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012d6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0096c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012d8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0096d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012da] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0096e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012dc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0096f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012de] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00970] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012e0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00971] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012e2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00972] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012e4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00973] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012e6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00974] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012e8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00975] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012ea] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00976] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012ec] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00977] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012ee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00978] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012f0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00979] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012f2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0097a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012f4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0097b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012f6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0097c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012f8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0097d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012fa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0097e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012fc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0097f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h012fe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00980] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01300] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00981] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01302] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00982] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01304] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00983] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01306] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00984] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01308] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00985] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0130a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00986] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0130c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00987] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0130e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00988] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01310] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00989] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01312] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0098a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01314] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0098b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01316] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0098c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01318] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0098d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0131a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0098e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0131c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0098f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0131e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00990] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01320] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00991] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01322] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00992] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01324] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00993] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01326] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00994] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01328] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00995] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0132a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00996] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0132c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00997] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0132e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00998] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01330] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00999] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01332] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0099a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01334] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0099b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01336] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0099c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01338] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0099d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0133a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0099e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0133c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0099f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0133e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009a0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01340] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009a1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01342] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009a2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01344] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009a3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01346] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009a4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01348] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009a5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0134a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009a6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0134c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009a7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0134e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009a8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01350] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009a9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01352] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009aa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01354] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009ab] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01356] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009ac] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01358] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009ad] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0135a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009ae] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0135c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009af] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0135e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009b0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01360] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009b1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01362] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009b2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01364] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009b3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01366] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009b4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01368] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009b5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0136a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009b6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0136c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009b7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0136e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009b8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01370] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009b9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01372] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009ba] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01374] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009bb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01376] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009bc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01378] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009bd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0137a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009be] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0137c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009bf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0137e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009c0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01380] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009c1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01382] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009c2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01384] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009c3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01386] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009c4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01388] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009c5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0138a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009c6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0138c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009c7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0138e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009c8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01390] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009c9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01392] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009ca] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01394] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009cb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01396] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009cc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01398] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009cd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0139a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009ce] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0139c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009cf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0139e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009d0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013a0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009d1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013a2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009d2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013a4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009d3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013a6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009d4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013a8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009d5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013aa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009d6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013ac] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009d7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013ae] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009d8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013b0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009d9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013b2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009da] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013b4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009db] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013b6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009dc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013b8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009dd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013ba] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009de] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013bc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009df] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013be] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009e0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013c0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009e1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013c2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009e2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013c4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009e3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013c6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009e4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013c8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009e5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013ca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009e6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013cc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009e7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013ce] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009e8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013d0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009e9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013d2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009ea] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013d4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009eb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013d6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009ec] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013d8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009ed] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013da] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009ee] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013dc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009ef] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013de] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009f0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013e0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009f1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013e2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009f2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013e4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009f3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013e6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009f4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013e8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009f5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013ea] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009f6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013ec] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009f7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013ee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009f8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013f0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009f9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013f2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009fa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013f4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009fb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013f6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009fc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013f8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009fd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013fa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009fe] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013fc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009ff] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h013fe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a00] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01400] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a01] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01402] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a02] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01404] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a03] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01406] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a04] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01408] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a05] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0140a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a06] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0140c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a07] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0140e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a08] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01410] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a09] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01412] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a0a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01414] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a0b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01416] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a0c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01418] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a0d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0141a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a0e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0141c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a0f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0141e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a10] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01420] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a11] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01422] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a12] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01424] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a13] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01426] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a14] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01428] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a15] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0142a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a16] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0142c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a17] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0142e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a18] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01430] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a19] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01432] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a1a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01434] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a1b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01436] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a1c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01438] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a1d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0143a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a1e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0143c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a1f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0143e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a20] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01440] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a21] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01442] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a22] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01444] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a23] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01446] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a24] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01448] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a25] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0144a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a26] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0144c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a27] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0144e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a28] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01450] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a29] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01452] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a2a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01454] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a2b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01456] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a2c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01458] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a2d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0145a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a2e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0145c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a2f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0145e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a30] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01460] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a31] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01462] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a32] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01464] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a33] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01466] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a34] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01468] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a35] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0146a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a36] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0146c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a37] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0146e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a38] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01470] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a39] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01472] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a3a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01474] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a3b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01476] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a3c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01478] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a3d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0147a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a3e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0147c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a3f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0147e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a40] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01480] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a41] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01482] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a42] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01484] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a43] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01486] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a44] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01488] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a45] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0148a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a46] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0148c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a47] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0148e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a48] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01490] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a49] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01492] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a4a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01494] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a4b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01496] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a4c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01498] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a4d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0149a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a4e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0149c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a4f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0149e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a50] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014a0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a51] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014a2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a52] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014a4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a53] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014a6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a54] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014a8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a55] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014aa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a56] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014ac] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a57] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014ae] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a58] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014b0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a59] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014b2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a5a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014b4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a5b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014b6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a5c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014b8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a5d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014ba] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a5e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014bc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a5f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014be] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a60] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014c0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a61] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014c2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a62] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014c4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a63] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014c6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a64] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014c8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a65] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014ca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a66] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014cc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a67] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014ce] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a68] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014d0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a69] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014d2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a6a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014d4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a6b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014d6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a6c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014d8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a6d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014da] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a6e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014dc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a6f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014de] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a70] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014e0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a71] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014e2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a72] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014e4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a73] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014e6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a74] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014e8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a75] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014ea] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a76] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014ec] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a77] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014ee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a78] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014f0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a79] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014f2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a7a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014f4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a7b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014f6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a7c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014f8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a7d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014fa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a7e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014fc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a7f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h014fe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a80] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01500] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a81] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01502] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a82] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01504] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a83] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01506] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a84] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01508] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a85] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0150a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a86] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0150c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a87] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0150e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a88] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01510] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a89] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01512] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a8a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01514] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a8b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01516] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a8c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01518] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a8d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0151a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a8e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0151c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a8f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0151e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a90] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01520] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a91] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01522] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a92] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01524] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a93] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01526] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a94] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01528] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a95] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0152a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a96] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0152c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a97] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0152e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a98] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01530] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a99] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01532] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a9a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01534] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a9b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01536] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a9c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01538] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a9d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0153a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a9e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0153c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a9f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0153e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aa0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01540] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aa1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01542] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aa2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01544] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aa3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01546] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aa4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01548] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aa5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0154a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aa6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0154c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aa7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0154e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aa8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01550] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aa9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01552] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aaa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01554] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aab] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01556] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aac] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01558] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aad] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0155a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aae] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0155c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aaf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0155e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ab0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01560] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ab1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01562] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ab2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01564] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ab3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01566] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ab4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01568] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ab5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0156a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ab6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0156c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ab7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0156e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ab8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01570] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ab9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01572] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aba] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01574] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00abb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01576] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00abc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01578] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00abd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0157a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00abe] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0157c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00abf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0157e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ac0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01580] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ac1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01582] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ac2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01584] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ac3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01586] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ac4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01588] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ac5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0158a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ac6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0158c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ac7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0158e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ac8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01590] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ac9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01592] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aca] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01594] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00acb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01596] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00acc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01598] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00acd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0159a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ace] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0159c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00acf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0159e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ad0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015a0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ad1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015a2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ad2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015a4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ad3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015a6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ad4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015a8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ad5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015aa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ad6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015ac] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ad7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015ae] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ad8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015b0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ad9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015b2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ada] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015b4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00adb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015b6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00adc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015b8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00add] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015ba] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ade] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015bc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00adf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015be] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ae0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015c0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ae1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015c2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ae2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015c4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ae3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015c6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ae4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015c8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ae5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015ca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ae6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015cc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ae7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015ce] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ae8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015d0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ae9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015d2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aea] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015d4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aeb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015d6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aec] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015d8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aed] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015da] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aee] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015dc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aef] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015de] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00af0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015e0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00af1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015e2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00af2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015e4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00af3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015e6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00af4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015e8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00af5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015ea] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00af6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015ec] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00af7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015ee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00af8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015f0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00af9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015f2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00afa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015f4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00afb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015f6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00afc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015f8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00afd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015fa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00afe] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015fc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aff] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h015fe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b00] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01600] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b01] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01602] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b02] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01604] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b03] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01606] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b04] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01608] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b05] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0160a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b06] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0160c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b07] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0160e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b08] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01610] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b09] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01612] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b0a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01614] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b0b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01616] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b0c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01618] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b0d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0161a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b0e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0161c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b0f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0161e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b10] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01620] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b11] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01622] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b12] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01624] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b13] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01626] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b14] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01628] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b15] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0162a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b16] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0162c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b17] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0162e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b18] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01630] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b19] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01632] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b1a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01634] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b1b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01636] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b1c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01638] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b1d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0163a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b1e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0163c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b1f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0163e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b20] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01640] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b21] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01642] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b22] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01644] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b23] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01646] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b24] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01648] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b25] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0164a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b26] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0164c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b27] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0164e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b28] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01650] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b29] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01652] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b2a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01654] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b2b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01656] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b2c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01658] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b2d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0165a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b2e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0165c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b2f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0165e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b30] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01660] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b31] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01662] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b32] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01664] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b33] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01666] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b34] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01668] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b35] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0166a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b36] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0166c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b37] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0166e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b38] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01670] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b39] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01672] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b3a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01674] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b3b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01676] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b3c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01678] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b3d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0167a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b3e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0167c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b3f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0167e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b40] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01680] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b41] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01682] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b42] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01684] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b43] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01686] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b44] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01688] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b45] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0168a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b46] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0168c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b47] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0168e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b48] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01690] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b49] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01692] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b4a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01694] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b4b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01696] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b4c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01698] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b4d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0169a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b4e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0169c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b4f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0169e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b50] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016a0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b51] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016a2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b52] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016a4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b53] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016a6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b54] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016a8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b55] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016aa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b56] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016ac] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b57] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016ae] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b58] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016b0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b59] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016b2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b5a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016b4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b5b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016b6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b5c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016b8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b5d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016ba] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b5e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016bc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b5f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016be] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b60] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016c0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b61] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016c2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b62] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016c4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b63] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016c6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b64] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016c8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b65] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016ca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b66] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016cc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b67] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016ce] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b68] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016d0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b69] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016d2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b6a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016d4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b6b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016d6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b6c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016d8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b6d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016da] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b6e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016dc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b6f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016de] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b70] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016e0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b71] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016e2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b72] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016e4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b73] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016e6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b74] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016e8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b75] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016ea] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b76] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016ec] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b77] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016ee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b78] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016f0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b79] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016f2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b7a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016f4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b7b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016f6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b7c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016f8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b7d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016fa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b7e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016fc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b7f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h016fe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b80] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01700] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b81] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01702] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b82] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01704] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b83] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01706] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b84] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01708] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b85] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0170a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b86] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0170c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b87] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0170e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b88] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01710] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b89] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01712] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b8a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01714] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b8b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01716] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b8c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01718] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b8d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0171a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b8e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0171c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b8f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0171e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b90] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01720] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b91] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01722] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b92] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01724] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b93] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01726] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b94] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01728] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b95] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0172a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b96] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0172c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b97] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0172e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b98] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01730] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b99] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01732] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b9a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01734] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b9b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01736] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b9c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01738] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b9d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0173a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b9e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0173c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b9f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0173e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ba0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01740] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ba1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01742] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ba2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01744] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ba3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01746] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ba4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01748] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ba5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0174a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ba6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0174c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ba7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0174e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ba8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01750] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ba9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01752] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00baa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01754] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bab] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01756] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bac] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01758] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bad] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0175a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bae] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0175c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00baf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0175e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bb0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01760] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bb1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01762] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bb2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01764] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bb3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01766] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bb4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01768] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bb5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0176a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bb6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0176c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bb7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0176e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bb8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01770] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bb9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01772] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bba] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01774] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bbb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01776] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bbc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01778] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bbd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0177a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bbe] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0177c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bbf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0177e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bc0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01780] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bc1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01782] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bc2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01784] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bc3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01786] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bc4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01788] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bc5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0178a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bc6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0178c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bc7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0178e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bc8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01790] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bc9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01792] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bca] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01794] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bcb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01796] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bcc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01798] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bcd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0179a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bce] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0179c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bcf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0179e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bd0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017a0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bd1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017a2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bd2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017a4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bd3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017a6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bd4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017a8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bd5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017aa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bd6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017ac] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bd7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017ae] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bd8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017b0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bd9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017b2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bda] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017b4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bdb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017b6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bdc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017b8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bdd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017ba] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bde] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017bc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bdf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017be] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00be0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017c0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00be1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017c2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00be2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017c4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00be3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017c6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00be4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017c8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00be5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017ca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00be6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017cc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00be7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017ce] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00be8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017d0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00be9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017d2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bea] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017d4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00beb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017d6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bec] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017d8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bed] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017da] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bee] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017dc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bef] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017de] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bf0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017e0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bf1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017e2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bf2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017e4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bf3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017e6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bf4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017e8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bf5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017ea] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bf6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017ec] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bf7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017ee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bf8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017f0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bf9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017f2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bfa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017f4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bfb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017f6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bfc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017f8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bfd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017fa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bfe] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017fc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bff] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h017fe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c00] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01800] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c01] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01802] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c02] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01804] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c03] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01806] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c04] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01808] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c05] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0180a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c06] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0180c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c07] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0180e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c08] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01810] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c09] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01812] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c0a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01814] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c0b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01816] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c0c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01818] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c0d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0181a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c0e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0181c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c0f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0181e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c10] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01820] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c11] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01822] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c12] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01824] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c13] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01826] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c14] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01828] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c15] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0182a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c16] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0182c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c17] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0182e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c18] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01830] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c19] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01832] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c1a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01834] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c1b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01836] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c1c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01838] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c1d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0183a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c1e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0183c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c1f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0183e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c20] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01840] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c21] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01842] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c22] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01844] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c23] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01846] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c24] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01848] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c25] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0184a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c26] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0184c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c27] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0184e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c28] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01850] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c29] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01852] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c2a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01854] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c2b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01856] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c2c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01858] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c2d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0185a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c2e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0185c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c2f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0185e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c30] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01860] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c31] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01862] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c32] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01864] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c33] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01866] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c34] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01868] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c35] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0186a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c36] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0186c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c37] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0186e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c38] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01870] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c39] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01872] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c3a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01874] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c3b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01876] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c3c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01878] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c3d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0187a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c3e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0187c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c3f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0187e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c40] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01880] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c41] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01882] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c42] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01884] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c43] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01886] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c44] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01888] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c45] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0188a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c46] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0188c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c47] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0188e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c48] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01890] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c49] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01892] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c4a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01894] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c4b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01896] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c4c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01898] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c4d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0189a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c4e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0189c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c4f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0189e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c50] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018a0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c51] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018a2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c52] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018a4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c53] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018a6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c54] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018a8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c55] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018aa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c56] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018ac] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c57] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018ae] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c58] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018b0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c59] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018b2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c5a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018b4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c5b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018b6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c5c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018b8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c5d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018ba] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c5e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018bc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c5f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018be] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c60] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018c0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c61] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018c2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c62] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018c4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c63] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018c6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c64] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018c8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c65] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018ca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c66] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018cc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c67] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018ce] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c68] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018d0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c69] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018d2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c6a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018d4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c6b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018d6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c6c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018d8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c6d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018da] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c6e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018dc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c6f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018de] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c70] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018e0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c71] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018e2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c72] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018e4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c73] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018e6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c74] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018e8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c75] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018ea] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c76] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018ec] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c77] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018ee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c78] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018f0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c79] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018f2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c7a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018f4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c7b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018f6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c7c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018f8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c7d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018fa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c7e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018fc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c7f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h018fe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c80] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01900] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c81] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01902] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c82] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01904] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c83] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01906] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c84] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01908] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c85] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0190a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c86] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0190c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c87] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0190e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c88] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01910] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c89] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01912] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c8a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01914] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c8b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01916] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c8c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01918] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c8d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0191a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c8e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0191c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c8f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0191e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c90] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01920] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c91] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01922] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c92] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01924] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c93] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01926] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c94] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01928] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c95] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0192a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c96] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0192c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c97] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0192e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c98] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01930] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c99] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01932] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c9a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01934] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c9b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01936] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c9c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01938] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c9d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0193a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c9e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0193c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c9f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0193e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ca0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01940] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ca1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01942] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ca2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01944] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ca3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01946] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ca4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01948] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ca5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0194a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ca6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0194c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ca7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0194e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ca8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01950] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ca9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01952] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00caa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01954] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cab] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01956] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cac] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01958] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cad] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0195a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cae] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0195c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00caf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0195e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cb0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01960] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cb1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01962] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cb2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01964] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cb3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01966] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cb4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01968] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cb5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0196a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cb6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0196c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cb7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0196e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cb8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01970] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cb9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01972] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cba] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01974] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cbb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01976] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cbc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01978] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cbd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0197a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cbe] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0197c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cbf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0197e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cc0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01980] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cc1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01982] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cc2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01984] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cc3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01986] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cc4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01988] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cc5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0198a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cc6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0198c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cc7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0198e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cc8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01990] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cc9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01992] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cca] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01994] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ccb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01996] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ccc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01998] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ccd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0199a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cce] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0199c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ccf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h0199e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cd0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019a0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cd1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019a2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cd2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019a4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cd3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019a6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cd4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019a8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cd5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019aa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cd6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019ac] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cd7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019ae] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cd8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019b0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cd9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019b2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cda] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019b4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cdb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019b6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cdc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019b8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cdd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019ba] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cde] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019bc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cdf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019be] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ce0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019c0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ce1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019c2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ce2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019c4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ce3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019c6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ce4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019c8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ce5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019ca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ce6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019cc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ce7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019ce] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ce8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019d0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ce9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019d2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cea] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019d4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ceb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019d6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cec] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019d8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ced] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019da] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cee] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019dc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cef] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019de] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cf0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019e0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cf1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019e2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cf2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019e4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cf3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019e6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cf4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019e8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cf5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019ea] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cf6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019ec] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cf7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019ee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cf8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019f0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cf9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019f2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cfa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019f4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cfb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019f6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cfc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019f8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cfd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019fa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cfe] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019fc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cff] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h019fe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d00] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a00] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d01] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a02] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d02] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a04] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d03] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a06] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d04] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a08] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d05] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a0a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d06] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a0c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d07] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a0e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d08] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a10] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d09] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a12] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d0a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a14] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d0b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a16] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d0c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a18] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d0d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a1a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d0e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a1c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d0f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a1e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d10] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a20] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d11] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a22] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d12] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a24] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d13] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a26] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d14] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a28] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d15] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a2a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d16] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a2c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d17] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a2e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d18] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a30] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d19] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a32] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d1a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a34] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d1b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a36] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d1c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a38] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d1d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a3a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d1e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a3c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d1f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a3e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d20] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a40] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d21] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a42] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d22] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a44] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d23] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a46] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d24] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a48] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d25] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a4a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d26] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a4c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d27] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a4e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d28] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a50] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d29] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a52] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d2a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a54] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d2b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a56] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d2c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a58] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d2d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a5a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d2e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a5c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d2f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a5e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d30] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a60] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d31] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a62] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d32] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a64] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d33] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a66] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d34] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a68] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d35] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a6a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d36] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a6c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d37] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a6e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d38] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a70] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d39] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a72] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d3a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a74] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d3b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a76] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d3c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a78] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d3d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a7a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d3e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a7c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d3f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a7e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d40] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a80] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d41] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a82] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d42] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a84] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d43] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a86] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d44] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a88] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d45] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a8a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d46] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a8c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d47] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a8e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d48] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a90] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d49] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a92] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d4a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a94] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d4b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a96] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d4c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a98] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d4d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a9a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d4e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a9c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d4f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01a9e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d50] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aa0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d51] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aa2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d52] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aa4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d53] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aa6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d54] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aa8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d55] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aaa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d56] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aac] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d57] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aae] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d58] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ab0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d59] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ab2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d5a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ab4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d5b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ab6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d5c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ab8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d5d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aba] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d5e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01abc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d5f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01abe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d60] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ac0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d61] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ac2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d62] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ac4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d63] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ac6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d64] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ac8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d65] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d66] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01acc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d67] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ace] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d68] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ad0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d69] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ad2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d6a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ad4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d6b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ad6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d6c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ad8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d6d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ada] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d6e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01adc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d6f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ade] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d70] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ae0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d71] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ae2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d72] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ae4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d73] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ae6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d74] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ae8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d75] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aea] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d76] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aec] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d77] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01aee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d78] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01af0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d79] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01af2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d7a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01af4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d7b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01af6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d7c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01af8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d7d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01afa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d7e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01afc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d7f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01afe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d80] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b00] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d81] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b02] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d82] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b04] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d83] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b06] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d84] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b08] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d85] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b0a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d86] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b0c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d87] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b0e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d88] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b10] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d89] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b12] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d8a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b14] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d8b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b16] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d8c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b18] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d8d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b1a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d8e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b1c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d8f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b1e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d90] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b20] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d91] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b22] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d92] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b24] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d93] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b26] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d94] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b28] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d95] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b2a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d96] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b2c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d97] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b2e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d98] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b30] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d99] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b32] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d9a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b34] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d9b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b36] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d9c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b38] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d9d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b3a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d9e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b3c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d9f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b3e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00da0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b40] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00da1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b42] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00da2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b44] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00da3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b46] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00da4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b48] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00da5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b4a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00da6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b4c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00da7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b4e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00da8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b50] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00da9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b52] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00daa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b54] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dab] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b56] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dac] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b58] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dad] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b5a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dae] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b5c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00daf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b5e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00db0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b60] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00db1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b62] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00db2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b64] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00db3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b66] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00db4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b68] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00db5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b6a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00db6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b6c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00db7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b6e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00db8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b70] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00db9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b72] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dba] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b74] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dbb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b76] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dbc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b78] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dbd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b7a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dbe] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b7c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dbf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b7e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dc0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b80] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dc1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b82] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dc2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b84] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dc3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b86] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dc4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b88] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dc5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b8a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dc6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b8c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dc7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b8e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dc8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b90] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dc9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b92] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dca] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b94] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dcb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b96] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dcc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b98] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dcd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b9a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dce] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b9c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dcf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01b9e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dd0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ba0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dd1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ba2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dd2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ba4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dd3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ba6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dd4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ba8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dd5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01baa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dd6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bac] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dd7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bae] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dd8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bb0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dd9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bb2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dda] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bb4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ddb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bb6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ddc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bb8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ddd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bba] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dde] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bbc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ddf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bbe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00de0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bc0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00de1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bc2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00de2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bc4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00de3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bc6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00de4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bc8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00de5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00de6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bcc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00de7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bce] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00de8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bd0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00de9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bd2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dea] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bd4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00deb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bd6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dec] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bd8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ded] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bda] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dee] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bdc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00def] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bde] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00df0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01be0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00df1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01be2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00df2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01be4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00df3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01be6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00df4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01be8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00df5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bea] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00df6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bec] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00df7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00df8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bf0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00df9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bf2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dfa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bf4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dfb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bf6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dfc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bf8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dfd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bfa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dfe] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bfc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dff] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01bfe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e00] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c00] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e01] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c02] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e02] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c04] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e03] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c06] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e04] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c08] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e05] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c0a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e06] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c0c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e07] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c0e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e08] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c10] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e09] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c12] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e0a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c14] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e0b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c16] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e0c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c18] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e0d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c1a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e0e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c1c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e0f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c1e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e10] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c20] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e11] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c22] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e12] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c24] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e13] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c26] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e14] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c28] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e15] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c2a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e16] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c2c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e17] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c2e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e18] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c30] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e19] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c32] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e1a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c34] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e1b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c36] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e1c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c38] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e1d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c3a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e1e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c3c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e1f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c3e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e20] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c40] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e21] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c42] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e22] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c44] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e23] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c46] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e24] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c48] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e25] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c4a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e26] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c4c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e27] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c4e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e28] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c50] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e29] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c52] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e2a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c54] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e2b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c56] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e2c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c58] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e2d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c5a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e2e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c5c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e2f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c5e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e30] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c60] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e31] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c62] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e32] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c64] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e33] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c66] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e34] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c68] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e35] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c6a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e36] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c6c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e37] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c6e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e38] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c70] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e39] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c72] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e3a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c74] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e3b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c76] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e3c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c78] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e3d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c7a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e3e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c7c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e3f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c7e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e40] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c80] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e41] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c82] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e42] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c84] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e43] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c86] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e44] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c88] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e45] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c8a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e46] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c8c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e47] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c8e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e48] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c90] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e49] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c92] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e4a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c94] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e4b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c96] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e4c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c98] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e4d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c9a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e4e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c9c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e4f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01c9e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e50] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ca0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e51] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ca2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e52] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ca4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e53] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ca6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e54] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ca8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e55] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01caa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e56] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cac] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e57] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cae] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e58] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cb0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e59] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cb2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e5a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cb4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e5b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cb6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e5c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cb8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e5d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cba] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e5e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cbc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e5f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cbe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e60] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cc0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e61] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cc2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e62] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cc4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e63] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cc6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e64] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cc8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e65] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e66] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ccc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e67] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cce] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e68] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cd0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e69] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cd2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e6a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cd4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e6b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cd6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e6c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cd8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e6d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cda] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e6e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cdc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e6f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cde] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e70] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ce0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e71] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ce2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e72] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ce4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e73] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ce6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e74] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ce8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e75] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cea] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e76] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cec] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e77] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e78] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cf0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e79] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cf2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e7a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cf4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e7b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cf6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e7c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cf8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e7d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cfa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e7e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cfc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e7f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01cfe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e80] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d00] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e81] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d02] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e82] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d04] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e83] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d06] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e84] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d08] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e85] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d0a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e86] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d0c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e87] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d0e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e88] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d10] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e89] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d12] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e8a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d14] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e8b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d16] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e8c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d18] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e8d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d1a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e8e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d1c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e8f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d1e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e90] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d20] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e91] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d22] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e92] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d24] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e93] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d26] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e94] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d28] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e95] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d2a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e96] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d2c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e97] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d2e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e98] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d30] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e99] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d32] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e9a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d34] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e9b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d36] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e9c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d38] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e9d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d3a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e9e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d3c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e9f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d3e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ea0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d40] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ea1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d42] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ea2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d44] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ea3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d46] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ea4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d48] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ea5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d4a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ea6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d4c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ea7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d4e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ea8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d50] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ea9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d52] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eaa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d54] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eab] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d56] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eac] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d58] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ead] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d5a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eae] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d5c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eaf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d5e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eb0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d60] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eb1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d62] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eb2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d64] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eb3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d66] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eb4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d68] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eb5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d6a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eb6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d6c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eb7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d6e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eb8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d70] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eb9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d72] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eba] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d74] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ebb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d76] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ebc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d78] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ebd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d7a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ebe] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d7c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ebf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d7e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ec0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d80] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ec1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d82] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ec2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d84] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ec3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d86] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ec4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d88] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ec5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d8a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ec6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d8c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ec7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d8e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ec8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d90] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ec9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d92] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eca] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d94] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ecb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d96] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ecc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d98] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ecd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d9a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ece] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d9c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ecf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01d9e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ed0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01da0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ed1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01da2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ed2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01da4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ed3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01da6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ed4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01da8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ed5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01daa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ed6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dac] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ed7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dae] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ed8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01db0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ed9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01db2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eda] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01db4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00edb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01db6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00edc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01db8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00edd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dba] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ede] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dbc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00edf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dbe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ee0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dc0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ee1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dc2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ee2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dc4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ee3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dc6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ee4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dc8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ee5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ee6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dcc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ee7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dce] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ee8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dd0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ee9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dd2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eea] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dd4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eeb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dd6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eec] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dd8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eed] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dda] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eee] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ddc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eef] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dde] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ef0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01de0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ef1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01de2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ef2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01de4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ef3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01de6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ef4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01de8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ef5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dea] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ef6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dec] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ef7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ef8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01df0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ef9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01df2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00efa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01df4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00efb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01df6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00efc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01df8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00efd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dfa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00efe] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dfc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eff] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01dfe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f00] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e00] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f01] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e02] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f02] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e04] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f03] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e06] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f04] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e08] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f05] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e0a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f06] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e0c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f07] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e0e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f08] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e10] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f09] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e12] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f0a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e14] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f0b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e16] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f0c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e18] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f0d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e1a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f0e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e1c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f0f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e1e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f10] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e20] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f11] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e22] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f12] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e24] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f13] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e26] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f14] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e28] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f15] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e2a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f16] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e2c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f17] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e2e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f18] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e30] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f19] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e32] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f1a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e34] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f1b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e36] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f1c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e38] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f1d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e3a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f1e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e3c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f1f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e3e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f20] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e40] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f21] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e42] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f22] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e44] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f23] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e46] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f24] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e48] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f25] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e4a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f26] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e4c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f27] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e4e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f28] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e50] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f29] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e52] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f2a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e54] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f2b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e56] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f2c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e58] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f2d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e5a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f2e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e5c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f2f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e5e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f30] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e60] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f31] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e62] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f32] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e64] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f33] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e66] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f34] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e68] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f35] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e6a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f36] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e6c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f37] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e6e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f38] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e70] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f39] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e72] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f3a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e74] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f3b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e76] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f3c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e78] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f3d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e7a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f3e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e7c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f3f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e7e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f40] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e80] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f41] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e82] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f42] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e84] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f43] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e86] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f44] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e88] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f45] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e8a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f46] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e8c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f47] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e8e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f48] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e90] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f49] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e92] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f4a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e94] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f4b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e96] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f4c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e98] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f4d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e9a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f4e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e9c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f4f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01e9e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f50] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ea0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f51] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ea2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f52] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ea4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f53] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ea6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f54] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ea8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f55] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eaa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f56] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eac] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f57] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eae] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f58] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eb0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f59] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eb2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f5a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eb4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f5b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eb6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f5c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eb8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f5d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eba] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f5e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ebc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f5f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ebe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f60] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ec0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f61] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ec2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f62] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ec4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f63] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ec6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f64] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ec8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f65] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f66] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ecc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f67] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ece] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f68] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ed0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f69] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ed2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f6a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ed4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f6b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ed6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f6c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ed8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f6d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eda] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f6e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01edc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f6f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ede] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f70] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ee0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f71] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ee2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f72] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ee4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f73] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ee6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f74] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ee8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f75] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eea] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f76] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eec] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f77] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01eee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f78] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ef0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f79] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ef2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f7a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ef4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f7b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ef6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f7c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ef8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f7d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01efa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f7e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01efc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f7f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01efe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f80] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f00] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f81] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f02] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f82] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f04] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f83] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f06] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f84] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f08] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f85] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f0a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f86] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f0c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f87] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f0e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f88] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f10] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f89] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f12] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f8a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f14] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f8b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f16] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f8c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f18] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f8d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f1a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f8e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f1c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f8f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f1e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f90] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f20] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f91] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f22] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f92] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f24] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f93] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f26] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f94] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f28] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f95] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f2a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f96] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f2c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f97] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f2e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f98] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f30] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f99] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f32] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f9a] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f34] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f9b] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f36] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f9c] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f38] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f9d] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f3a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f9e] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f3c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f9f] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f3e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fa0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f40] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fa1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f42] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fa2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f44] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fa3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f46] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fa4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f48] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fa5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f4a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fa6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f4c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fa7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f4e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fa8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f50] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fa9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f52] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00faa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f54] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fab] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f56] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fac] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f58] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fad] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f5a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fae] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f5c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00faf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f5e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fb0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f60] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fb1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f62] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fb2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f64] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fb3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f66] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fb4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f68] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fb5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f6a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fb6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f6c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fb7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f6e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fb8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f70] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fb9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f72] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fba] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f74] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fbb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f76] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fbc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f78] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fbd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f7a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fbe] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f7c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fbf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f7e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fc0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f80] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fc1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f82] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fc2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f84] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fc3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f86] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fc4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f88] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fc5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f8a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fc6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f8c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fc7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f8e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fc8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f90] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fc9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f92] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fca] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f94] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fcb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f96] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fcc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f98] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fcd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f9a] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fce] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f9c] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fcf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01f9e] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fd0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fa0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fd1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fa2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fd2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fa4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fd3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fa6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fd4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fa8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fd5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01faa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fd6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fac] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fd7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fae] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fd8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fb0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fd9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fb2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fda] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fb4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fdb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fb6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fdc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fb8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fdd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fba] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fde] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fbc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fdf] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fbe] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fe0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fc0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fe1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fc2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fe2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fc4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fe3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fc6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fe4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fc8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fe5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fca] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fe6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fcc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fe7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fce] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fe8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fd0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fe9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fd2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fea] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fd4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00feb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fd6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fec] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fd8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fed] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fda] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fee] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fdc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fef] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fde] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ff0] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fe0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ff1] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fe2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ff2] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fe4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ff3] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fe6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ff4] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fe8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ff5] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fea] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ff6] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fec] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ff7] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01fee] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ff8] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ff0] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ff9] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ff2] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ffa] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ff4] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ffb] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ff6] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ffc] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ff8] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ffd] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ffa] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ffe] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ffc] ;
//end
//always_comb begin // 
               I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fff] =  Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f['h01ffe] ;
//end
