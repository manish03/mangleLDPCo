 reg  ['h7fff:0] [$clog2('h7000+1)-1:0] I6eb3a3e04397efbe48cc2f5809bfcb98 ;
