              Ia7d34a5c48214f2a621b50e8ab83b8ed = 
          (!fgallag_sel[6]) ? 
                       I999768f7a0479b93e065e98bb8d71bb7: 
                       I6668f7bb8dc077f0ff1cac6d088185c3;
              Ia8a2a18441971a3b4fdc380de8e51678 = 
          (!fgallag_sel[6]) ? 
                       I99ce11aaea6da1dfb5d0567597b95ef4: 
                       I75b52e5dd015a0e0cfc2f7d453857ccd;
              I543147506272c69e234afd12a1d222ca = 
          (!fgallag_sel[6]) ? 
                       If01ebfc5e8f0038e0fd309e8b69f89e4: 
                       Id265f18fa76b685483b0694a5bb7ed43;
               I3b387622a3b87ba5f2e9cbe3841ea8eb =  0;
