         I0b93aca5ef7c84ffba0064eb4a53ec4f =   'h00380 ;
         Id37ee8cb85e5cd05bbe92dd90fd22777 =   'h0013a ;
         I41450c30addcb3bb1d2c1c036dc26d2f =   'h0011c ;
         I078a7802a3340b0c207a002a4046a4e3 =   'h000fa ;
         I5a33c28f0bc44840136790663423bd48 =   'h000e4 ;
         I777e21d17f74d2fe893977e1654e2c2d =   'h000d4 ;
         I0b457f5bce1ac08077d7c061655dd03f =   'h000c8 ;
         I8d508a837624b899a748b9152f4a787d =   'h000bd ;
         Ib226330c1225db758177402a9bcb4848 =   'h000b4 ;
         Ic9d6b4cdd3bfef73660bcd8319a9a7be =   'h000ad ;
         I8e094e0c0b13b04dee8f4f70fdee87c4 =   'h000a6 ;
         I5469abe94b035be8eb8713d061774eb5 =   'h0009f ;
         Ic6dd18ea6082a83222edb24cff9873da =   'h0009a ;
         If46aa2c29de75a5a44a4d629204b0963 =   'h00094 ;
         I86f471de37f4d7f2599425d1f7ae60b9 =   'h0008f ;
         Id4063c01903ecbf60f39cc2a65c5b73e =   'h0008b ;
         I1be4f732652b930e60cb6bf53fbb7132 =   'h00087 ;
         I64355c5e822a8d545c6fded925a984b6 =   'h00083 ;
         I865085332575d46654188a23e78a5ab5 =   'h0007f ;
         I5a3af3b67e01e19177daaa19b995b876 =   'h0007c ;
         Ic82f2a7d5019f0912c100d6336dfb3a8 =   'h00078 ;
         Icaa4f34ed9aaa9f1690a03ff7c374de4 =   'h00075 ;
         I7662e29bd142424284880f29b6d32038 =   'h00072 ;
         Ib9befe6fabe9ca87ddb96713b6c6e0d4 =   'h0006f ;
         I69bd49e2f242a3c2a32d182a32cf39f8 =   'h0006d ;
         I820044a9516905bcd63a9e6d98ec961d =   'h0006a ;
         I4b1cce4cb416fc1776b09254d2589bfe =   'h00068 ;
         I9cae305381503e9d92a4a8240bb2aac0 =   'h00065 ;
         I5a1301cdc00c141cd57b0c4b90d7dd7a =   'h00063 ;
         I98abd404eafd5efdc2a990f2760fb0d9 =   'h00061 ;
         I3e8a5169cec2e8120a2ba6b6dc0f5742 =   'h0005f ;
         I8b50f6cf167c2ec62d739f294512c324 =   'h0005d ;
         Ib0fffb83f9af51787fff93443dd10287 =   'h0005b ;
         I3e4d4fb93b28d431849e2dd307f91197 =   'h00059 ;
         I85b43efcd6de020aceb66ed5948fd901 =   'h00057 ;
         Ibf4c9739576bfc4c8d79dcdbdb629a6d =   'h00055 ;
         Ib96063e5603755f2354a15d573374fe0 =   'h00053 ;
         I5f07fe122c1bb26c6805a7f9d31218db =   'h00052 ;
         I0ed871a78ca4e2815ce45133571353a1 =   'h00050 ;
         Ib0ba4dc6303dade812ab25816938899e =   'h0004f ;
         Iea7ffe40a13deb5bfe2903c2965e4b63 =   'h0004d ;
         Iad7d1d253ed65347182adf53486dc1de =   'h0004b ;
         Ie4cc734fa69e1b46577b5df885ba3592 =   'h0004a ;
         I75554ec87598151940cd118e6ee59741 =   'h00049 ;
         Ifec751297668f80d860a9d6cc176e5f8 =   'h00047 ;
         I8fcbbdfd901920672268b4d6ca269849 =   'h00046 ;
         Id16656f72b76591b0bd03a3c2750684c =   'h00045 ;
         Iefa235bdb6e83afe1f793787d8dfca2f =   'h00043 ;
         Id4fc19c089fa63c1b901fb64c9c0e064 =   'h00042 ;
         Ib22f4bce6db16f279ad4085901174664 =   'h00041 ;
         I432b06e788f0047c5e66cac253186eca =   'h00040 ;
         I51d270bbc6e26272e0d6998307c33272 =   'h0003f ;
         I7f0c42c0c3c63ba11cdd3c26093bc3f5 =   'h0003d ;
         Ibe2e871186cde032e6ce4de65c0fbf75 =   'h0003c ;
         I9aaab4112c129c0563c8983c3cb372ba =   'h0003b ;
         I58b6cde8739d1e98ccbdd13b1a963c8f =   'h0003a ;
         I6d3d948976b4f578039a6dbaa8f08642 =   'h00039 ;
         I714b8ce615cf088e1ac52a7e22eb69df =   'h00038 ;
         I7672fb8749f7573c27144fffd1721ef7 =   'h00037 ;
         I5fa7ef4e8130409885342236b9f60fcd =   'h00036 ;
         I2ab7e691bb0a2f89f9cdbfbad80d7120 =   'h00035 ;
         Idc22eb4529d6e2f82fd6c23a113809da =   'h00034 ;
         I449ee1a89494568e104c9e29f66d4262 =   'h00033 ;
         I5e8f226f92643e61ad527be4f148de00 =   'h00033 ;
         I56a2b51825ae20cd1d9b434aa976b4dd =   'h00032 ;
         I580e0ae47b151812c4373cb1f268e4fe =   'h00031 ;
         I69e6eeed488ce445421bf458f3d1baaf =   'h00030 ;
         Ie3781ac0023a6e8091d66990ee3983ff =   'h0002f ;
         Ia6a4c1e9dcb6ab1ad0114e2da7a396bc =   'h0002e ;
         I91ed400a23a8aa771dbb930317b63466 =   'h0002e ;
         I15c7e1315b03dc87984424245b7e6dab =   'h0002d ;
         I4ae2e6ccef3d457713203f83eb10d60d =   'h0002c ;
         I08a273aa764a26045fd205007493d27a =   'h0002b ;
         Ifae99596becf8c2c7b69fc3e508a362a =   'h0002b ;
         Ib080cdead060a391cb67c54d97c7fb0b =   'h0002a ;
         Ie14db629163bf8c01b457b0df3bbb634 =   'h00029 ;
         Ib4c7a688661be990227b9902dcaa0721 =   'h00029 ;
         I4b33852fd89354d5eeaaf75dcb84e726 =   'h00028 ;
         I982d1672a39f86bf7da5bb7844bd57f9 =   'h00027 ;
         I29949584d0bbd464970883cc5724f8a4 =   'h00027 ;
         I03ec49385def83a3f577d847012976fc =   'h00026 ;
         I6bb12bbec43b6315c92ac22f43ef5a60 =   'h00025 ;
         I5c49372712967408ed819ba89624dc98 =   'h00025 ;
         I477fb86a2ad5f7ed4f225b0c85609bee =   'h00024 ;
         I67099935c6636fc80d472f193753ba55 =   'h00024 ;
         Icf692082f362b6bb08f320e2b27853c7 =   'h00023 ;
         Iae5385d0436fb1f5c949c0d1e8c3aa96 =   'h00022 ;
         I6951d4063e974375523406edae080570 =   'h00022 ;
         I54e637eae832d289eeba34eda853a657 =   'h00021 ;
         I89479946789730c4000d8166356cb964 =   'h00021 ;
         Ide9c460b12322a14105bd0484d4b9135 =   'h00020 ;
         Icb6633d32c69b880dea230dbae0896cd =   'h00020 ;
         Icc91b46df090bdc04306996433be6136 =   'h0001f ;
         I5ac7c7696f008ebbaf6019fa5ad57302 =   'h0001f ;
         Iab7f04bf5075b64439bff52f4779ca67 =   'h0001e ;
         I9c3e9f415a26edb9fedf25288a8fa453 =   'h0001e ;
         If0e39a30beb041d9c6b3c168e965a1af =   'h0001d ;
         Ibb59c086a89025918626f18799e73605 =   'h0001d ;
         Ic436ebe8aa48c3e6e935f6ce0b3f43d5 =   'h0001c ;
         I05239dbfe2cd2ef57477ecb654880bf4 =   'h0001c ;
         I1765216a10c88b6081f34198e8a5d26f =   'h0001b ;
         I37b9f75cb896a9e45a650b6dadd0b2ff =   'h0001b ;
         Ib9eeab393231e41cca081394b036bde6 =   'h0001b ;
         I499fb85792bd0c5a73022ac96ac27f13 =   'h0001a ;
         I3da1d9759bbad87b216b2bc8afc19f8e =   'h0001a ;
         Ie220bafbf40ee68b7591948b607fcaa0 =   'h00019 ;
         I34b7451c43eee381ab7b3f1e2a816b99 =   'h00019 ;
         I5a3b2767a2c2b41984b6f2a7f05dfcbc =   'h00018 ;
         I8ad73072ca340501c2b14404b9353b08 =   'h00018 ;
         Id3987a88bcc92458973c9ee529f52a56 =   'h00018 ;
         I49666607354671cb5d6ec9c3e6354f42 =   'h00017 ;
         I4da0ec3a6c662f7e76bd3f6c43b40722 =   'h00017 ;
         I039f5eff8e87d37a9cf7d754a82df849 =   'h00017 ;
         Ia6fa92e40471f5741d59b8515c67c24b =   'h00016 ;
         Ib4ce242cd8f88c4eb147129be5e6785c =   'h00016 ;
         Icc28fa9f2f20d09b439a9553b6e592fa =   'h00016 ;
         I8b4b437c18f15ae386e0c12371151913 =   'h00015 ;
         I7c34ca74407090b532ec5f0f65e5dc74 =   'h00015 ;
         I1f69904e43d7fb93f39873efcbbb558b =   'h00015 ;
         Ie1f3985459b6de4b08d14263f5b1aa18 =   'h00014 ;
         I3640c422ee8389926afc8108564b593b =   'h00014 ;
         Ie11fa9bb26231d41be8646707525d022 =   'h00014 ;
         Ibabb39952458fdb3127ed17f3909e043 =   'h00013 ;
         I8b1452ad1732c78b5397caddc0d43daa =   'h00013 ;
         I5adc876cca35af9714a2cb9ca0eb3ae1 =   'h00013 ;
         Ia2848a15587c0e23eef1de69c2a238b1 =   'h00012 ;
         Ic4119a74d5a813a98baede5515be91bc =   'h00012 ;
         Id3b3231272ef7b602acb9b7dcd5033e8 =   'h00012 ;
         I05e604f9ffc573b44538d9d864dd4e92 =   'h00012 ;
         I116d21ad2753927dbf389f373bb1a344 =   'h00011 ;
         I3805a70a8e257eeea2bdc179fba1d185 =   'h00011 ;
         Ie2d31cc4673f92faf8545984e9b52031 =   'h00011 ;
         I5bbb1e57ed53613e06ba3fe1cc4fd266 =   'h00010 ;
         Ic4e117cdda2e62382412fb1dfb9c850d =   'h00010 ;
         Iab33d8521b7118693333cb5f624f3904 =   'h00010 ;
         I4183bbdffed2418b9190d610ef9c85a5 =   'h00010 ;
         Ibee805f0c9d18428759c5ce6c61f4dee =   'h0000f ;
         Ic8255e62414174e60282be5b4d63c494 =   'h0000f ;
         Ie76911ee442cfab80022b3a534438350 =   'h0000f ;
         Ie9d09a2059dea91a80a00bdeb56940f2 =   'h0000f ;
         I86ecfe340941ed77c09fd4c69f5c272a =   'h0000e ;
         I511c8519304a31c10313838c1a053f85 =   'h0000e ;
         I8824abf0eb1a4d6b48a26abae23d0bff =   'h0000e ;
         I5d8953fa34cb14027d8375d02999f132 =   'h0000e ;
         I0d8e31fd51ec5b82c5206c307e0d53f7 =   'h0000e ;
         Ie1ea3318d114c790e9343e45555755ab =   'h0000d ;
         I495a91d95803df2b5cfca5053bf13a9b =   'h0000d ;
         Ide9b85fb8d57bdfbf9b8de9c18e9c5cd =   'h0000d ;
         I9cd4f5d3b10c25759e7993f9292a7390 =   'h0000d ;
         I5ea9ea2fd34572dc6833ccf368e52ccb =   'h0000d ;
         If3883c5646540cf78aee0589c3cd3022 =   'h0000c ;
         I61df05bea32eda79ed88930bbc84a13f =   'h0000c ;
         I7f1a2ad313f7af4a0f9eb4311f35ac12 =   'h0000c ;
         I685601482e2bded73351f69f3f5c21b2 =   'h0000c ;
         I484b91ff2256c38308e18bc50afed4ef =   'h0000c ;
         Id86467d5f10985a00ab65a8b029a8c82 =   'h0000b ;
         I56110e27931a312345e239eaf42781a2 =   'h0000b ;
         Iee57da8134718b73f0598a1884ecf424 =   'h0000b ;
         I7de0f163ab38efee6f9c2f362708f4a0 =   'h0000b ;
         Id397e815fb86c38fbb509692ec4dab0b =   'h0000b ;
         I2c5e75d48e9ca1a198d70980900bdc41 =   'h0000b ;
         If728db81c67f83aab133c8ceaa3a5c7b =   'h0000a ;
         I80d54bec914a5b89de0f5296459b152d =   'h0000a ;
         Ic99c4503bcbcad1099d0c26d3d9161b9 =   'h0000a ;
         I36119b67ff8b6471d47a6681ce27666b =   'h0000a ;
         I29103484cf42c813700bcc89a04146c8 =   'h0000a ;
         I3cef2dada2657f2140d9bdc43f83057b =   'h0000a ;
         I23abb9c83aae42b4b3a330f277ce3c5a =   'h00009 ;
         I79b6e7abe2503f1f13195584805dfcb6 =   'h00009 ;
         I4d042a3d0026d6b93b5b394034174b00 =   'h00009 ;
         I92d347131e209dc81a8321d27d38a69e =   'h00009 ;
         I79c6fd3ceb89abc93f49a67d913505ae =   'h00009 ;
         Ieb5038840ac4ab2ebdd9cf6222c15750 =   'h00009 ;
         Id81b8442322f6bdc3728f5459a830aeb =   'h00009 ;
         Ie3a852b81ccaf2d520d024dd989caa47 =   'h00008 ;
         I33b0bd948bf4495908c59c2d8f58cf2c =   'h00008 ;
         I09a19721c1644f9d1a6eaab84d8dddbe =   'h00008 ;
         I7065b10d4533cd967733d262d5e5777e =   'h00008 ;
         Ie75d8156129eb98d76783e3a6ade280e =   'h00008 ;
         Id3d25ba968ed699bd0b61ee32695edee =   'h00008 ;
         Ic560d519645177df445db05bad34e60e =   'h00008 ;
         Ia5720f57dcae8ac0b00ac4e4a3c89657 =   'h00008 ;
         I8cfcf912f60acfc715c63291a8c04729 =   'h00007 ;
         I6e5f2896cda9b8db3638d2b14cd6ac00 =   'h00007 ;
         I349da988b53307693f1e74a98fa686b6 =   'h00007 ;
         I47ec23a2e834f9c66f23f1e89eaf8679 =   'h00007 ;
         If03782abea72e6519c530636040d2291 =   'h00007 ;
         I512ac9f87b0fc7590f5434fc1e3f0372 =   'h00007 ;
         Ia0d98d1391069c78a92be189e60cec14 =   'h00007 ;
         Ic75a566d180368ca17dac6f967fe397d =   'h00007 ;
         Id9acaf5c4d2e0ff41de104ab47e77756 =   'h00007 ;
         Ic0a4f0637df63f87635fa78c21b2e99e =   'h00007 ;
         I4a61d91e170ec3b767be88ccb343f1ca =   'h00006 ;
         I12a049b431155546b8663137cc66bb9a =   'h00006 ;
         Ia019f222e96881e643709af1eb85011a =   'h00006 ;
         I09be79fb5efca2f460b667770755191b =   'h00006 ;
         I53f09f16c58b346a02997b021f882363 =   'h00006 ;
         I19b06a7f2c499994044c7dae5057d8a1 =   'h00006 ;
         Idb57cc9ee60ae36bf3c0117776a46d70 =   'h00006 ;
         I8c056925751f5cbfd61b1195817d25b1 =   'h00006 ;
         I8b92da1d7f30fa71249623b2bc87b462 =   'h00006 ;
         I020b3d3e1109655d6f795fd1ecc0a322 =   'h00006 ;
         If0e90362af64ee2a20b44f61aa766fb4 =   'h00005 ;
         Ie192f4f4088d17d1f7840213009ca3be =   'h00005 ;
         Ic72e05f3be735d52d9354cb8f43c1cc0 =   'h00005 ;
         I76141646fbd2efad1e121c6e08ac174e =   'h00005 ;
         I4ac4e1dec3801e462a47f80276b42397 =   'h00005 ;
         Ifefb5a209dde348266eb66805c0a7d2e =   'h00005 ;
         I92c5b8b76f0000bfffa0120f70f1991a =   'h00005 ;
         Ia94fc30c06efdb8ae6f388149d0dad5c =   'h00005 ;
         Ifdb73b22fe15d17de645cf8aa3da99e2 =   'h00005 ;
         I0b0e5a5734bd09dfad80a75fca5a763c =   'h00005 ;
         I73354f6673afdd64f94fe36e146cace0 =   'h00005 ;
         Ibe0a9cbd6da728e5f7e53081af472ea9 =   'h00005 ;
         I0edeae6c95ab6198047ded7f3b41efee =   'h00005 ;
         I473cf664c81394c8dab1d7f145b3804b =   'h00004 ;
         I7201b831890988766bc871eb0fa6e19d =   'h00004 ;
         Ic772d12c6a9f51ff6cb51bf7d54d1b21 =   'h00004 ;
         I16120aeff10370316421751a8f4e9505 =   'h00004 ;
         I77146070f8693370d971ec3a91e18f84 =   'h00004 ;
         I784fb1f69095ccb95c4bb705539970d8 =   'h00004 ;
         I2b2174ba9f0956782a3ab584fd11777a =   'h00004 ;
         I8f31a3afb2cc62773332f251278c1153 =   'h00004 ;
         Ib2cdf1583fe14fd7b16229572511fd7c =   'h00004 ;
         Ib04043dbfa7a17abbb728899e2459398 =   'h00004 ;
         Ib1eaa856a32de8ec5107bb40c8611700 =   'h00004 ;
         I04ac748d74a312f05ede4d4665042de6 =   'h00004 ;
         I70ef81ae751a5a7640ce2d4b0ac381c7 =   'h00004 ;
         I6c64c351f3b91838c0c3c25f3b06d201 =   'h00004 ;
         I146352e56b780e8cc0f10ac09cee3a2d =   'h00004 ;
         I966ffe439dac9390e18e84a65e4b6f11 =   'h00004 ;
         Ief16bdfba3e4ab746af015310ebbb6b8 =   'h00003 ;
         I0bb8923bb50a4fc7278094a514c79fb6 =   'h00003 ;
         I9e93a476f9669fb72f7999a6f0a05c16 =   'h00003 ;
         I0442bb2973db673118791e504be846e4 =   'h00003 ;
         Ib00b860d9b3981465aa3bb1f18cfc627 =   'h00003 ;
         I6ddab9f5aca020985482b76c25f2f81e =   'h00003 ;
         Idaa6aa87b597a3bcc6275f5f40444057 =   'h00003 ;
         I1e2ca5efd6735a6e241f9bcade3c2b60 =   'h00003 ;
         I50da8ce0a49993e0b7c16710e68da821 =   'h00003 ;
         Ief43e8dc88393e5a4015033c4021a8e5 =   'h00003 ;
         Idc4a8277aa0ac4ac35b9fa6b37f198f9 =   'h00003 ;
         I4f555c0f5b4b6f79ad394e0f196c8e9f =   'h00003 ;
         I7ddabcd95dfd2719f9e9925598e0cd80 =   'h00003 ;
         I007d2500c173825191e1243fc0758203 =   'h00003 ;
         Icee24ae7d32c16a6b5dd7089f6a63d18 =   'h00003 ;
         I0d5ad201c17a461d16a13675a0abf874 =   'h00003 ;
         I8cdcb20840d2cafe54bf1a40bb5fdb1c =   'h00003 ;
         I5dce978811c8a3680684eb168992afe7 =   'h00003 ;
         Ied4802a1ff9e40f97bd6ed7e5c9af351 =   'h00003 ;
         I54c34254efd813baebdff01bb5d9100a =   'h00003 ;
         Idf998c5802562dd8ba5cbbe2d8f4eca3 =   'h00003 ;
         I5140c93c2312dc879b408cce4db484d3 =   'h00003 ;
         I0110a5e1c6faa19f5d97ee4b4f763285 =   'h00002 ;
         I923c20fa85b752d9f31a3476e863c4c5 =   'h00002 ;
         I0eb29e587012701bb6ff57aa27d71ecc =   'h00002 ;
         Ib3668e1656878dd9ba2862b988011686 =   'h00002 ;
         Id7a758f960bb811f4ebb46662228c33c =   'h00002 ;
         I271fa5cfca7bbdafb091c3afcc3a7a41 =   'h00002 ;
         I864329472b61fb8580558865bcee6de1 =   'h00002 ;
         I78527503b3be9fca973ab9fb7f987f27 =   'h00002 ;
         I3f50edcfbffa653e39523fb6125d4fd5 =   'h00002 ;
         Ib5dd6975eedeed971f4aeaef77f28f1e =   'h00002 ;
         Ica77a9f6eb020b850ed2fa38021f33fe =   'h00002 ;
         I783f912ad4fff3731add8abca943629c =   'h00002 ;
         I1d7c0387f65da7d2ae51250edfc764de =   'h00002 ;
         I809a5efeed0db403579d08d520c2c9f1 =   'h00002 ;
         I7649e3988149218a8845000ffe68477f =   'h00002 ;
         Iad53806231a0e21d8b1e6b8a22fe3dfb =   'h00002 ;
         I9dcd325f9d12b6495d5b9f050af3c72e =   'h00002 ;
         Ib0d29b4d3693a1487dd507cd4610006f =   'h00002 ;
         Ide3d8fa67f76ce3a1762381698b59301 =   'h00002 ;
         I85818659b37457732130fef9b829758e =   'h00002 ;
         Ia8d5826890b3ca20e13dfa917300631b =   'h00002 ;
         I6b7c6fa01374134b230ebe6de1602785 =   'h00002 ;
         I4ebeea8273995c7ccb406a5cfedc3ef8 =   'h00002 ;
         I6521570d5f202bce800b1c49adf3f2ca =   'h00002 ;
         Iec61267ecdecf9fe305142fe095a21bb =   'h00002 ;
         Idd383af878d242f7be34d1c9d3efa0e8 =   'h00002 ;
         I44107557054891b33135a13058e00649 =   'h00002 ;
         I013496291a38e851842de8ea28b540ba =   'h00002 ;
         I54e8b21c865654527ee0720a72ef1cd0 =   'h00002 ;
         Ia40d6a1517b7b0a79c88646d209263dc =   'h00002 ;
         I1e10e22806a41d12b8c6328dbd9471df =   'h00002 ;
         If96824bc7f67bd2bce941ce96559867e =   'h00002 ;
         Ib252f7e32a3780abfb1a3e9285d0ed56 =   'h00001 ;
         I192fd55ca87b7cb2277aca900d015b04 =   'h00001 ;
         Ie973db372fd3127653d6c63a551a8c0c =   'h00001 ;
         I3446695b823b258ade0a7ac2aa9d61d7 =   'h00001 ;
         Iea584b5174273f9082695eec0d7a8ab1 =   'h00001 ;
         I6d7f0d64776ea582e326ca3b008f2b35 =   'h00001 ;
         Ifc32a10a9fcddca15eeef7d093d1401a =   'h00001 ;
         I84db677284b3e4bf9feddc2af30e9ad3 =   'h00001 ;
         Ia04c9bc6fc469c62a3645e0e691b3897 =   'h00001 ;
         Ib7457f82785a56cbcb5be6c0432641b7 =   'h00001 ;
         I42a4d0da5f0b890624310c94b32f1a27 =   'h00001 ;
         I08a589b0a34d88ac456d6cf40da0f5ae =   'h00001 ;
         I2f1e3460880499c961fcb244ca935f3b =   'h00001 ;
         Ie7f199c3586f87a1cdba687bd880497e =   'h00001 ;
         Ia3518f4b7c1b0aa2a864d5ce53158ce8 =   'h00001 ;
         Id2616c8625d0a75ea0946506034955ca =   'h00001 ;
         Ic3c6cbf9171a81f229a0fb9efd57b000 =   'h00001 ;
         If63bcb026b347506aff08fda75ac7c43 =   'h00001 ;
         Ia79c0c66c81e60806fe3df0addd5608d =   'h00001 ;
         I0695fe1981c8019decb9873e186934ae =   'h00001 ;
         Ic334a0e64e305848782becce03c85d2b =   'h00001 ;
         If737be717332ee2670d2c6736d9e0a2f =   'h00001 ;
         I66316458bfbdf6b24cdc0cd7396c84f6 =   'h00001 ;
         Ib23a5c11d42408a0f4a6d314a670da51 =   'h00001 ;
         I792738baad12910007da8123fa0ac415 =   'h00001 ;
         I64f43975f3065e3c7cfed15d5dbc8d72 =   'h00001 ;
         I4c0a3a24dcfac4edcdf29847761a8fb8 =   'h00001 ;
         I65fa0e67f8ee4669bba74ece0c565a0d =   'h00001 ;
         I6bea44d0467b461aa22c3ddcb1d8f886 =   'h00001 ;
         I582cb5f8b17099f479f297c5475542c1 =   'h00001 ;
         I6cba6eca48f199379e62726b4ac271f8 =   'h00001 ;
         I57cfe42eafe8357ec85906472dec3f36 =   'h00001 ;
         Iec7bf02aeaa8630497275c7eccab7667 =   'h00001 ;
         I388c7af9494f4c425621d3abfdf72b63 =   'h00001 ;
         I2622bb3685a7d6a297506eac3efb9c08 =   'h00001 ;
         If025bad83549d872a3fc9c44248174c8 =   'h00001 ;
         I3440574538a5d7dd250fbc98d574548b =   'h00001 ;
         Ibe30f2ceb078297737ce1444c1e6c524 =   'h00001 ;
         Ifbd6f1ac3bb594aad652d4e3cac018e1 =   'h00001 ;
         Ie41d26b8a9ac93a09ece53b2af8c855e =   'h00001 ;
         I497c3961e446544a8031e8013ca80ad5 =   'h00001 ;
         I6ab9d8eb7b8e3454b01a8e67a410624c =   'h00001 ;
         Icd351f2625b163cee904fa4e446d0cc4 =   'h00001 ;
         I79c9be2982685762d0907583f9f459e2 =   'h00001 ;
         Idc20427e979f3d5c03d7dd947cb4df84 =   'h00001 ;
         Ie8abbb597c8132b8e23936a5bc035041 =   'h00001 ;
         I42b0c89a558950f658440d8f9916b42f =   'h00001 ;
         I5a4d5a128b1fedabfdc39cb019359106 =   'h00001 ;
         I8227a9907c39647a4cef8e883d487913 =   'h00001 ;
         Icb2a399b8ac8449ff9ff8e5986aac03d =   'h00001 ;
         I933a5eb08d4d1445f167a74db5fbdc75 =   'h00001 ;
         I9c046caddde3b171774d3eba258190f0 =   'h00001 ;
         Ic8f12fefb9c055923e2842aeca48765f =   'h00001 ;
         I26631e7940eb983e49a9313da628e23a =   'h00001 ;
         I7fac6686ca9a63213ec3cdee4b812daa =   'h00001 ;
         I1960eba710ca20ef749501b02fd3b0bd =   'h00001 ;
         Ie1f5cc89163ee091f938a4c3edaca65b =   'h00001 ;
         I63e7cf958a0de50d3299d2077d8cb192 =   'h00001 ;
         I50c2132c2b5e60af7ba2b9be8c90d9a4 =   'h00001 ;
         If1243756e31d0a56b6666cad5b21f731 =   'h00001 ;
         I92c03e59c3f96f63800051762f6949c0 =   'h00001 ;
         I488d337ed967adebd6c580b7203991b5 =   'h00001 ;
         I32aa0d9a082eb6a595467f3c7f36a3f7 =   'h00001 ;
         Iec440f37d189fbcd4c06cf34344c4439 =   'h00001 ;
         I66d815daa51bcda0d549dbcc9c027195 =   'h00001 ;
         I192d10feae906d5ef90b4a90398d3ced =   'h00001 ;
         I1d8d269f64d0d3041bc69d879a3654ab =   'h00001 ;
         I5fce715f064098fe4685479aede832e7 =   'h00001 ;
         I1b65989684c087f328e3fb58d3a3395e =   'h00001 ;
         I5352562c002801df06f847362d347180 =   'h00001 ;
         I176397bab05ee39f7d54a28c5f74c3cc =   'h00001 ;
