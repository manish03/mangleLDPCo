//`include "GF2_LDPC_fgallag_0x00009_assign_inc.sv"
//always_comb begin
              If9057226a42b596a6dd2c84a37efff79['h00000] = 
          (!fgallag_sel['h00009]) ? 
                       Icff8af1f5c3ae89ef95ed8451273154b['h00000] : //%
                       Icff8af1f5c3ae89ef95ed8451273154b['h00001] ;
//end
//always_comb begin
              If9057226a42b596a6dd2c84a37efff79['h00001] = 
          (!fgallag_sel['h00009]) ? 
                       Icff8af1f5c3ae89ef95ed8451273154b['h00002] : //%
                       Icff8af1f5c3ae89ef95ed8451273154b['h00003] ;
//end
//always_comb begin
              If9057226a42b596a6dd2c84a37efff79['h00002] = 
          (!fgallag_sel['h00009]) ? 
                       Icff8af1f5c3ae89ef95ed8451273154b['h00004] : //%
                       Icff8af1f5c3ae89ef95ed8451273154b['h00005] ;
//end
//always_comb begin
              If9057226a42b596a6dd2c84a37efff79['h00003] = 
          (!fgallag_sel['h00009]) ? 
                       Icff8af1f5c3ae89ef95ed8451273154b['h00006] : //%
                       Icff8af1f5c3ae89ef95ed8451273154b['h00007] ;
//end
//always_comb begin
              If9057226a42b596a6dd2c84a37efff79['h00004] = 
          (!fgallag_sel['h00009]) ? 
                       Icff8af1f5c3ae89ef95ed8451273154b['h00008] : //%
                       Icff8af1f5c3ae89ef95ed8451273154b['h00009] ;
//end
//always_comb begin
              If9057226a42b596a6dd2c84a37efff79['h00005] = 
          (!fgallag_sel['h00009]) ? 
                       Icff8af1f5c3ae89ef95ed8451273154b['h0000a] : //%
                       Icff8af1f5c3ae89ef95ed8451273154b['h0000b] ;
//end
//always_comb begin
              If9057226a42b596a6dd2c84a37efff79['h00006] = 
          (!fgallag_sel['h00009]) ? 
                       Icff8af1f5c3ae89ef95ed8451273154b['h0000c] : //%
                       Icff8af1f5c3ae89ef95ed8451273154b['h0000d] ;
//end
//always_comb begin
              If9057226a42b596a6dd2c84a37efff79['h00007] = 
          (!fgallag_sel['h00009]) ? 
                       Icff8af1f5c3ae89ef95ed8451273154b['h0000e] : //%
                       Icff8af1f5c3ae89ef95ed8451273154b['h0000f] ;
//end
//always_comb begin
              If9057226a42b596a6dd2c84a37efff79['h00008] = 
          (!fgallag_sel['h00009]) ? 
                       Icff8af1f5c3ae89ef95ed8451273154b['h00010] : //%
                       Icff8af1f5c3ae89ef95ed8451273154b['h00011] ;
//end
//always_comb begin
              If9057226a42b596a6dd2c84a37efff79['h00009] = 
          (!fgallag_sel['h00009]) ? 
                       Icff8af1f5c3ae89ef95ed8451273154b['h00012] : //%
                       Icff8af1f5c3ae89ef95ed8451273154b['h00013] ;
//end
//always_comb begin
              If9057226a42b596a6dd2c84a37efff79['h0000a] = 
          (!fgallag_sel['h00009]) ? 
                       Icff8af1f5c3ae89ef95ed8451273154b['h00014] : //%
                       Icff8af1f5c3ae89ef95ed8451273154b['h00015] ;
//end
//always_comb begin
              If9057226a42b596a6dd2c84a37efff79['h0000b] = 
          (!fgallag_sel['h00009]) ? 
                       Icff8af1f5c3ae89ef95ed8451273154b['h00016] : //%
                       Icff8af1f5c3ae89ef95ed8451273154b['h00017] ;
//end
//always_comb begin
              If9057226a42b596a6dd2c84a37efff79['h0000c] = 
          (!fgallag_sel['h00009]) ? 
                       Icff8af1f5c3ae89ef95ed8451273154b['h00018] : //%
                       Icff8af1f5c3ae89ef95ed8451273154b['h00019] ;
//end
//always_comb begin
              If9057226a42b596a6dd2c84a37efff79['h0000d] = 
          (!fgallag_sel['h00009]) ? 
                       Icff8af1f5c3ae89ef95ed8451273154b['h0001a] : //%
                       Icff8af1f5c3ae89ef95ed8451273154b['h0001b] ;
//end
//always_comb begin
              If9057226a42b596a6dd2c84a37efff79['h0000e] = 
          (!fgallag_sel['h00009]) ? 
                       Icff8af1f5c3ae89ef95ed8451273154b['h0001c] : //%
                       Icff8af1f5c3ae89ef95ed8451273154b['h0001d] ;
//end
//always_comb begin
              If9057226a42b596a6dd2c84a37efff79['h0000f] = 
          (!fgallag_sel['h00009]) ? 
                       Icff8af1f5c3ae89ef95ed8451273154b['h0001e] : //%
                       Icff8af1f5c3ae89ef95ed8451273154b['h0001f] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00010] =  Icff8af1f5c3ae89ef95ed8451273154b['h00020] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00011] =  Icff8af1f5c3ae89ef95ed8451273154b['h00022] ;
//end
//always_comb begin
              If9057226a42b596a6dd2c84a37efff79['h00012] = 
          (!fgallag_sel['h00009]) ? 
                       Icff8af1f5c3ae89ef95ed8451273154b['h00024] : //%
                       Icff8af1f5c3ae89ef95ed8451273154b['h00025] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00013] =  Icff8af1f5c3ae89ef95ed8451273154b['h00026] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00014] =  Icff8af1f5c3ae89ef95ed8451273154b['h00028] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00015] =  Icff8af1f5c3ae89ef95ed8451273154b['h0002a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00016] =  Icff8af1f5c3ae89ef95ed8451273154b['h0002c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00017] =  Icff8af1f5c3ae89ef95ed8451273154b['h0002e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00018] =  Icff8af1f5c3ae89ef95ed8451273154b['h00030] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00019] =  Icff8af1f5c3ae89ef95ed8451273154b['h00032] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0001a] =  Icff8af1f5c3ae89ef95ed8451273154b['h00034] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0001b] =  Icff8af1f5c3ae89ef95ed8451273154b['h00036] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0001c] =  Icff8af1f5c3ae89ef95ed8451273154b['h00038] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0001d] =  Icff8af1f5c3ae89ef95ed8451273154b['h0003a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0001e] =  Icff8af1f5c3ae89ef95ed8451273154b['h0003c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0001f] =  Icff8af1f5c3ae89ef95ed8451273154b['h0003e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00020] =  Icff8af1f5c3ae89ef95ed8451273154b['h00040] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00021] =  Icff8af1f5c3ae89ef95ed8451273154b['h00042] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00022] =  Icff8af1f5c3ae89ef95ed8451273154b['h00044] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00023] =  Icff8af1f5c3ae89ef95ed8451273154b['h00046] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00024] =  Icff8af1f5c3ae89ef95ed8451273154b['h00048] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00025] =  Icff8af1f5c3ae89ef95ed8451273154b['h0004a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00026] =  Icff8af1f5c3ae89ef95ed8451273154b['h0004c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00027] =  Icff8af1f5c3ae89ef95ed8451273154b['h0004e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00028] =  Icff8af1f5c3ae89ef95ed8451273154b['h00050] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00029] =  Icff8af1f5c3ae89ef95ed8451273154b['h00052] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0002a] =  Icff8af1f5c3ae89ef95ed8451273154b['h00054] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0002b] =  Icff8af1f5c3ae89ef95ed8451273154b['h00056] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0002c] =  Icff8af1f5c3ae89ef95ed8451273154b['h00058] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0002d] =  Icff8af1f5c3ae89ef95ed8451273154b['h0005a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0002e] =  Icff8af1f5c3ae89ef95ed8451273154b['h0005c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0002f] =  Icff8af1f5c3ae89ef95ed8451273154b['h0005e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00030] =  Icff8af1f5c3ae89ef95ed8451273154b['h00060] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00031] =  Icff8af1f5c3ae89ef95ed8451273154b['h00062] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00032] =  Icff8af1f5c3ae89ef95ed8451273154b['h00064] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00033] =  Icff8af1f5c3ae89ef95ed8451273154b['h00066] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00034] =  Icff8af1f5c3ae89ef95ed8451273154b['h00068] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00035] =  Icff8af1f5c3ae89ef95ed8451273154b['h0006a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00036] =  Icff8af1f5c3ae89ef95ed8451273154b['h0006c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00037] =  Icff8af1f5c3ae89ef95ed8451273154b['h0006e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00038] =  Icff8af1f5c3ae89ef95ed8451273154b['h00070] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00039] =  Icff8af1f5c3ae89ef95ed8451273154b['h00072] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0003a] =  Icff8af1f5c3ae89ef95ed8451273154b['h00074] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0003b] =  Icff8af1f5c3ae89ef95ed8451273154b['h00076] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0003c] =  Icff8af1f5c3ae89ef95ed8451273154b['h00078] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0003d] =  Icff8af1f5c3ae89ef95ed8451273154b['h0007a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0003e] =  Icff8af1f5c3ae89ef95ed8451273154b['h0007c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0003f] =  Icff8af1f5c3ae89ef95ed8451273154b['h0007e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00040] =  Icff8af1f5c3ae89ef95ed8451273154b['h00080] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00041] =  Icff8af1f5c3ae89ef95ed8451273154b['h00082] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00042] =  Icff8af1f5c3ae89ef95ed8451273154b['h00084] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00043] =  Icff8af1f5c3ae89ef95ed8451273154b['h00086] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00044] =  Icff8af1f5c3ae89ef95ed8451273154b['h00088] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00045] =  Icff8af1f5c3ae89ef95ed8451273154b['h0008a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00046] =  Icff8af1f5c3ae89ef95ed8451273154b['h0008c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00047] =  Icff8af1f5c3ae89ef95ed8451273154b['h0008e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00048] =  Icff8af1f5c3ae89ef95ed8451273154b['h00090] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00049] =  Icff8af1f5c3ae89ef95ed8451273154b['h00092] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0004a] =  Icff8af1f5c3ae89ef95ed8451273154b['h00094] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0004b] =  Icff8af1f5c3ae89ef95ed8451273154b['h00096] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0004c] =  Icff8af1f5c3ae89ef95ed8451273154b['h00098] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0004d] =  Icff8af1f5c3ae89ef95ed8451273154b['h0009a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0004e] =  Icff8af1f5c3ae89ef95ed8451273154b['h0009c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0004f] =  Icff8af1f5c3ae89ef95ed8451273154b['h0009e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00050] =  Icff8af1f5c3ae89ef95ed8451273154b['h000a0] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00051] =  Icff8af1f5c3ae89ef95ed8451273154b['h000a2] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00052] =  Icff8af1f5c3ae89ef95ed8451273154b['h000a4] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00053] =  Icff8af1f5c3ae89ef95ed8451273154b['h000a6] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00054] =  Icff8af1f5c3ae89ef95ed8451273154b['h000a8] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00055] =  Icff8af1f5c3ae89ef95ed8451273154b['h000aa] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00056] =  Icff8af1f5c3ae89ef95ed8451273154b['h000ac] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00057] =  Icff8af1f5c3ae89ef95ed8451273154b['h000ae] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00058] =  Icff8af1f5c3ae89ef95ed8451273154b['h000b0] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00059] =  Icff8af1f5c3ae89ef95ed8451273154b['h000b2] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0005a] =  Icff8af1f5c3ae89ef95ed8451273154b['h000b4] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0005b] =  Icff8af1f5c3ae89ef95ed8451273154b['h000b6] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0005c] =  Icff8af1f5c3ae89ef95ed8451273154b['h000b8] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0005d] =  Icff8af1f5c3ae89ef95ed8451273154b['h000ba] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0005e] =  Icff8af1f5c3ae89ef95ed8451273154b['h000bc] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0005f] =  Icff8af1f5c3ae89ef95ed8451273154b['h000be] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00060] =  Icff8af1f5c3ae89ef95ed8451273154b['h000c0] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00061] =  Icff8af1f5c3ae89ef95ed8451273154b['h000c2] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00062] =  Icff8af1f5c3ae89ef95ed8451273154b['h000c4] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00063] =  Icff8af1f5c3ae89ef95ed8451273154b['h000c6] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00064] =  Icff8af1f5c3ae89ef95ed8451273154b['h000c8] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00065] =  Icff8af1f5c3ae89ef95ed8451273154b['h000ca] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00066] =  Icff8af1f5c3ae89ef95ed8451273154b['h000cc] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00067] =  Icff8af1f5c3ae89ef95ed8451273154b['h000ce] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00068] =  Icff8af1f5c3ae89ef95ed8451273154b['h000d0] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00069] =  Icff8af1f5c3ae89ef95ed8451273154b['h000d2] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0006a] =  Icff8af1f5c3ae89ef95ed8451273154b['h000d4] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0006b] =  Icff8af1f5c3ae89ef95ed8451273154b['h000d6] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0006c] =  Icff8af1f5c3ae89ef95ed8451273154b['h000d8] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0006d] =  Icff8af1f5c3ae89ef95ed8451273154b['h000da] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0006e] =  Icff8af1f5c3ae89ef95ed8451273154b['h000dc] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0006f] =  Icff8af1f5c3ae89ef95ed8451273154b['h000de] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00070] =  Icff8af1f5c3ae89ef95ed8451273154b['h000e0] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00071] =  Icff8af1f5c3ae89ef95ed8451273154b['h000e2] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00072] =  Icff8af1f5c3ae89ef95ed8451273154b['h000e4] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00073] =  Icff8af1f5c3ae89ef95ed8451273154b['h000e6] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00074] =  Icff8af1f5c3ae89ef95ed8451273154b['h000e8] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00075] =  Icff8af1f5c3ae89ef95ed8451273154b['h000ea] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00076] =  Icff8af1f5c3ae89ef95ed8451273154b['h000ec] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00077] =  Icff8af1f5c3ae89ef95ed8451273154b['h000ee] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00078] =  Icff8af1f5c3ae89ef95ed8451273154b['h000f0] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00079] =  Icff8af1f5c3ae89ef95ed8451273154b['h000f2] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0007a] =  Icff8af1f5c3ae89ef95ed8451273154b['h000f4] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0007b] =  Icff8af1f5c3ae89ef95ed8451273154b['h000f6] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0007c] =  Icff8af1f5c3ae89ef95ed8451273154b['h000f8] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0007d] =  Icff8af1f5c3ae89ef95ed8451273154b['h000fa] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0007e] =  Icff8af1f5c3ae89ef95ed8451273154b['h000fc] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0007f] =  Icff8af1f5c3ae89ef95ed8451273154b['h000fe] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00080] =  Icff8af1f5c3ae89ef95ed8451273154b['h00100] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00081] =  Icff8af1f5c3ae89ef95ed8451273154b['h00102] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00082] =  Icff8af1f5c3ae89ef95ed8451273154b['h00104] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00083] =  Icff8af1f5c3ae89ef95ed8451273154b['h00106] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00084] =  Icff8af1f5c3ae89ef95ed8451273154b['h00108] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00085] =  Icff8af1f5c3ae89ef95ed8451273154b['h0010a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00086] =  Icff8af1f5c3ae89ef95ed8451273154b['h0010c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00087] =  Icff8af1f5c3ae89ef95ed8451273154b['h0010e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00088] =  Icff8af1f5c3ae89ef95ed8451273154b['h00110] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00089] =  Icff8af1f5c3ae89ef95ed8451273154b['h00112] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0008a] =  Icff8af1f5c3ae89ef95ed8451273154b['h00114] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0008b] =  Icff8af1f5c3ae89ef95ed8451273154b['h00116] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0008c] =  Icff8af1f5c3ae89ef95ed8451273154b['h00118] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0008d] =  Icff8af1f5c3ae89ef95ed8451273154b['h0011a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0008e] =  Icff8af1f5c3ae89ef95ed8451273154b['h0011c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0008f] =  Icff8af1f5c3ae89ef95ed8451273154b['h0011e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00090] =  Icff8af1f5c3ae89ef95ed8451273154b['h00120] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00091] =  Icff8af1f5c3ae89ef95ed8451273154b['h00122] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00092] =  Icff8af1f5c3ae89ef95ed8451273154b['h00124] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00093] =  Icff8af1f5c3ae89ef95ed8451273154b['h00126] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00094] =  Icff8af1f5c3ae89ef95ed8451273154b['h00128] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00095] =  Icff8af1f5c3ae89ef95ed8451273154b['h0012a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00096] =  Icff8af1f5c3ae89ef95ed8451273154b['h0012c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00097] =  Icff8af1f5c3ae89ef95ed8451273154b['h0012e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00098] =  Icff8af1f5c3ae89ef95ed8451273154b['h00130] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00099] =  Icff8af1f5c3ae89ef95ed8451273154b['h00132] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0009a] =  Icff8af1f5c3ae89ef95ed8451273154b['h00134] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0009b] =  Icff8af1f5c3ae89ef95ed8451273154b['h00136] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0009c] =  Icff8af1f5c3ae89ef95ed8451273154b['h00138] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0009d] =  Icff8af1f5c3ae89ef95ed8451273154b['h0013a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0009e] =  Icff8af1f5c3ae89ef95ed8451273154b['h0013c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0009f] =  Icff8af1f5c3ae89ef95ed8451273154b['h0013e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000a0] =  Icff8af1f5c3ae89ef95ed8451273154b['h00140] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000a1] =  Icff8af1f5c3ae89ef95ed8451273154b['h00142] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000a2] =  Icff8af1f5c3ae89ef95ed8451273154b['h00144] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000a3] =  Icff8af1f5c3ae89ef95ed8451273154b['h00146] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000a4] =  Icff8af1f5c3ae89ef95ed8451273154b['h00148] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000a5] =  Icff8af1f5c3ae89ef95ed8451273154b['h0014a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000a6] =  Icff8af1f5c3ae89ef95ed8451273154b['h0014c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000a7] =  Icff8af1f5c3ae89ef95ed8451273154b['h0014e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000a8] =  Icff8af1f5c3ae89ef95ed8451273154b['h00150] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000a9] =  Icff8af1f5c3ae89ef95ed8451273154b['h00152] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000aa] =  Icff8af1f5c3ae89ef95ed8451273154b['h00154] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000ab] =  Icff8af1f5c3ae89ef95ed8451273154b['h00156] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000ac] =  Icff8af1f5c3ae89ef95ed8451273154b['h00158] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000ad] =  Icff8af1f5c3ae89ef95ed8451273154b['h0015a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000ae] =  Icff8af1f5c3ae89ef95ed8451273154b['h0015c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000af] =  Icff8af1f5c3ae89ef95ed8451273154b['h0015e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000b0] =  Icff8af1f5c3ae89ef95ed8451273154b['h00160] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000b1] =  Icff8af1f5c3ae89ef95ed8451273154b['h00162] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000b2] =  Icff8af1f5c3ae89ef95ed8451273154b['h00164] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000b3] =  Icff8af1f5c3ae89ef95ed8451273154b['h00166] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000b4] =  Icff8af1f5c3ae89ef95ed8451273154b['h00168] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000b5] =  Icff8af1f5c3ae89ef95ed8451273154b['h0016a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000b6] =  Icff8af1f5c3ae89ef95ed8451273154b['h0016c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000b7] =  Icff8af1f5c3ae89ef95ed8451273154b['h0016e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000b8] =  Icff8af1f5c3ae89ef95ed8451273154b['h00170] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000b9] =  Icff8af1f5c3ae89ef95ed8451273154b['h00172] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000ba] =  Icff8af1f5c3ae89ef95ed8451273154b['h00174] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000bb] =  Icff8af1f5c3ae89ef95ed8451273154b['h00176] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000bc] =  Icff8af1f5c3ae89ef95ed8451273154b['h00178] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000bd] =  Icff8af1f5c3ae89ef95ed8451273154b['h0017a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000be] =  Icff8af1f5c3ae89ef95ed8451273154b['h0017c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000bf] =  Icff8af1f5c3ae89ef95ed8451273154b['h0017e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000c0] =  Icff8af1f5c3ae89ef95ed8451273154b['h00180] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000c1] =  Icff8af1f5c3ae89ef95ed8451273154b['h00182] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000c2] =  Icff8af1f5c3ae89ef95ed8451273154b['h00184] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000c3] =  Icff8af1f5c3ae89ef95ed8451273154b['h00186] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000c4] =  Icff8af1f5c3ae89ef95ed8451273154b['h00188] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000c5] =  Icff8af1f5c3ae89ef95ed8451273154b['h0018a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000c6] =  Icff8af1f5c3ae89ef95ed8451273154b['h0018c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000c7] =  Icff8af1f5c3ae89ef95ed8451273154b['h0018e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000c8] =  Icff8af1f5c3ae89ef95ed8451273154b['h00190] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000c9] =  Icff8af1f5c3ae89ef95ed8451273154b['h00192] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000ca] =  Icff8af1f5c3ae89ef95ed8451273154b['h00194] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000cb] =  Icff8af1f5c3ae89ef95ed8451273154b['h00196] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000cc] =  Icff8af1f5c3ae89ef95ed8451273154b['h00198] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000cd] =  Icff8af1f5c3ae89ef95ed8451273154b['h0019a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000ce] =  Icff8af1f5c3ae89ef95ed8451273154b['h0019c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000cf] =  Icff8af1f5c3ae89ef95ed8451273154b['h0019e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000d0] =  Icff8af1f5c3ae89ef95ed8451273154b['h001a0] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000d1] =  Icff8af1f5c3ae89ef95ed8451273154b['h001a2] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000d2] =  Icff8af1f5c3ae89ef95ed8451273154b['h001a4] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000d3] =  Icff8af1f5c3ae89ef95ed8451273154b['h001a6] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000d4] =  Icff8af1f5c3ae89ef95ed8451273154b['h001a8] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000d5] =  Icff8af1f5c3ae89ef95ed8451273154b['h001aa] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000d6] =  Icff8af1f5c3ae89ef95ed8451273154b['h001ac] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000d7] =  Icff8af1f5c3ae89ef95ed8451273154b['h001ae] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000d8] =  Icff8af1f5c3ae89ef95ed8451273154b['h001b0] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000d9] =  Icff8af1f5c3ae89ef95ed8451273154b['h001b2] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000da] =  Icff8af1f5c3ae89ef95ed8451273154b['h001b4] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000db] =  Icff8af1f5c3ae89ef95ed8451273154b['h001b6] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000dc] =  Icff8af1f5c3ae89ef95ed8451273154b['h001b8] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000dd] =  Icff8af1f5c3ae89ef95ed8451273154b['h001ba] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000de] =  Icff8af1f5c3ae89ef95ed8451273154b['h001bc] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000df] =  Icff8af1f5c3ae89ef95ed8451273154b['h001be] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000e0] =  Icff8af1f5c3ae89ef95ed8451273154b['h001c0] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000e1] =  Icff8af1f5c3ae89ef95ed8451273154b['h001c2] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000e2] =  Icff8af1f5c3ae89ef95ed8451273154b['h001c4] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000e3] =  Icff8af1f5c3ae89ef95ed8451273154b['h001c6] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000e4] =  Icff8af1f5c3ae89ef95ed8451273154b['h001c8] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000e5] =  Icff8af1f5c3ae89ef95ed8451273154b['h001ca] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000e6] =  Icff8af1f5c3ae89ef95ed8451273154b['h001cc] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000e7] =  Icff8af1f5c3ae89ef95ed8451273154b['h001ce] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000e8] =  Icff8af1f5c3ae89ef95ed8451273154b['h001d0] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000e9] =  Icff8af1f5c3ae89ef95ed8451273154b['h001d2] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000ea] =  Icff8af1f5c3ae89ef95ed8451273154b['h001d4] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000eb] =  Icff8af1f5c3ae89ef95ed8451273154b['h001d6] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000ec] =  Icff8af1f5c3ae89ef95ed8451273154b['h001d8] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000ed] =  Icff8af1f5c3ae89ef95ed8451273154b['h001da] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000ee] =  Icff8af1f5c3ae89ef95ed8451273154b['h001dc] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000ef] =  Icff8af1f5c3ae89ef95ed8451273154b['h001de] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000f0] =  Icff8af1f5c3ae89ef95ed8451273154b['h001e0] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000f1] =  Icff8af1f5c3ae89ef95ed8451273154b['h001e2] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000f2] =  Icff8af1f5c3ae89ef95ed8451273154b['h001e4] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000f3] =  Icff8af1f5c3ae89ef95ed8451273154b['h001e6] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000f4] =  Icff8af1f5c3ae89ef95ed8451273154b['h001e8] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000f5] =  Icff8af1f5c3ae89ef95ed8451273154b['h001ea] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000f6] =  Icff8af1f5c3ae89ef95ed8451273154b['h001ec] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000f7] =  Icff8af1f5c3ae89ef95ed8451273154b['h001ee] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000f8] =  Icff8af1f5c3ae89ef95ed8451273154b['h001f0] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000f9] =  Icff8af1f5c3ae89ef95ed8451273154b['h001f2] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000fa] =  Icff8af1f5c3ae89ef95ed8451273154b['h001f4] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000fb] =  Icff8af1f5c3ae89ef95ed8451273154b['h001f6] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000fc] =  Icff8af1f5c3ae89ef95ed8451273154b['h001f8] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000fd] =  Icff8af1f5c3ae89ef95ed8451273154b['h001fa] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000fe] =  Icff8af1f5c3ae89ef95ed8451273154b['h001fc] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h000ff] =  Icff8af1f5c3ae89ef95ed8451273154b['h001fe] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00100] =  Icff8af1f5c3ae89ef95ed8451273154b['h00200] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00101] =  Icff8af1f5c3ae89ef95ed8451273154b['h00202] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00102] =  Icff8af1f5c3ae89ef95ed8451273154b['h00204] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00103] =  Icff8af1f5c3ae89ef95ed8451273154b['h00206] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00104] =  Icff8af1f5c3ae89ef95ed8451273154b['h00208] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00105] =  Icff8af1f5c3ae89ef95ed8451273154b['h0020a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00106] =  Icff8af1f5c3ae89ef95ed8451273154b['h0020c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00107] =  Icff8af1f5c3ae89ef95ed8451273154b['h0020e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00108] =  Icff8af1f5c3ae89ef95ed8451273154b['h00210] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00109] =  Icff8af1f5c3ae89ef95ed8451273154b['h00212] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0010a] =  Icff8af1f5c3ae89ef95ed8451273154b['h00214] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0010b] =  Icff8af1f5c3ae89ef95ed8451273154b['h00216] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0010c] =  Icff8af1f5c3ae89ef95ed8451273154b['h00218] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0010d] =  Icff8af1f5c3ae89ef95ed8451273154b['h0021a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0010e] =  Icff8af1f5c3ae89ef95ed8451273154b['h0021c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0010f] =  Icff8af1f5c3ae89ef95ed8451273154b['h0021e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00110] =  Icff8af1f5c3ae89ef95ed8451273154b['h00220] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00111] =  Icff8af1f5c3ae89ef95ed8451273154b['h00222] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00112] =  Icff8af1f5c3ae89ef95ed8451273154b['h00224] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00113] =  Icff8af1f5c3ae89ef95ed8451273154b['h00226] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00114] =  Icff8af1f5c3ae89ef95ed8451273154b['h00228] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00115] =  Icff8af1f5c3ae89ef95ed8451273154b['h0022a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00116] =  Icff8af1f5c3ae89ef95ed8451273154b['h0022c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00117] =  Icff8af1f5c3ae89ef95ed8451273154b['h0022e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00118] =  Icff8af1f5c3ae89ef95ed8451273154b['h00230] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00119] =  Icff8af1f5c3ae89ef95ed8451273154b['h00232] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0011a] =  Icff8af1f5c3ae89ef95ed8451273154b['h00234] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0011b] =  Icff8af1f5c3ae89ef95ed8451273154b['h00236] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0011c] =  Icff8af1f5c3ae89ef95ed8451273154b['h00238] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0011d] =  Icff8af1f5c3ae89ef95ed8451273154b['h0023a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0011e] =  Icff8af1f5c3ae89ef95ed8451273154b['h0023c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0011f] =  Icff8af1f5c3ae89ef95ed8451273154b['h0023e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00120] =  Icff8af1f5c3ae89ef95ed8451273154b['h00240] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00121] =  Icff8af1f5c3ae89ef95ed8451273154b['h00242] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00122] =  Icff8af1f5c3ae89ef95ed8451273154b['h00244] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00123] =  Icff8af1f5c3ae89ef95ed8451273154b['h00246] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00124] =  Icff8af1f5c3ae89ef95ed8451273154b['h00248] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00125] =  Icff8af1f5c3ae89ef95ed8451273154b['h0024a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00126] =  Icff8af1f5c3ae89ef95ed8451273154b['h0024c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00127] =  Icff8af1f5c3ae89ef95ed8451273154b['h0024e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00128] =  Icff8af1f5c3ae89ef95ed8451273154b['h00250] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00129] =  Icff8af1f5c3ae89ef95ed8451273154b['h00252] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0012a] =  Icff8af1f5c3ae89ef95ed8451273154b['h00254] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0012b] =  Icff8af1f5c3ae89ef95ed8451273154b['h00256] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0012c] =  Icff8af1f5c3ae89ef95ed8451273154b['h00258] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0012d] =  Icff8af1f5c3ae89ef95ed8451273154b['h0025a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0012e] =  Icff8af1f5c3ae89ef95ed8451273154b['h0025c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0012f] =  Icff8af1f5c3ae89ef95ed8451273154b['h0025e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00130] =  Icff8af1f5c3ae89ef95ed8451273154b['h00260] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00131] =  Icff8af1f5c3ae89ef95ed8451273154b['h00262] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00132] =  Icff8af1f5c3ae89ef95ed8451273154b['h00264] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00133] =  Icff8af1f5c3ae89ef95ed8451273154b['h00266] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00134] =  Icff8af1f5c3ae89ef95ed8451273154b['h00268] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00135] =  Icff8af1f5c3ae89ef95ed8451273154b['h0026a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00136] =  Icff8af1f5c3ae89ef95ed8451273154b['h0026c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00137] =  Icff8af1f5c3ae89ef95ed8451273154b['h0026e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00138] =  Icff8af1f5c3ae89ef95ed8451273154b['h00270] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00139] =  Icff8af1f5c3ae89ef95ed8451273154b['h00272] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0013a] =  Icff8af1f5c3ae89ef95ed8451273154b['h00274] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0013b] =  Icff8af1f5c3ae89ef95ed8451273154b['h00276] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0013c] =  Icff8af1f5c3ae89ef95ed8451273154b['h00278] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0013d] =  Icff8af1f5c3ae89ef95ed8451273154b['h0027a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0013e] =  Icff8af1f5c3ae89ef95ed8451273154b['h0027c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0013f] =  Icff8af1f5c3ae89ef95ed8451273154b['h0027e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00140] =  Icff8af1f5c3ae89ef95ed8451273154b['h00280] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00141] =  Icff8af1f5c3ae89ef95ed8451273154b['h00282] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00142] =  Icff8af1f5c3ae89ef95ed8451273154b['h00284] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00143] =  Icff8af1f5c3ae89ef95ed8451273154b['h00286] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00144] =  Icff8af1f5c3ae89ef95ed8451273154b['h00288] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00145] =  Icff8af1f5c3ae89ef95ed8451273154b['h0028a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00146] =  Icff8af1f5c3ae89ef95ed8451273154b['h0028c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00147] =  Icff8af1f5c3ae89ef95ed8451273154b['h0028e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00148] =  Icff8af1f5c3ae89ef95ed8451273154b['h00290] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00149] =  Icff8af1f5c3ae89ef95ed8451273154b['h00292] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0014a] =  Icff8af1f5c3ae89ef95ed8451273154b['h00294] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0014b] =  Icff8af1f5c3ae89ef95ed8451273154b['h00296] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0014c] =  Icff8af1f5c3ae89ef95ed8451273154b['h00298] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0014d] =  Icff8af1f5c3ae89ef95ed8451273154b['h0029a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0014e] =  Icff8af1f5c3ae89ef95ed8451273154b['h0029c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0014f] =  Icff8af1f5c3ae89ef95ed8451273154b['h0029e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00150] =  Icff8af1f5c3ae89ef95ed8451273154b['h002a0] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00151] =  Icff8af1f5c3ae89ef95ed8451273154b['h002a2] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00152] =  Icff8af1f5c3ae89ef95ed8451273154b['h002a4] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00153] =  Icff8af1f5c3ae89ef95ed8451273154b['h002a6] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00154] =  Icff8af1f5c3ae89ef95ed8451273154b['h002a8] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00155] =  Icff8af1f5c3ae89ef95ed8451273154b['h002aa] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00156] =  Icff8af1f5c3ae89ef95ed8451273154b['h002ac] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00157] =  Icff8af1f5c3ae89ef95ed8451273154b['h002ae] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00158] =  Icff8af1f5c3ae89ef95ed8451273154b['h002b0] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00159] =  Icff8af1f5c3ae89ef95ed8451273154b['h002b2] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0015a] =  Icff8af1f5c3ae89ef95ed8451273154b['h002b4] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0015b] =  Icff8af1f5c3ae89ef95ed8451273154b['h002b6] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0015c] =  Icff8af1f5c3ae89ef95ed8451273154b['h002b8] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0015d] =  Icff8af1f5c3ae89ef95ed8451273154b['h002ba] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0015e] =  Icff8af1f5c3ae89ef95ed8451273154b['h002bc] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0015f] =  Icff8af1f5c3ae89ef95ed8451273154b['h002be] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00160] =  Icff8af1f5c3ae89ef95ed8451273154b['h002c0] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00161] =  Icff8af1f5c3ae89ef95ed8451273154b['h002c2] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00162] =  Icff8af1f5c3ae89ef95ed8451273154b['h002c4] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00163] =  Icff8af1f5c3ae89ef95ed8451273154b['h002c6] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00164] =  Icff8af1f5c3ae89ef95ed8451273154b['h002c8] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00165] =  Icff8af1f5c3ae89ef95ed8451273154b['h002ca] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00166] =  Icff8af1f5c3ae89ef95ed8451273154b['h002cc] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00167] =  Icff8af1f5c3ae89ef95ed8451273154b['h002ce] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00168] =  Icff8af1f5c3ae89ef95ed8451273154b['h002d0] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00169] =  Icff8af1f5c3ae89ef95ed8451273154b['h002d2] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0016a] =  Icff8af1f5c3ae89ef95ed8451273154b['h002d4] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0016b] =  Icff8af1f5c3ae89ef95ed8451273154b['h002d6] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0016c] =  Icff8af1f5c3ae89ef95ed8451273154b['h002d8] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0016d] =  Icff8af1f5c3ae89ef95ed8451273154b['h002da] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0016e] =  Icff8af1f5c3ae89ef95ed8451273154b['h002dc] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0016f] =  Icff8af1f5c3ae89ef95ed8451273154b['h002de] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00170] =  Icff8af1f5c3ae89ef95ed8451273154b['h002e0] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00171] =  Icff8af1f5c3ae89ef95ed8451273154b['h002e2] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00172] =  Icff8af1f5c3ae89ef95ed8451273154b['h002e4] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00173] =  Icff8af1f5c3ae89ef95ed8451273154b['h002e6] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00174] =  Icff8af1f5c3ae89ef95ed8451273154b['h002e8] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00175] =  Icff8af1f5c3ae89ef95ed8451273154b['h002ea] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00176] =  Icff8af1f5c3ae89ef95ed8451273154b['h002ec] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00177] =  Icff8af1f5c3ae89ef95ed8451273154b['h002ee] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00178] =  Icff8af1f5c3ae89ef95ed8451273154b['h002f0] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00179] =  Icff8af1f5c3ae89ef95ed8451273154b['h002f2] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0017a] =  Icff8af1f5c3ae89ef95ed8451273154b['h002f4] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0017b] =  Icff8af1f5c3ae89ef95ed8451273154b['h002f6] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0017c] =  Icff8af1f5c3ae89ef95ed8451273154b['h002f8] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0017d] =  Icff8af1f5c3ae89ef95ed8451273154b['h002fa] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0017e] =  Icff8af1f5c3ae89ef95ed8451273154b['h002fc] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0017f] =  Icff8af1f5c3ae89ef95ed8451273154b['h002fe] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00180] =  Icff8af1f5c3ae89ef95ed8451273154b['h00300] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00181] =  Icff8af1f5c3ae89ef95ed8451273154b['h00302] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00182] =  Icff8af1f5c3ae89ef95ed8451273154b['h00304] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00183] =  Icff8af1f5c3ae89ef95ed8451273154b['h00306] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00184] =  Icff8af1f5c3ae89ef95ed8451273154b['h00308] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00185] =  Icff8af1f5c3ae89ef95ed8451273154b['h0030a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00186] =  Icff8af1f5c3ae89ef95ed8451273154b['h0030c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00187] =  Icff8af1f5c3ae89ef95ed8451273154b['h0030e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00188] =  Icff8af1f5c3ae89ef95ed8451273154b['h00310] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00189] =  Icff8af1f5c3ae89ef95ed8451273154b['h00312] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0018a] =  Icff8af1f5c3ae89ef95ed8451273154b['h00314] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0018b] =  Icff8af1f5c3ae89ef95ed8451273154b['h00316] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0018c] =  Icff8af1f5c3ae89ef95ed8451273154b['h00318] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0018d] =  Icff8af1f5c3ae89ef95ed8451273154b['h0031a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0018e] =  Icff8af1f5c3ae89ef95ed8451273154b['h0031c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0018f] =  Icff8af1f5c3ae89ef95ed8451273154b['h0031e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00190] =  Icff8af1f5c3ae89ef95ed8451273154b['h00320] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00191] =  Icff8af1f5c3ae89ef95ed8451273154b['h00322] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00192] =  Icff8af1f5c3ae89ef95ed8451273154b['h00324] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00193] =  Icff8af1f5c3ae89ef95ed8451273154b['h00326] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00194] =  Icff8af1f5c3ae89ef95ed8451273154b['h00328] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00195] =  Icff8af1f5c3ae89ef95ed8451273154b['h0032a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00196] =  Icff8af1f5c3ae89ef95ed8451273154b['h0032c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00197] =  Icff8af1f5c3ae89ef95ed8451273154b['h0032e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00198] =  Icff8af1f5c3ae89ef95ed8451273154b['h00330] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h00199] =  Icff8af1f5c3ae89ef95ed8451273154b['h00332] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0019a] =  Icff8af1f5c3ae89ef95ed8451273154b['h00334] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0019b] =  Icff8af1f5c3ae89ef95ed8451273154b['h00336] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0019c] =  Icff8af1f5c3ae89ef95ed8451273154b['h00338] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0019d] =  Icff8af1f5c3ae89ef95ed8451273154b['h0033a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0019e] =  Icff8af1f5c3ae89ef95ed8451273154b['h0033c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h0019f] =  Icff8af1f5c3ae89ef95ed8451273154b['h0033e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001a0] =  Icff8af1f5c3ae89ef95ed8451273154b['h00340] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001a1] =  Icff8af1f5c3ae89ef95ed8451273154b['h00342] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001a2] =  Icff8af1f5c3ae89ef95ed8451273154b['h00344] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001a3] =  Icff8af1f5c3ae89ef95ed8451273154b['h00346] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001a4] =  Icff8af1f5c3ae89ef95ed8451273154b['h00348] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001a5] =  Icff8af1f5c3ae89ef95ed8451273154b['h0034a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001a6] =  Icff8af1f5c3ae89ef95ed8451273154b['h0034c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001a7] =  Icff8af1f5c3ae89ef95ed8451273154b['h0034e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001a8] =  Icff8af1f5c3ae89ef95ed8451273154b['h00350] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001a9] =  Icff8af1f5c3ae89ef95ed8451273154b['h00352] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001aa] =  Icff8af1f5c3ae89ef95ed8451273154b['h00354] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001ab] =  Icff8af1f5c3ae89ef95ed8451273154b['h00356] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001ac] =  Icff8af1f5c3ae89ef95ed8451273154b['h00358] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001ad] =  Icff8af1f5c3ae89ef95ed8451273154b['h0035a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001ae] =  Icff8af1f5c3ae89ef95ed8451273154b['h0035c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001af] =  Icff8af1f5c3ae89ef95ed8451273154b['h0035e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001b0] =  Icff8af1f5c3ae89ef95ed8451273154b['h00360] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001b1] =  Icff8af1f5c3ae89ef95ed8451273154b['h00362] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001b2] =  Icff8af1f5c3ae89ef95ed8451273154b['h00364] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001b3] =  Icff8af1f5c3ae89ef95ed8451273154b['h00366] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001b4] =  Icff8af1f5c3ae89ef95ed8451273154b['h00368] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001b5] =  Icff8af1f5c3ae89ef95ed8451273154b['h0036a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001b6] =  Icff8af1f5c3ae89ef95ed8451273154b['h0036c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001b7] =  Icff8af1f5c3ae89ef95ed8451273154b['h0036e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001b8] =  Icff8af1f5c3ae89ef95ed8451273154b['h00370] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001b9] =  Icff8af1f5c3ae89ef95ed8451273154b['h00372] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001ba] =  Icff8af1f5c3ae89ef95ed8451273154b['h00374] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001bb] =  Icff8af1f5c3ae89ef95ed8451273154b['h00376] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001bc] =  Icff8af1f5c3ae89ef95ed8451273154b['h00378] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001bd] =  Icff8af1f5c3ae89ef95ed8451273154b['h0037a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001be] =  Icff8af1f5c3ae89ef95ed8451273154b['h0037c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001bf] =  Icff8af1f5c3ae89ef95ed8451273154b['h0037e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001c0] =  Icff8af1f5c3ae89ef95ed8451273154b['h00380] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001c1] =  Icff8af1f5c3ae89ef95ed8451273154b['h00382] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001c2] =  Icff8af1f5c3ae89ef95ed8451273154b['h00384] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001c3] =  Icff8af1f5c3ae89ef95ed8451273154b['h00386] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001c4] =  Icff8af1f5c3ae89ef95ed8451273154b['h00388] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001c5] =  Icff8af1f5c3ae89ef95ed8451273154b['h0038a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001c6] =  Icff8af1f5c3ae89ef95ed8451273154b['h0038c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001c7] =  Icff8af1f5c3ae89ef95ed8451273154b['h0038e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001c8] =  Icff8af1f5c3ae89ef95ed8451273154b['h00390] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001c9] =  Icff8af1f5c3ae89ef95ed8451273154b['h00392] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001ca] =  Icff8af1f5c3ae89ef95ed8451273154b['h00394] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001cb] =  Icff8af1f5c3ae89ef95ed8451273154b['h00396] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001cc] =  Icff8af1f5c3ae89ef95ed8451273154b['h00398] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001cd] =  Icff8af1f5c3ae89ef95ed8451273154b['h0039a] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001ce] =  Icff8af1f5c3ae89ef95ed8451273154b['h0039c] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001cf] =  Icff8af1f5c3ae89ef95ed8451273154b['h0039e] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001d0] =  Icff8af1f5c3ae89ef95ed8451273154b['h003a0] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001d1] =  Icff8af1f5c3ae89ef95ed8451273154b['h003a2] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001d2] =  Icff8af1f5c3ae89ef95ed8451273154b['h003a4] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001d3] =  Icff8af1f5c3ae89ef95ed8451273154b['h003a6] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001d4] =  Icff8af1f5c3ae89ef95ed8451273154b['h003a8] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001d5] =  Icff8af1f5c3ae89ef95ed8451273154b['h003aa] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001d6] =  Icff8af1f5c3ae89ef95ed8451273154b['h003ac] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001d7] =  Icff8af1f5c3ae89ef95ed8451273154b['h003ae] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001d8] =  Icff8af1f5c3ae89ef95ed8451273154b['h003b0] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001d9] =  Icff8af1f5c3ae89ef95ed8451273154b['h003b2] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001da] =  Icff8af1f5c3ae89ef95ed8451273154b['h003b4] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001db] =  Icff8af1f5c3ae89ef95ed8451273154b['h003b6] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001dc] =  Icff8af1f5c3ae89ef95ed8451273154b['h003b8] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001dd] =  Icff8af1f5c3ae89ef95ed8451273154b['h003ba] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001de] =  Icff8af1f5c3ae89ef95ed8451273154b['h003bc] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001df] =  Icff8af1f5c3ae89ef95ed8451273154b['h003be] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001e0] =  Icff8af1f5c3ae89ef95ed8451273154b['h003c0] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001e1] =  Icff8af1f5c3ae89ef95ed8451273154b['h003c2] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001e2] =  Icff8af1f5c3ae89ef95ed8451273154b['h003c4] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001e3] =  Icff8af1f5c3ae89ef95ed8451273154b['h003c6] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001e4] =  Icff8af1f5c3ae89ef95ed8451273154b['h003c8] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001e5] =  Icff8af1f5c3ae89ef95ed8451273154b['h003ca] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001e6] =  Icff8af1f5c3ae89ef95ed8451273154b['h003cc] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001e7] =  Icff8af1f5c3ae89ef95ed8451273154b['h003ce] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001e8] =  Icff8af1f5c3ae89ef95ed8451273154b['h003d0] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001e9] =  Icff8af1f5c3ae89ef95ed8451273154b['h003d2] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001ea] =  Icff8af1f5c3ae89ef95ed8451273154b['h003d4] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001eb] =  Icff8af1f5c3ae89ef95ed8451273154b['h003d6] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001ec] =  Icff8af1f5c3ae89ef95ed8451273154b['h003d8] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001ed] =  Icff8af1f5c3ae89ef95ed8451273154b['h003da] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001ee] =  Icff8af1f5c3ae89ef95ed8451273154b['h003dc] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001ef] =  Icff8af1f5c3ae89ef95ed8451273154b['h003de] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001f0] =  Icff8af1f5c3ae89ef95ed8451273154b['h003e0] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001f1] =  Icff8af1f5c3ae89ef95ed8451273154b['h003e2] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001f2] =  Icff8af1f5c3ae89ef95ed8451273154b['h003e4] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001f3] =  Icff8af1f5c3ae89ef95ed8451273154b['h003e6] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001f4] =  Icff8af1f5c3ae89ef95ed8451273154b['h003e8] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001f5] =  Icff8af1f5c3ae89ef95ed8451273154b['h003ea] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001f6] =  Icff8af1f5c3ae89ef95ed8451273154b['h003ec] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001f7] =  Icff8af1f5c3ae89ef95ed8451273154b['h003ee] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001f8] =  Icff8af1f5c3ae89ef95ed8451273154b['h003f0] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001f9] =  Icff8af1f5c3ae89ef95ed8451273154b['h003f2] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001fa] =  Icff8af1f5c3ae89ef95ed8451273154b['h003f4] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001fb] =  Icff8af1f5c3ae89ef95ed8451273154b['h003f6] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001fc] =  Icff8af1f5c3ae89ef95ed8451273154b['h003f8] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001fd] =  Icff8af1f5c3ae89ef95ed8451273154b['h003fa] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001fe] =  Icff8af1f5c3ae89ef95ed8451273154b['h003fc] ;
//end
//always_comb begin // 
               If9057226a42b596a6dd2c84a37efff79['h001ff] =  Icff8af1f5c3ae89ef95ed8451273154b['h003fe] ;
//end
