//`include "GF2_LDPC_flogtanh_0x0000f_assign_inc.sv"
//always_comb begin
              Iae34f8e78093d5bcc3db929580c94da8015f69b8c6dd2133f36668c2d4b1e0c7['h00000] = 
          (!flogtanh_sel['h0000f]) ? 
                       Ica808b9c1910a49740bb889b7521538bc786bf51f6b2c7c3ad1af9712127147b['h00000] : //%
                       Ica808b9c1910a49740bb889b7521538bc786bf51f6b2c7c3ad1af9712127147b['h00001] ;
//end
//always_comb begin // 
               Iae34f8e78093d5bcc3db929580c94da8015f69b8c6dd2133f36668c2d4b1e0c7['h00001] =  Ica808b9c1910a49740bb889b7521538bc786bf51f6b2c7c3ad1af9712127147b['h00002] ;
//end
//always_comb begin // 
               Iae34f8e78093d5bcc3db929580c94da8015f69b8c6dd2133f36668c2d4b1e0c7['h00002] =  Ica808b9c1910a49740bb889b7521538bc786bf51f6b2c7c3ad1af9712127147b['h00004] ;
//end
//always_comb begin // 
               Iae34f8e78093d5bcc3db929580c94da8015f69b8c6dd2133f36668c2d4b1e0c7['h00003] =  Ica808b9c1910a49740bb889b7521538bc786bf51f6b2c7c3ad1af9712127147b['h00006] ;
//end
//always_comb begin // 
               Iae34f8e78093d5bcc3db929580c94da8015f69b8c6dd2133f36668c2d4b1e0c7['h00004] =  Ica808b9c1910a49740bb889b7521538bc786bf51f6b2c7c3ad1af9712127147b['h00008] ;
//end
//always_comb begin // 
               Iae34f8e78093d5bcc3db929580c94da8015f69b8c6dd2133f36668c2d4b1e0c7['h00005] =  Ica808b9c1910a49740bb889b7521538bc786bf51f6b2c7c3ad1af9712127147b['h0000a] ;
//end
//always_comb begin // 
               Iae34f8e78093d5bcc3db929580c94da8015f69b8c6dd2133f36668c2d4b1e0c7['h00006] =  Ica808b9c1910a49740bb889b7521538bc786bf51f6b2c7c3ad1af9712127147b['h0000c] ;
//end
//always_comb begin // 
               Iae34f8e78093d5bcc3db929580c94da8015f69b8c6dd2133f36668c2d4b1e0c7['h00007] =  Ica808b9c1910a49740bb889b7521538bc786bf51f6b2c7c3ad1af9712127147b['h0000e] ;
//end
