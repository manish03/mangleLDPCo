//`include "GF2_LDPC_fgallag_0x0000d_assign_inc.sv"
//always_comb begin
              I1f3af771a6bf6da6d9e448fb87a2d186['h00000] = 
          (!fgallag_sel['h0000d]) ? 
                       Ia2f891646e6ab8d9fb9ea77d93148790['h00000] : //%
                       Ia2f891646e6ab8d9fb9ea77d93148790['h00001] ;
//end
//always_comb begin
              I1f3af771a6bf6da6d9e448fb87a2d186['h00001] = 
          (!fgallag_sel['h0000d]) ? 
                       Ia2f891646e6ab8d9fb9ea77d93148790['h00002] : //%
                       Ia2f891646e6ab8d9fb9ea77d93148790['h00003] ;
//end
//always_comb begin // 
               I1f3af771a6bf6da6d9e448fb87a2d186['h00002] =  Ia2f891646e6ab8d9fb9ea77d93148790['h00004] ;
//end
//always_comb begin // 
               I1f3af771a6bf6da6d9e448fb87a2d186['h00003] =  Ia2f891646e6ab8d9fb9ea77d93148790['h00006] ;
//end
//always_comb begin // 
               I1f3af771a6bf6da6d9e448fb87a2d186['h00004] =  Ia2f891646e6ab8d9fb9ea77d93148790['h00008] ;
//end
//always_comb begin // 
               I1f3af771a6bf6da6d9e448fb87a2d186['h00005] =  Ia2f891646e6ab8d9fb9ea77d93148790['h0000a] ;
//end
//always_comb begin // 
               I1f3af771a6bf6da6d9e448fb87a2d186['h00006] =  Ia2f891646e6ab8d9fb9ea77d93148790['h0000c] ;
//end
//always_comb begin // 
               I1f3af771a6bf6da6d9e448fb87a2d186['h00007] =  Ia2f891646e6ab8d9fb9ea77d93148790['h0000e] ;
//end
//always_comb begin // 
               I1f3af771a6bf6da6d9e448fb87a2d186['h00008] =  Ia2f891646e6ab8d9fb9ea77d93148790['h00010] ;
//end
//always_comb begin // 
               I1f3af771a6bf6da6d9e448fb87a2d186['h00009] =  Ia2f891646e6ab8d9fb9ea77d93148790['h00012] ;
//end
//always_comb begin // 
               I1f3af771a6bf6da6d9e448fb87a2d186['h0000a] =  Ia2f891646e6ab8d9fb9ea77d93148790['h00014] ;
//end
//always_comb begin // 
               I1f3af771a6bf6da6d9e448fb87a2d186['h0000b] =  Ia2f891646e6ab8d9fb9ea77d93148790['h00016] ;
//end
//always_comb begin // 
               I1f3af771a6bf6da6d9e448fb87a2d186['h0000c] =  Ia2f891646e6ab8d9fb9ea77d93148790['h00018] ;
//end
//always_comb begin // 
               I1f3af771a6bf6da6d9e448fb87a2d186['h0000d] =  Ia2f891646e6ab8d9fb9ea77d93148790['h0001a] ;
//end
//always_comb begin // 
               I1f3af771a6bf6da6d9e448fb87a2d186['h0000e] =  Ia2f891646e6ab8d9fb9ea77d93148790['h0001c] ;
//end
//always_comb begin // 
               I1f3af771a6bf6da6d9e448fb87a2d186['h0000f] =  Ia2f891646e6ab8d9fb9ea77d93148790['h0001e] ;
//end
//always_comb begin // 
               I1f3af771a6bf6da6d9e448fb87a2d186['h00010] =  Ia2f891646e6ab8d9fb9ea77d93148790['h00020] ;
//end
//always_comb begin // 
               I1f3af771a6bf6da6d9e448fb87a2d186['h00011] =  Ia2f891646e6ab8d9fb9ea77d93148790['h00022] ;
//end
//always_comb begin // 
               I1f3af771a6bf6da6d9e448fb87a2d186['h00012] =  Ia2f891646e6ab8d9fb9ea77d93148790['h00024] ;
//end
//always_comb begin // 
               I1f3af771a6bf6da6d9e448fb87a2d186['h00013] =  Ia2f891646e6ab8d9fb9ea77d93148790['h00026] ;
//end
//always_comb begin // 
               I1f3af771a6bf6da6d9e448fb87a2d186['h00014] =  Ia2f891646e6ab8d9fb9ea77d93148790['h00028] ;
//end
//always_comb begin // 
               I1f3af771a6bf6da6d9e448fb87a2d186['h00015] =  Ia2f891646e6ab8d9fb9ea77d93148790['h0002a] ;
//end
//always_comb begin // 
               I1f3af771a6bf6da6d9e448fb87a2d186['h00016] =  Ia2f891646e6ab8d9fb9ea77d93148790['h0002c] ;
//end
//always_comb begin // 
               I1f3af771a6bf6da6d9e448fb87a2d186['h00017] =  Ia2f891646e6ab8d9fb9ea77d93148790['h0002e] ;
//end
//always_comb begin // 
               I1f3af771a6bf6da6d9e448fb87a2d186['h00018] =  Ia2f891646e6ab8d9fb9ea77d93148790['h00030] ;
//end
//always_comb begin // 
               I1f3af771a6bf6da6d9e448fb87a2d186['h00019] =  Ia2f891646e6ab8d9fb9ea77d93148790['h00032] ;
//end
//always_comb begin // 
               I1f3af771a6bf6da6d9e448fb87a2d186['h0001a] =  Ia2f891646e6ab8d9fb9ea77d93148790['h00034] ;
//end
//always_comb begin // 
               I1f3af771a6bf6da6d9e448fb87a2d186['h0001b] =  Ia2f891646e6ab8d9fb9ea77d93148790['h00036] ;
//end
//always_comb begin // 
               I1f3af771a6bf6da6d9e448fb87a2d186['h0001c] =  Ia2f891646e6ab8d9fb9ea77d93148790['h00038] ;
//end
//always_comb begin // 
               I1f3af771a6bf6da6d9e448fb87a2d186['h0001d] =  Ia2f891646e6ab8d9fb9ea77d93148790['h0003a] ;
//end
//always_comb begin // 
               I1f3af771a6bf6da6d9e448fb87a2d186['h0001e] =  Ia2f891646e6ab8d9fb9ea77d93148790['h0003c] ;
//end
//always_comb begin // 
               I1f3af771a6bf6da6d9e448fb87a2d186['h0001f] =  Ia2f891646e6ab8d9fb9ea77d93148790['h0003e] ;
//end
