 reg  ['h7fff:0] [$clog2('h7000+1)-1:0] I2827cdce2a636f7c98629379745844a40e270ed3c43c15a22ae4dfb130ceba7e ;
