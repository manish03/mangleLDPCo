 reg  ['h7:0] [$clog2('h7000+1)-1:0] Ice223344c1d41676e20d7b2668ccff71 ;
