reg [fgallag_WDTH -1:0] fgallag0x00003_0, fgallag0x00003_0_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_1, fgallag0x00003_1_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_2, fgallag0x00003_2_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_3, fgallag0x00003_3_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_4, fgallag0x00003_4_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_5, fgallag0x00003_5_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_6, fgallag0x00003_6_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_7, fgallag0x00003_7_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_8, fgallag0x00003_8_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_9, fgallag0x00003_9_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_10, fgallag0x00003_10_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_11, fgallag0x00003_11_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_12, fgallag0x00003_12_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_13, fgallag0x00003_13_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_14, fgallag0x00003_14_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_15, fgallag0x00003_15_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_16, fgallag0x00003_16_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_17, fgallag0x00003_17_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_18, fgallag0x00003_18_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_19, fgallag0x00003_19_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_20, fgallag0x00003_20_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_21, fgallag0x00003_21_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_22, fgallag0x00003_22_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_23, fgallag0x00003_23_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_24, fgallag0x00003_24_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_25, fgallag0x00003_25_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_26, fgallag0x00003_26_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_27, fgallag0x00003_27_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_28, fgallag0x00003_28_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_29, fgallag0x00003_29_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_30, fgallag0x00003_30_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_31, fgallag0x00003_31_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_32, fgallag0x00003_32_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_33, fgallag0x00003_33_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_34, fgallag0x00003_34_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_35, fgallag0x00003_35_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_36, fgallag0x00003_36_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_37, fgallag0x00003_37_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_38, fgallag0x00003_38_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_39, fgallag0x00003_39_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_40, fgallag0x00003_40_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_41, fgallag0x00003_41_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_42, fgallag0x00003_42_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_43, fgallag0x00003_43_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_44, fgallag0x00003_44_q;
reg [fgallag_WDTH -1:0] fgallag0x00003_45, fgallag0x00003_45_q;
reg start_d_fgallag0x00003_q ;
always @(posedge clk or negedge rstn)
if (!rstn) begin
 fgallag0x00003_0_q <= 'h0;
 fgallag0x00003_1_q <= 'h0;
 fgallag0x00003_2_q <= 'h0;
 fgallag0x00003_3_q <= 'h0;
 fgallag0x00003_4_q <= 'h0;
 fgallag0x00003_5_q <= 'h0;
 fgallag0x00003_6_q <= 'h0;
 fgallag0x00003_7_q <= 'h0;
 fgallag0x00003_8_q <= 'h0;
 fgallag0x00003_9_q <= 'h0;
 fgallag0x00003_10_q <= 'h0;
 fgallag0x00003_11_q <= 'h0;
 fgallag0x00003_12_q <= 'h0;
 fgallag0x00003_13_q <= 'h0;
 fgallag0x00003_14_q <= 'h0;
 fgallag0x00003_15_q <= 'h0;
 fgallag0x00003_16_q <= 'h0;
 fgallag0x00003_17_q <= 'h0;
 fgallag0x00003_18_q <= 'h0;
 fgallag0x00003_19_q <= 'h0;
 fgallag0x00003_20_q <= 'h0;
 fgallag0x00003_21_q <= 'h0;
 fgallag0x00003_22_q <= 'h0;
 fgallag0x00003_23_q <= 'h0;
 fgallag0x00003_24_q <= 'h0;
 fgallag0x00003_25_q <= 'h0;
 fgallag0x00003_26_q <= 'h0;
 fgallag0x00003_27_q <= 'h0;
 fgallag0x00003_28_q <= 'h0;
 fgallag0x00003_29_q <= 'h0;
 fgallag0x00003_30_q <= 'h0;
 fgallag0x00003_31_q <= 'h0;
 fgallag0x00003_32_q <= 'h0;
 fgallag0x00003_33_q <= 'h0;
 fgallag0x00003_34_q <= 'h0;
 fgallag0x00003_35_q <= 'h0;
 fgallag0x00003_36_q <= 'h0;
 fgallag0x00003_37_q <= 'h0;
 fgallag0x00003_38_q <= 'h0;
 fgallag0x00003_39_q <= 'h0;
 fgallag0x00003_40_q <= 'h0;
 fgallag0x00003_41_q <= 'h0;
 fgallag0x00003_42_q <= 'h0;
 fgallag0x00003_43_q <= 'h0;
 fgallag0x00003_44_q <= 'h0;
 fgallag0x00003_45_q <= 'h0;
 start_d_fgallag0x00003_q <= 'h0;
end
else
begin
 fgallag0x00003_0_q <=  fgallag0x00003_0;
 fgallag0x00003_1_q <=  fgallag0x00003_1;
 fgallag0x00003_2_q <=  fgallag0x00003_2;
 fgallag0x00003_3_q <=  fgallag0x00003_3;
 fgallag0x00003_4_q <=  fgallag0x00003_4;
 fgallag0x00003_5_q <=  fgallag0x00003_5;
 fgallag0x00003_6_q <=  fgallag0x00003_6;
 fgallag0x00003_7_q <=  fgallag0x00003_7;
 fgallag0x00003_8_q <=  fgallag0x00003_8;
 fgallag0x00003_9_q <=  fgallag0x00003_9;
 fgallag0x00003_10_q <=  fgallag0x00003_10;
 fgallag0x00003_11_q <=  fgallag0x00003_11;
 fgallag0x00003_12_q <=  fgallag0x00003_12;
 fgallag0x00003_13_q <=  fgallag0x00003_13;
 fgallag0x00003_14_q <=  fgallag0x00003_14;
 fgallag0x00003_15_q <=  fgallag0x00003_15;
 fgallag0x00003_16_q <=  fgallag0x00003_16;
 fgallag0x00003_17_q <=  fgallag0x00003_17;
 fgallag0x00003_18_q <=  fgallag0x00003_18;
 fgallag0x00003_19_q <=  fgallag0x00003_19;
 fgallag0x00003_20_q <=  fgallag0x00003_20;
 fgallag0x00003_21_q <=  fgallag0x00003_21;
 fgallag0x00003_22_q <=  fgallag0x00003_22;
 fgallag0x00003_23_q <=  fgallag0x00003_23;
 fgallag0x00003_24_q <=  fgallag0x00003_24;
 fgallag0x00003_25_q <=  fgallag0x00003_25;
 fgallag0x00003_26_q <=  fgallag0x00003_26;
 fgallag0x00003_27_q <=  fgallag0x00003_27;
 fgallag0x00003_28_q <=  fgallag0x00003_28;
 fgallag0x00003_29_q <=  fgallag0x00003_29;
 fgallag0x00003_30_q <=  fgallag0x00003_30;
 fgallag0x00003_31_q <=  fgallag0x00003_31;
 fgallag0x00003_32_q <=  fgallag0x00003_32;
 fgallag0x00003_33_q <=  fgallag0x00003_33;
 fgallag0x00003_34_q <=  fgallag0x00003_34;
 fgallag0x00003_35_q <=  fgallag0x00003_35;
 fgallag0x00003_36_q <=  fgallag0x00003_36;
 fgallag0x00003_37_q <=  fgallag0x00003_37;
 fgallag0x00003_38_q <=  fgallag0x00003_38;
 fgallag0x00003_39_q <=  fgallag0x00003_39;
 fgallag0x00003_40_q <=  fgallag0x00003_40;
 fgallag0x00003_41_q <=  fgallag0x00003_41;
 fgallag0x00003_42_q <=  fgallag0x00003_42;
 fgallag0x00003_43_q <=  fgallag0x00003_43;
 fgallag0x00003_44_q <=  fgallag0x00003_44;
 fgallag0x00003_45_q <=  fgallag0x00003_45;
 start_d_fgallag0x00003_q <=  start_d_fgallag0x00002_q;
end
