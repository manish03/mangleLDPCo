reg [flogtanh_WDTH -1:0] flogtanh0x00002_0, flogtanh0x00002_0_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_1, flogtanh0x00002_1_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_2, flogtanh0x00002_2_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_3, flogtanh0x00002_3_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_4, flogtanh0x00002_4_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_5, flogtanh0x00002_5_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_6, flogtanh0x00002_6_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_7, flogtanh0x00002_7_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_8, flogtanh0x00002_8_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_9, flogtanh0x00002_9_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_10, flogtanh0x00002_10_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_11, flogtanh0x00002_11_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_12, flogtanh0x00002_12_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_13, flogtanh0x00002_13_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_14, flogtanh0x00002_14_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_15, flogtanh0x00002_15_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_16, flogtanh0x00002_16_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_17, flogtanh0x00002_17_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_18, flogtanh0x00002_18_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_19, flogtanh0x00002_19_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_20, flogtanh0x00002_20_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_21, flogtanh0x00002_21_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_22, flogtanh0x00002_22_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_23, flogtanh0x00002_23_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_24, flogtanh0x00002_24_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_25, flogtanh0x00002_25_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_26, flogtanh0x00002_26_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_27, flogtanh0x00002_27_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_28, flogtanh0x00002_28_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_29, flogtanh0x00002_29_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_30, flogtanh0x00002_30_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_31, flogtanh0x00002_31_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_32, flogtanh0x00002_32_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_33, flogtanh0x00002_33_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_34, flogtanh0x00002_34_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_35, flogtanh0x00002_35_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_36, flogtanh0x00002_36_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_37, flogtanh0x00002_37_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_38, flogtanh0x00002_38_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_39, flogtanh0x00002_39_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_40, flogtanh0x00002_40_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_41, flogtanh0x00002_41_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_42, flogtanh0x00002_42_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_43, flogtanh0x00002_43_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_44, flogtanh0x00002_44_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_45, flogtanh0x00002_45_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_46, flogtanh0x00002_46_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_47, flogtanh0x00002_47_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_48, flogtanh0x00002_48_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_49, flogtanh0x00002_49_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_50, flogtanh0x00002_50_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_51, flogtanh0x00002_51_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_52, flogtanh0x00002_52_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_53, flogtanh0x00002_53_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_54, flogtanh0x00002_54_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_55, flogtanh0x00002_55_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_56, flogtanh0x00002_56_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_57, flogtanh0x00002_57_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_58, flogtanh0x00002_58_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_59, flogtanh0x00002_59_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_60, flogtanh0x00002_60_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_61, flogtanh0x00002_61_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_62, flogtanh0x00002_62_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_63, flogtanh0x00002_63_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_64, flogtanh0x00002_64_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_65, flogtanh0x00002_65_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_66, flogtanh0x00002_66_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_67, flogtanh0x00002_67_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_68, flogtanh0x00002_68_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_69, flogtanh0x00002_69_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_70, flogtanh0x00002_70_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_71, flogtanh0x00002_71_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_72, flogtanh0x00002_72_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_73, flogtanh0x00002_73_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_74, flogtanh0x00002_74_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_75, flogtanh0x00002_75_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_76, flogtanh0x00002_76_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_77, flogtanh0x00002_77_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_78, flogtanh0x00002_78_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_79, flogtanh0x00002_79_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_80, flogtanh0x00002_80_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_81, flogtanh0x00002_81_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_82, flogtanh0x00002_82_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_83, flogtanh0x00002_83_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_84, flogtanh0x00002_84_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_85, flogtanh0x00002_85_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_86, flogtanh0x00002_86_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_87, flogtanh0x00002_87_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_88, flogtanh0x00002_88_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00002_89, flogtanh0x00002_89_q;
reg start_d_flogtanh0x00002_q ;
always @(posedge clk or negedge rstn)
if (!rstn) begin
 flogtanh0x00002_0_q <= 'h0;
 flogtanh0x00002_1_q <= 'h0;
 flogtanh0x00002_2_q <= 'h0;
 flogtanh0x00002_3_q <= 'h0;
 flogtanh0x00002_4_q <= 'h0;
 flogtanh0x00002_5_q <= 'h0;
 flogtanh0x00002_6_q <= 'h0;
 flogtanh0x00002_7_q <= 'h0;
 flogtanh0x00002_8_q <= 'h0;
 flogtanh0x00002_9_q <= 'h0;
 flogtanh0x00002_10_q <= 'h0;
 flogtanh0x00002_11_q <= 'h0;
 flogtanh0x00002_12_q <= 'h0;
 flogtanh0x00002_13_q <= 'h0;
 flogtanh0x00002_14_q <= 'h0;
 flogtanh0x00002_15_q <= 'h0;
 flogtanh0x00002_16_q <= 'h0;
 flogtanh0x00002_17_q <= 'h0;
 flogtanh0x00002_18_q <= 'h0;
 flogtanh0x00002_19_q <= 'h0;
 flogtanh0x00002_20_q <= 'h0;
 flogtanh0x00002_21_q <= 'h0;
 flogtanh0x00002_22_q <= 'h0;
 flogtanh0x00002_23_q <= 'h0;
 flogtanh0x00002_24_q <= 'h0;
 flogtanh0x00002_25_q <= 'h0;
 flogtanh0x00002_26_q <= 'h0;
 flogtanh0x00002_27_q <= 'h0;
 flogtanh0x00002_28_q <= 'h0;
 flogtanh0x00002_29_q <= 'h0;
 flogtanh0x00002_30_q <= 'h0;
 flogtanh0x00002_31_q <= 'h0;
 flogtanh0x00002_32_q <= 'h0;
 flogtanh0x00002_33_q <= 'h0;
 flogtanh0x00002_34_q <= 'h0;
 flogtanh0x00002_35_q <= 'h0;
 flogtanh0x00002_36_q <= 'h0;
 flogtanh0x00002_37_q <= 'h0;
 flogtanh0x00002_38_q <= 'h0;
 flogtanh0x00002_39_q <= 'h0;
 flogtanh0x00002_40_q <= 'h0;
 flogtanh0x00002_41_q <= 'h0;
 flogtanh0x00002_42_q <= 'h0;
 flogtanh0x00002_43_q <= 'h0;
 flogtanh0x00002_44_q <= 'h0;
 flogtanh0x00002_45_q <= 'h0;
 flogtanh0x00002_46_q <= 'h0;
 flogtanh0x00002_47_q <= 'h0;
 flogtanh0x00002_48_q <= 'h0;
 flogtanh0x00002_49_q <= 'h0;
 flogtanh0x00002_50_q <= 'h0;
 flogtanh0x00002_51_q <= 'h0;
 flogtanh0x00002_52_q <= 'h0;
 flogtanh0x00002_53_q <= 'h0;
 flogtanh0x00002_54_q <= 'h0;
 flogtanh0x00002_55_q <= 'h0;
 flogtanh0x00002_56_q <= 'h0;
 flogtanh0x00002_57_q <= 'h0;
 flogtanh0x00002_58_q <= 'h0;
 flogtanh0x00002_59_q <= 'h0;
 flogtanh0x00002_60_q <= 'h0;
 flogtanh0x00002_61_q <= 'h0;
 flogtanh0x00002_62_q <= 'h0;
 flogtanh0x00002_63_q <= 'h0;
 flogtanh0x00002_64_q <= 'h0;
 flogtanh0x00002_65_q <= 'h0;
 flogtanh0x00002_66_q <= 'h0;
 flogtanh0x00002_67_q <= 'h0;
 flogtanh0x00002_68_q <= 'h0;
 flogtanh0x00002_69_q <= 'h0;
 flogtanh0x00002_70_q <= 'h0;
 flogtanh0x00002_71_q <= 'h0;
 flogtanh0x00002_72_q <= 'h0;
 flogtanh0x00002_73_q <= 'h0;
 flogtanh0x00002_74_q <= 'h0;
 flogtanh0x00002_75_q <= 'h0;
 flogtanh0x00002_76_q <= 'h0;
 flogtanh0x00002_77_q <= 'h0;
 flogtanh0x00002_78_q <= 'h0;
 flogtanh0x00002_79_q <= 'h0;
 flogtanh0x00002_80_q <= 'h0;
 flogtanh0x00002_81_q <= 'h0;
 flogtanh0x00002_82_q <= 'h0;
 flogtanh0x00002_83_q <= 'h0;
 flogtanh0x00002_84_q <= 'h0;
 flogtanh0x00002_85_q <= 'h0;
 flogtanh0x00002_86_q <= 'h0;
 flogtanh0x00002_87_q <= 'h0;
 flogtanh0x00002_88_q <= 'h0;
 flogtanh0x00002_89_q <= 'h0;
 start_d_flogtanh0x00002_q <= 'h0;
end
else
begin
 flogtanh0x00002_0_q <=  flogtanh0x00002_0;
 flogtanh0x00002_1_q <=  flogtanh0x00002_1;
 flogtanh0x00002_2_q <=  flogtanh0x00002_2;
 flogtanh0x00002_3_q <=  flogtanh0x00002_3;
 flogtanh0x00002_4_q <=  flogtanh0x00002_4;
 flogtanh0x00002_5_q <=  flogtanh0x00002_5;
 flogtanh0x00002_6_q <=  flogtanh0x00002_6;
 flogtanh0x00002_7_q <=  flogtanh0x00002_7;
 flogtanh0x00002_8_q <=  flogtanh0x00002_8;
 flogtanh0x00002_9_q <=  flogtanh0x00002_9;
 flogtanh0x00002_10_q <=  flogtanh0x00002_10;
 flogtanh0x00002_11_q <=  flogtanh0x00002_11;
 flogtanh0x00002_12_q <=  flogtanh0x00002_12;
 flogtanh0x00002_13_q <=  flogtanh0x00002_13;
 flogtanh0x00002_14_q <=  flogtanh0x00002_14;
 flogtanh0x00002_15_q <=  flogtanh0x00002_15;
 flogtanh0x00002_16_q <=  flogtanh0x00002_16;
 flogtanh0x00002_17_q <=  flogtanh0x00002_17;
 flogtanh0x00002_18_q <=  flogtanh0x00002_18;
 flogtanh0x00002_19_q <=  flogtanh0x00002_19;
 flogtanh0x00002_20_q <=  flogtanh0x00002_20;
 flogtanh0x00002_21_q <=  flogtanh0x00002_21;
 flogtanh0x00002_22_q <=  flogtanh0x00002_22;
 flogtanh0x00002_23_q <=  flogtanh0x00002_23;
 flogtanh0x00002_24_q <=  flogtanh0x00002_24;
 flogtanh0x00002_25_q <=  flogtanh0x00002_25;
 flogtanh0x00002_26_q <=  flogtanh0x00002_26;
 flogtanh0x00002_27_q <=  flogtanh0x00002_27;
 flogtanh0x00002_28_q <=  flogtanh0x00002_28;
 flogtanh0x00002_29_q <=  flogtanh0x00002_29;
 flogtanh0x00002_30_q <=  flogtanh0x00002_30;
 flogtanh0x00002_31_q <=  flogtanh0x00002_31;
 flogtanh0x00002_32_q <=  flogtanh0x00002_32;
 flogtanh0x00002_33_q <=  flogtanh0x00002_33;
 flogtanh0x00002_34_q <=  flogtanh0x00002_34;
 flogtanh0x00002_35_q <=  flogtanh0x00002_35;
 flogtanh0x00002_36_q <=  flogtanh0x00002_36;
 flogtanh0x00002_37_q <=  flogtanh0x00002_37;
 flogtanh0x00002_38_q <=  flogtanh0x00002_38;
 flogtanh0x00002_39_q <=  flogtanh0x00002_39;
 flogtanh0x00002_40_q <=  flogtanh0x00002_40;
 flogtanh0x00002_41_q <=  flogtanh0x00002_41;
 flogtanh0x00002_42_q <=  flogtanh0x00002_42;
 flogtanh0x00002_43_q <=  flogtanh0x00002_43;
 flogtanh0x00002_44_q <=  flogtanh0x00002_44;
 flogtanh0x00002_45_q <=  flogtanh0x00002_45;
 flogtanh0x00002_46_q <=  flogtanh0x00002_46;
 flogtanh0x00002_47_q <=  flogtanh0x00002_47;
 flogtanh0x00002_48_q <=  flogtanh0x00002_48;
 flogtanh0x00002_49_q <=  flogtanh0x00002_49;
 flogtanh0x00002_50_q <=  flogtanh0x00002_50;
 flogtanh0x00002_51_q <=  flogtanh0x00002_51;
 flogtanh0x00002_52_q <=  flogtanh0x00002_52;
 flogtanh0x00002_53_q <=  flogtanh0x00002_53;
 flogtanh0x00002_54_q <=  flogtanh0x00002_54;
 flogtanh0x00002_55_q <=  flogtanh0x00002_55;
 flogtanh0x00002_56_q <=  flogtanh0x00002_56;
 flogtanh0x00002_57_q <=  flogtanh0x00002_57;
 flogtanh0x00002_58_q <=  flogtanh0x00002_58;
 flogtanh0x00002_59_q <=  flogtanh0x00002_59;
 flogtanh0x00002_60_q <=  flogtanh0x00002_60;
 flogtanh0x00002_61_q <=  flogtanh0x00002_61;
 flogtanh0x00002_62_q <=  flogtanh0x00002_62;
 flogtanh0x00002_63_q <=  flogtanh0x00002_63;
 flogtanh0x00002_64_q <=  flogtanh0x00002_64;
 flogtanh0x00002_65_q <=  flogtanh0x00002_65;
 flogtanh0x00002_66_q <=  flogtanh0x00002_66;
 flogtanh0x00002_67_q <=  flogtanh0x00002_67;
 flogtanh0x00002_68_q <=  flogtanh0x00002_68;
 flogtanh0x00002_69_q <=  flogtanh0x00002_69;
 flogtanh0x00002_70_q <=  flogtanh0x00002_70;
 flogtanh0x00002_71_q <=  flogtanh0x00002_71;
 flogtanh0x00002_72_q <=  flogtanh0x00002_72;
 flogtanh0x00002_73_q <=  flogtanh0x00002_73;
 flogtanh0x00002_74_q <=  flogtanh0x00002_74;
 flogtanh0x00002_75_q <=  flogtanh0x00002_75;
 flogtanh0x00002_76_q <=  flogtanh0x00002_76;
 flogtanh0x00002_77_q <=  flogtanh0x00002_77;
 flogtanh0x00002_78_q <=  flogtanh0x00002_78;
 flogtanh0x00002_79_q <=  flogtanh0x00002_79;
 flogtanh0x00002_80_q <=  flogtanh0x00002_80;
 flogtanh0x00002_81_q <=  flogtanh0x00002_81;
 flogtanh0x00002_82_q <=  flogtanh0x00002_82;
 flogtanh0x00002_83_q <=  flogtanh0x00002_83;
 flogtanh0x00002_84_q <=  flogtanh0x00002_84;
 flogtanh0x00002_85_q <=  flogtanh0x00002_85;
 flogtanh0x00002_86_q <=  flogtanh0x00002_86;
 flogtanh0x00002_87_q <=  flogtanh0x00002_87;
 flogtanh0x00002_88_q <=  flogtanh0x00002_88;
 flogtanh0x00002_89_q <=  flogtanh0x00002_89;
 start_d_flogtanh0x00002_q <=  start_d_flogtanh0x00001_q;
end
