 reg  ['hf:0] [$clog2('h7000+1)-1:0] Ica808b9c1910a49740bb889b7521538bc786bf51f6b2c7c3ad1af9712127147b ;
