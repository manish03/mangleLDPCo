//`include "GF2_LDPC_flogtanh_0x00008_assign_inc.sv"
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h00000] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h00000] : //%
                       I38e438ab568822a1c40149a2acc5d876['h00001] ;
//end
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h00001] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h00002] : //%
                       I38e438ab568822a1c40149a2acc5d876['h00003] ;
//end
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h00002] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h00004] : //%
                       I38e438ab568822a1c40149a2acc5d876['h00005] ;
//end
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h00003] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h00006] : //%
                       I38e438ab568822a1c40149a2acc5d876['h00007] ;
//end
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h00004] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h00008] : //%
                       I38e438ab568822a1c40149a2acc5d876['h00009] ;
//end
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h00005] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h0000a] : //%
                       I38e438ab568822a1c40149a2acc5d876['h0000b] ;
//end
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h00006] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h0000c] : //%
                       I38e438ab568822a1c40149a2acc5d876['h0000d] ;
//end
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h00007] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h0000e] : //%
                       I38e438ab568822a1c40149a2acc5d876['h0000f] ;
//end
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h00008] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h00010] : //%
                       I38e438ab568822a1c40149a2acc5d876['h00011] ;
//end
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h00009] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h00012] : //%
                       I38e438ab568822a1c40149a2acc5d876['h00013] ;
//end
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h0000a] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h00014] : //%
                       I38e438ab568822a1c40149a2acc5d876['h00015] ;
//end
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h0000b] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h00016] : //%
                       I38e438ab568822a1c40149a2acc5d876['h00017] ;
//end
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h0000c] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h00018] : //%
                       I38e438ab568822a1c40149a2acc5d876['h00019] ;
//end
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h0000d] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h0001a] : //%
                       I38e438ab568822a1c40149a2acc5d876['h0001b] ;
//end
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h0000e] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h0001c] : //%
                       I38e438ab568822a1c40149a2acc5d876['h0001d] ;
//end
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h0000f] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h0001e] : //%
                       I38e438ab568822a1c40149a2acc5d876['h0001f] ;
//end
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h00010] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h00020] : //%
                       I38e438ab568822a1c40149a2acc5d876['h00021] ;
//end
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h00011] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h00022] : //%
                       I38e438ab568822a1c40149a2acc5d876['h00023] ;
//end
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h00012] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h00024] : //%
                       I38e438ab568822a1c40149a2acc5d876['h00025] ;
//end
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h00013] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h00026] : //%
                       I38e438ab568822a1c40149a2acc5d876['h00027] ;
//end
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h00014] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h00028] : //%
                       I38e438ab568822a1c40149a2acc5d876['h00029] ;
//end
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h00015] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h0002a] : //%
                       I38e438ab568822a1c40149a2acc5d876['h0002b] ;
//end
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h00016] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h0002c] : //%
                       I38e438ab568822a1c40149a2acc5d876['h0002d] ;
//end
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h00017] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h0002e] : //%
                       I38e438ab568822a1c40149a2acc5d876['h0002f] ;
//end
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h00018] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h00030] : //%
                       I38e438ab568822a1c40149a2acc5d876['h00031] ;
//end
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h00019] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h00032] : //%
                       I38e438ab568822a1c40149a2acc5d876['h00033] ;
//end
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h0001a] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h00034] : //%
                       I38e438ab568822a1c40149a2acc5d876['h00035] ;
//end
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h0001b] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h00036] : //%
                       I38e438ab568822a1c40149a2acc5d876['h00037] ;
//end
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h0001c] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h00038] : //%
                       I38e438ab568822a1c40149a2acc5d876['h00039] ;
//end
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h0001d] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h0003a] : //%
                       I38e438ab568822a1c40149a2acc5d876['h0003b] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0001e] =  I38e438ab568822a1c40149a2acc5d876['h0003c] ;
//end
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h0001f] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h0003e] : //%
                       I38e438ab568822a1c40149a2acc5d876['h0003f] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00020] =  I38e438ab568822a1c40149a2acc5d876['h00040] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00021] =  I38e438ab568822a1c40149a2acc5d876['h00042] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00022] =  I38e438ab568822a1c40149a2acc5d876['h00044] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00023] =  I38e438ab568822a1c40149a2acc5d876['h00046] ;
//end
//always_comb begin
              I810764ca41a2b12d686e115c79b0578f['h00024] = 
          (!flogtanh_sel['h00008]) ? 
                       I38e438ab568822a1c40149a2acc5d876['h00048] : //%
                       I38e438ab568822a1c40149a2acc5d876['h00049] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00025] =  I38e438ab568822a1c40149a2acc5d876['h0004a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00026] =  I38e438ab568822a1c40149a2acc5d876['h0004c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00027] =  I38e438ab568822a1c40149a2acc5d876['h0004e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00028] =  I38e438ab568822a1c40149a2acc5d876['h00050] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00029] =  I38e438ab568822a1c40149a2acc5d876['h00052] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0002a] =  I38e438ab568822a1c40149a2acc5d876['h00054] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0002b] =  I38e438ab568822a1c40149a2acc5d876['h00056] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0002c] =  I38e438ab568822a1c40149a2acc5d876['h00058] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0002d] =  I38e438ab568822a1c40149a2acc5d876['h0005a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0002e] =  I38e438ab568822a1c40149a2acc5d876['h0005c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0002f] =  I38e438ab568822a1c40149a2acc5d876['h0005e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00030] =  I38e438ab568822a1c40149a2acc5d876['h00060] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00031] =  I38e438ab568822a1c40149a2acc5d876['h00062] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00032] =  I38e438ab568822a1c40149a2acc5d876['h00064] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00033] =  I38e438ab568822a1c40149a2acc5d876['h00066] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00034] =  I38e438ab568822a1c40149a2acc5d876['h00068] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00035] =  I38e438ab568822a1c40149a2acc5d876['h0006a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00036] =  I38e438ab568822a1c40149a2acc5d876['h0006c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00037] =  I38e438ab568822a1c40149a2acc5d876['h0006e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00038] =  I38e438ab568822a1c40149a2acc5d876['h00070] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00039] =  I38e438ab568822a1c40149a2acc5d876['h00072] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0003a] =  I38e438ab568822a1c40149a2acc5d876['h00074] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0003b] =  I38e438ab568822a1c40149a2acc5d876['h00076] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0003c] =  I38e438ab568822a1c40149a2acc5d876['h00078] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0003d] =  I38e438ab568822a1c40149a2acc5d876['h0007a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0003e] =  I38e438ab568822a1c40149a2acc5d876['h0007c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0003f] =  I38e438ab568822a1c40149a2acc5d876['h0007e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00040] =  I38e438ab568822a1c40149a2acc5d876['h00080] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00041] =  I38e438ab568822a1c40149a2acc5d876['h00082] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00042] =  I38e438ab568822a1c40149a2acc5d876['h00084] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00043] =  I38e438ab568822a1c40149a2acc5d876['h00086] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00044] =  I38e438ab568822a1c40149a2acc5d876['h00088] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00045] =  I38e438ab568822a1c40149a2acc5d876['h0008a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00046] =  I38e438ab568822a1c40149a2acc5d876['h0008c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00047] =  I38e438ab568822a1c40149a2acc5d876['h0008e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00048] =  I38e438ab568822a1c40149a2acc5d876['h00090] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00049] =  I38e438ab568822a1c40149a2acc5d876['h00092] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0004a] =  I38e438ab568822a1c40149a2acc5d876['h00094] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0004b] =  I38e438ab568822a1c40149a2acc5d876['h00096] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0004c] =  I38e438ab568822a1c40149a2acc5d876['h00098] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0004d] =  I38e438ab568822a1c40149a2acc5d876['h0009a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0004e] =  I38e438ab568822a1c40149a2acc5d876['h0009c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0004f] =  I38e438ab568822a1c40149a2acc5d876['h0009e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00050] =  I38e438ab568822a1c40149a2acc5d876['h000a0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00051] =  I38e438ab568822a1c40149a2acc5d876['h000a2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00052] =  I38e438ab568822a1c40149a2acc5d876['h000a4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00053] =  I38e438ab568822a1c40149a2acc5d876['h000a6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00054] =  I38e438ab568822a1c40149a2acc5d876['h000a8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00055] =  I38e438ab568822a1c40149a2acc5d876['h000aa] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00056] =  I38e438ab568822a1c40149a2acc5d876['h000ac] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00057] =  I38e438ab568822a1c40149a2acc5d876['h000ae] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00058] =  I38e438ab568822a1c40149a2acc5d876['h000b0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00059] =  I38e438ab568822a1c40149a2acc5d876['h000b2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0005a] =  I38e438ab568822a1c40149a2acc5d876['h000b4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0005b] =  I38e438ab568822a1c40149a2acc5d876['h000b6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0005c] =  I38e438ab568822a1c40149a2acc5d876['h000b8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0005d] =  I38e438ab568822a1c40149a2acc5d876['h000ba] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0005e] =  I38e438ab568822a1c40149a2acc5d876['h000bc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0005f] =  I38e438ab568822a1c40149a2acc5d876['h000be] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00060] =  I38e438ab568822a1c40149a2acc5d876['h000c0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00061] =  I38e438ab568822a1c40149a2acc5d876['h000c2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00062] =  I38e438ab568822a1c40149a2acc5d876['h000c4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00063] =  I38e438ab568822a1c40149a2acc5d876['h000c6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00064] =  I38e438ab568822a1c40149a2acc5d876['h000c8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00065] =  I38e438ab568822a1c40149a2acc5d876['h000ca] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00066] =  I38e438ab568822a1c40149a2acc5d876['h000cc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00067] =  I38e438ab568822a1c40149a2acc5d876['h000ce] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00068] =  I38e438ab568822a1c40149a2acc5d876['h000d0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00069] =  I38e438ab568822a1c40149a2acc5d876['h000d2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0006a] =  I38e438ab568822a1c40149a2acc5d876['h000d4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0006b] =  I38e438ab568822a1c40149a2acc5d876['h000d6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0006c] =  I38e438ab568822a1c40149a2acc5d876['h000d8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0006d] =  I38e438ab568822a1c40149a2acc5d876['h000da] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0006e] =  I38e438ab568822a1c40149a2acc5d876['h000dc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0006f] =  I38e438ab568822a1c40149a2acc5d876['h000de] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00070] =  I38e438ab568822a1c40149a2acc5d876['h000e0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00071] =  I38e438ab568822a1c40149a2acc5d876['h000e2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00072] =  I38e438ab568822a1c40149a2acc5d876['h000e4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00073] =  I38e438ab568822a1c40149a2acc5d876['h000e6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00074] =  I38e438ab568822a1c40149a2acc5d876['h000e8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00075] =  I38e438ab568822a1c40149a2acc5d876['h000ea] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00076] =  I38e438ab568822a1c40149a2acc5d876['h000ec] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00077] =  I38e438ab568822a1c40149a2acc5d876['h000ee] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00078] =  I38e438ab568822a1c40149a2acc5d876['h000f0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00079] =  I38e438ab568822a1c40149a2acc5d876['h000f2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0007a] =  I38e438ab568822a1c40149a2acc5d876['h000f4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0007b] =  I38e438ab568822a1c40149a2acc5d876['h000f6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0007c] =  I38e438ab568822a1c40149a2acc5d876['h000f8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0007d] =  I38e438ab568822a1c40149a2acc5d876['h000fa] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0007e] =  I38e438ab568822a1c40149a2acc5d876['h000fc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0007f] =  I38e438ab568822a1c40149a2acc5d876['h000fe] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00080] =  I38e438ab568822a1c40149a2acc5d876['h00100] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00081] =  I38e438ab568822a1c40149a2acc5d876['h00102] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00082] =  I38e438ab568822a1c40149a2acc5d876['h00104] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00083] =  I38e438ab568822a1c40149a2acc5d876['h00106] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00084] =  I38e438ab568822a1c40149a2acc5d876['h00108] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00085] =  I38e438ab568822a1c40149a2acc5d876['h0010a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00086] =  I38e438ab568822a1c40149a2acc5d876['h0010c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00087] =  I38e438ab568822a1c40149a2acc5d876['h0010e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00088] =  I38e438ab568822a1c40149a2acc5d876['h00110] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00089] =  I38e438ab568822a1c40149a2acc5d876['h00112] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0008a] =  I38e438ab568822a1c40149a2acc5d876['h00114] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0008b] =  I38e438ab568822a1c40149a2acc5d876['h00116] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0008c] =  I38e438ab568822a1c40149a2acc5d876['h00118] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0008d] =  I38e438ab568822a1c40149a2acc5d876['h0011a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0008e] =  I38e438ab568822a1c40149a2acc5d876['h0011c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0008f] =  I38e438ab568822a1c40149a2acc5d876['h0011e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00090] =  I38e438ab568822a1c40149a2acc5d876['h00120] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00091] =  I38e438ab568822a1c40149a2acc5d876['h00122] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00092] =  I38e438ab568822a1c40149a2acc5d876['h00124] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00093] =  I38e438ab568822a1c40149a2acc5d876['h00126] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00094] =  I38e438ab568822a1c40149a2acc5d876['h00128] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00095] =  I38e438ab568822a1c40149a2acc5d876['h0012a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00096] =  I38e438ab568822a1c40149a2acc5d876['h0012c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00097] =  I38e438ab568822a1c40149a2acc5d876['h0012e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00098] =  I38e438ab568822a1c40149a2acc5d876['h00130] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00099] =  I38e438ab568822a1c40149a2acc5d876['h00132] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0009a] =  I38e438ab568822a1c40149a2acc5d876['h00134] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0009b] =  I38e438ab568822a1c40149a2acc5d876['h00136] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0009c] =  I38e438ab568822a1c40149a2acc5d876['h00138] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0009d] =  I38e438ab568822a1c40149a2acc5d876['h0013a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0009e] =  I38e438ab568822a1c40149a2acc5d876['h0013c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0009f] =  I38e438ab568822a1c40149a2acc5d876['h0013e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000a0] =  I38e438ab568822a1c40149a2acc5d876['h00140] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000a1] =  I38e438ab568822a1c40149a2acc5d876['h00142] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000a2] =  I38e438ab568822a1c40149a2acc5d876['h00144] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000a3] =  I38e438ab568822a1c40149a2acc5d876['h00146] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000a4] =  I38e438ab568822a1c40149a2acc5d876['h00148] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000a5] =  I38e438ab568822a1c40149a2acc5d876['h0014a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000a6] =  I38e438ab568822a1c40149a2acc5d876['h0014c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000a7] =  I38e438ab568822a1c40149a2acc5d876['h0014e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000a8] =  I38e438ab568822a1c40149a2acc5d876['h00150] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000a9] =  I38e438ab568822a1c40149a2acc5d876['h00152] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000aa] =  I38e438ab568822a1c40149a2acc5d876['h00154] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000ab] =  I38e438ab568822a1c40149a2acc5d876['h00156] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000ac] =  I38e438ab568822a1c40149a2acc5d876['h00158] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000ad] =  I38e438ab568822a1c40149a2acc5d876['h0015a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000ae] =  I38e438ab568822a1c40149a2acc5d876['h0015c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000af] =  I38e438ab568822a1c40149a2acc5d876['h0015e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000b0] =  I38e438ab568822a1c40149a2acc5d876['h00160] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000b1] =  I38e438ab568822a1c40149a2acc5d876['h00162] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000b2] =  I38e438ab568822a1c40149a2acc5d876['h00164] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000b3] =  I38e438ab568822a1c40149a2acc5d876['h00166] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000b4] =  I38e438ab568822a1c40149a2acc5d876['h00168] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000b5] =  I38e438ab568822a1c40149a2acc5d876['h0016a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000b6] =  I38e438ab568822a1c40149a2acc5d876['h0016c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000b7] =  I38e438ab568822a1c40149a2acc5d876['h0016e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000b8] =  I38e438ab568822a1c40149a2acc5d876['h00170] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000b9] =  I38e438ab568822a1c40149a2acc5d876['h00172] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000ba] =  I38e438ab568822a1c40149a2acc5d876['h00174] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000bb] =  I38e438ab568822a1c40149a2acc5d876['h00176] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000bc] =  I38e438ab568822a1c40149a2acc5d876['h00178] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000bd] =  I38e438ab568822a1c40149a2acc5d876['h0017a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000be] =  I38e438ab568822a1c40149a2acc5d876['h0017c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000bf] =  I38e438ab568822a1c40149a2acc5d876['h0017e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000c0] =  I38e438ab568822a1c40149a2acc5d876['h00180] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000c1] =  I38e438ab568822a1c40149a2acc5d876['h00182] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000c2] =  I38e438ab568822a1c40149a2acc5d876['h00184] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000c3] =  I38e438ab568822a1c40149a2acc5d876['h00186] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000c4] =  I38e438ab568822a1c40149a2acc5d876['h00188] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000c5] =  I38e438ab568822a1c40149a2acc5d876['h0018a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000c6] =  I38e438ab568822a1c40149a2acc5d876['h0018c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000c7] =  I38e438ab568822a1c40149a2acc5d876['h0018e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000c8] =  I38e438ab568822a1c40149a2acc5d876['h00190] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000c9] =  I38e438ab568822a1c40149a2acc5d876['h00192] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000ca] =  I38e438ab568822a1c40149a2acc5d876['h00194] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000cb] =  I38e438ab568822a1c40149a2acc5d876['h00196] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000cc] =  I38e438ab568822a1c40149a2acc5d876['h00198] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000cd] =  I38e438ab568822a1c40149a2acc5d876['h0019a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000ce] =  I38e438ab568822a1c40149a2acc5d876['h0019c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000cf] =  I38e438ab568822a1c40149a2acc5d876['h0019e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000d0] =  I38e438ab568822a1c40149a2acc5d876['h001a0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000d1] =  I38e438ab568822a1c40149a2acc5d876['h001a2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000d2] =  I38e438ab568822a1c40149a2acc5d876['h001a4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000d3] =  I38e438ab568822a1c40149a2acc5d876['h001a6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000d4] =  I38e438ab568822a1c40149a2acc5d876['h001a8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000d5] =  I38e438ab568822a1c40149a2acc5d876['h001aa] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000d6] =  I38e438ab568822a1c40149a2acc5d876['h001ac] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000d7] =  I38e438ab568822a1c40149a2acc5d876['h001ae] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000d8] =  I38e438ab568822a1c40149a2acc5d876['h001b0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000d9] =  I38e438ab568822a1c40149a2acc5d876['h001b2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000da] =  I38e438ab568822a1c40149a2acc5d876['h001b4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000db] =  I38e438ab568822a1c40149a2acc5d876['h001b6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000dc] =  I38e438ab568822a1c40149a2acc5d876['h001b8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000dd] =  I38e438ab568822a1c40149a2acc5d876['h001ba] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000de] =  I38e438ab568822a1c40149a2acc5d876['h001bc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000df] =  I38e438ab568822a1c40149a2acc5d876['h001be] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000e0] =  I38e438ab568822a1c40149a2acc5d876['h001c0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000e1] =  I38e438ab568822a1c40149a2acc5d876['h001c2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000e2] =  I38e438ab568822a1c40149a2acc5d876['h001c4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000e3] =  I38e438ab568822a1c40149a2acc5d876['h001c6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000e4] =  I38e438ab568822a1c40149a2acc5d876['h001c8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000e5] =  I38e438ab568822a1c40149a2acc5d876['h001ca] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000e6] =  I38e438ab568822a1c40149a2acc5d876['h001cc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000e7] =  I38e438ab568822a1c40149a2acc5d876['h001ce] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000e8] =  I38e438ab568822a1c40149a2acc5d876['h001d0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000e9] =  I38e438ab568822a1c40149a2acc5d876['h001d2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000ea] =  I38e438ab568822a1c40149a2acc5d876['h001d4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000eb] =  I38e438ab568822a1c40149a2acc5d876['h001d6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000ec] =  I38e438ab568822a1c40149a2acc5d876['h001d8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000ed] =  I38e438ab568822a1c40149a2acc5d876['h001da] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000ee] =  I38e438ab568822a1c40149a2acc5d876['h001dc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000ef] =  I38e438ab568822a1c40149a2acc5d876['h001de] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000f0] =  I38e438ab568822a1c40149a2acc5d876['h001e0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000f1] =  I38e438ab568822a1c40149a2acc5d876['h001e2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000f2] =  I38e438ab568822a1c40149a2acc5d876['h001e4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000f3] =  I38e438ab568822a1c40149a2acc5d876['h001e6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000f4] =  I38e438ab568822a1c40149a2acc5d876['h001e8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000f5] =  I38e438ab568822a1c40149a2acc5d876['h001ea] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000f6] =  I38e438ab568822a1c40149a2acc5d876['h001ec] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000f7] =  I38e438ab568822a1c40149a2acc5d876['h001ee] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000f8] =  I38e438ab568822a1c40149a2acc5d876['h001f0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000f9] =  I38e438ab568822a1c40149a2acc5d876['h001f2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000fa] =  I38e438ab568822a1c40149a2acc5d876['h001f4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000fb] =  I38e438ab568822a1c40149a2acc5d876['h001f6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000fc] =  I38e438ab568822a1c40149a2acc5d876['h001f8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000fd] =  I38e438ab568822a1c40149a2acc5d876['h001fa] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000fe] =  I38e438ab568822a1c40149a2acc5d876['h001fc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h000ff] =  I38e438ab568822a1c40149a2acc5d876['h001fe] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00100] =  I38e438ab568822a1c40149a2acc5d876['h00200] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00101] =  I38e438ab568822a1c40149a2acc5d876['h00202] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00102] =  I38e438ab568822a1c40149a2acc5d876['h00204] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00103] =  I38e438ab568822a1c40149a2acc5d876['h00206] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00104] =  I38e438ab568822a1c40149a2acc5d876['h00208] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00105] =  I38e438ab568822a1c40149a2acc5d876['h0020a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00106] =  I38e438ab568822a1c40149a2acc5d876['h0020c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00107] =  I38e438ab568822a1c40149a2acc5d876['h0020e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00108] =  I38e438ab568822a1c40149a2acc5d876['h00210] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00109] =  I38e438ab568822a1c40149a2acc5d876['h00212] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0010a] =  I38e438ab568822a1c40149a2acc5d876['h00214] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0010b] =  I38e438ab568822a1c40149a2acc5d876['h00216] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0010c] =  I38e438ab568822a1c40149a2acc5d876['h00218] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0010d] =  I38e438ab568822a1c40149a2acc5d876['h0021a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0010e] =  I38e438ab568822a1c40149a2acc5d876['h0021c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0010f] =  I38e438ab568822a1c40149a2acc5d876['h0021e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00110] =  I38e438ab568822a1c40149a2acc5d876['h00220] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00111] =  I38e438ab568822a1c40149a2acc5d876['h00222] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00112] =  I38e438ab568822a1c40149a2acc5d876['h00224] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00113] =  I38e438ab568822a1c40149a2acc5d876['h00226] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00114] =  I38e438ab568822a1c40149a2acc5d876['h00228] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00115] =  I38e438ab568822a1c40149a2acc5d876['h0022a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00116] =  I38e438ab568822a1c40149a2acc5d876['h0022c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00117] =  I38e438ab568822a1c40149a2acc5d876['h0022e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00118] =  I38e438ab568822a1c40149a2acc5d876['h00230] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00119] =  I38e438ab568822a1c40149a2acc5d876['h00232] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0011a] =  I38e438ab568822a1c40149a2acc5d876['h00234] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0011b] =  I38e438ab568822a1c40149a2acc5d876['h00236] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0011c] =  I38e438ab568822a1c40149a2acc5d876['h00238] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0011d] =  I38e438ab568822a1c40149a2acc5d876['h0023a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0011e] =  I38e438ab568822a1c40149a2acc5d876['h0023c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0011f] =  I38e438ab568822a1c40149a2acc5d876['h0023e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00120] =  I38e438ab568822a1c40149a2acc5d876['h00240] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00121] =  I38e438ab568822a1c40149a2acc5d876['h00242] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00122] =  I38e438ab568822a1c40149a2acc5d876['h00244] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00123] =  I38e438ab568822a1c40149a2acc5d876['h00246] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00124] =  I38e438ab568822a1c40149a2acc5d876['h00248] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00125] =  I38e438ab568822a1c40149a2acc5d876['h0024a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00126] =  I38e438ab568822a1c40149a2acc5d876['h0024c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00127] =  I38e438ab568822a1c40149a2acc5d876['h0024e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00128] =  I38e438ab568822a1c40149a2acc5d876['h00250] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00129] =  I38e438ab568822a1c40149a2acc5d876['h00252] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0012a] =  I38e438ab568822a1c40149a2acc5d876['h00254] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0012b] =  I38e438ab568822a1c40149a2acc5d876['h00256] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0012c] =  I38e438ab568822a1c40149a2acc5d876['h00258] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0012d] =  I38e438ab568822a1c40149a2acc5d876['h0025a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0012e] =  I38e438ab568822a1c40149a2acc5d876['h0025c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0012f] =  I38e438ab568822a1c40149a2acc5d876['h0025e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00130] =  I38e438ab568822a1c40149a2acc5d876['h00260] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00131] =  I38e438ab568822a1c40149a2acc5d876['h00262] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00132] =  I38e438ab568822a1c40149a2acc5d876['h00264] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00133] =  I38e438ab568822a1c40149a2acc5d876['h00266] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00134] =  I38e438ab568822a1c40149a2acc5d876['h00268] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00135] =  I38e438ab568822a1c40149a2acc5d876['h0026a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00136] =  I38e438ab568822a1c40149a2acc5d876['h0026c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00137] =  I38e438ab568822a1c40149a2acc5d876['h0026e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00138] =  I38e438ab568822a1c40149a2acc5d876['h00270] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00139] =  I38e438ab568822a1c40149a2acc5d876['h00272] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0013a] =  I38e438ab568822a1c40149a2acc5d876['h00274] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0013b] =  I38e438ab568822a1c40149a2acc5d876['h00276] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0013c] =  I38e438ab568822a1c40149a2acc5d876['h00278] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0013d] =  I38e438ab568822a1c40149a2acc5d876['h0027a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0013e] =  I38e438ab568822a1c40149a2acc5d876['h0027c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0013f] =  I38e438ab568822a1c40149a2acc5d876['h0027e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00140] =  I38e438ab568822a1c40149a2acc5d876['h00280] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00141] =  I38e438ab568822a1c40149a2acc5d876['h00282] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00142] =  I38e438ab568822a1c40149a2acc5d876['h00284] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00143] =  I38e438ab568822a1c40149a2acc5d876['h00286] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00144] =  I38e438ab568822a1c40149a2acc5d876['h00288] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00145] =  I38e438ab568822a1c40149a2acc5d876['h0028a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00146] =  I38e438ab568822a1c40149a2acc5d876['h0028c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00147] =  I38e438ab568822a1c40149a2acc5d876['h0028e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00148] =  I38e438ab568822a1c40149a2acc5d876['h00290] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00149] =  I38e438ab568822a1c40149a2acc5d876['h00292] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0014a] =  I38e438ab568822a1c40149a2acc5d876['h00294] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0014b] =  I38e438ab568822a1c40149a2acc5d876['h00296] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0014c] =  I38e438ab568822a1c40149a2acc5d876['h00298] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0014d] =  I38e438ab568822a1c40149a2acc5d876['h0029a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0014e] =  I38e438ab568822a1c40149a2acc5d876['h0029c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0014f] =  I38e438ab568822a1c40149a2acc5d876['h0029e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00150] =  I38e438ab568822a1c40149a2acc5d876['h002a0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00151] =  I38e438ab568822a1c40149a2acc5d876['h002a2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00152] =  I38e438ab568822a1c40149a2acc5d876['h002a4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00153] =  I38e438ab568822a1c40149a2acc5d876['h002a6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00154] =  I38e438ab568822a1c40149a2acc5d876['h002a8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00155] =  I38e438ab568822a1c40149a2acc5d876['h002aa] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00156] =  I38e438ab568822a1c40149a2acc5d876['h002ac] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00157] =  I38e438ab568822a1c40149a2acc5d876['h002ae] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00158] =  I38e438ab568822a1c40149a2acc5d876['h002b0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00159] =  I38e438ab568822a1c40149a2acc5d876['h002b2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0015a] =  I38e438ab568822a1c40149a2acc5d876['h002b4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0015b] =  I38e438ab568822a1c40149a2acc5d876['h002b6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0015c] =  I38e438ab568822a1c40149a2acc5d876['h002b8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0015d] =  I38e438ab568822a1c40149a2acc5d876['h002ba] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0015e] =  I38e438ab568822a1c40149a2acc5d876['h002bc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0015f] =  I38e438ab568822a1c40149a2acc5d876['h002be] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00160] =  I38e438ab568822a1c40149a2acc5d876['h002c0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00161] =  I38e438ab568822a1c40149a2acc5d876['h002c2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00162] =  I38e438ab568822a1c40149a2acc5d876['h002c4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00163] =  I38e438ab568822a1c40149a2acc5d876['h002c6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00164] =  I38e438ab568822a1c40149a2acc5d876['h002c8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00165] =  I38e438ab568822a1c40149a2acc5d876['h002ca] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00166] =  I38e438ab568822a1c40149a2acc5d876['h002cc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00167] =  I38e438ab568822a1c40149a2acc5d876['h002ce] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00168] =  I38e438ab568822a1c40149a2acc5d876['h002d0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00169] =  I38e438ab568822a1c40149a2acc5d876['h002d2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0016a] =  I38e438ab568822a1c40149a2acc5d876['h002d4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0016b] =  I38e438ab568822a1c40149a2acc5d876['h002d6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0016c] =  I38e438ab568822a1c40149a2acc5d876['h002d8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0016d] =  I38e438ab568822a1c40149a2acc5d876['h002da] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0016e] =  I38e438ab568822a1c40149a2acc5d876['h002dc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0016f] =  I38e438ab568822a1c40149a2acc5d876['h002de] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00170] =  I38e438ab568822a1c40149a2acc5d876['h002e0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00171] =  I38e438ab568822a1c40149a2acc5d876['h002e2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00172] =  I38e438ab568822a1c40149a2acc5d876['h002e4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00173] =  I38e438ab568822a1c40149a2acc5d876['h002e6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00174] =  I38e438ab568822a1c40149a2acc5d876['h002e8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00175] =  I38e438ab568822a1c40149a2acc5d876['h002ea] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00176] =  I38e438ab568822a1c40149a2acc5d876['h002ec] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00177] =  I38e438ab568822a1c40149a2acc5d876['h002ee] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00178] =  I38e438ab568822a1c40149a2acc5d876['h002f0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00179] =  I38e438ab568822a1c40149a2acc5d876['h002f2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0017a] =  I38e438ab568822a1c40149a2acc5d876['h002f4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0017b] =  I38e438ab568822a1c40149a2acc5d876['h002f6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0017c] =  I38e438ab568822a1c40149a2acc5d876['h002f8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0017d] =  I38e438ab568822a1c40149a2acc5d876['h002fa] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0017e] =  I38e438ab568822a1c40149a2acc5d876['h002fc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0017f] =  I38e438ab568822a1c40149a2acc5d876['h002fe] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00180] =  I38e438ab568822a1c40149a2acc5d876['h00300] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00181] =  I38e438ab568822a1c40149a2acc5d876['h00302] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00182] =  I38e438ab568822a1c40149a2acc5d876['h00304] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00183] =  I38e438ab568822a1c40149a2acc5d876['h00306] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00184] =  I38e438ab568822a1c40149a2acc5d876['h00308] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00185] =  I38e438ab568822a1c40149a2acc5d876['h0030a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00186] =  I38e438ab568822a1c40149a2acc5d876['h0030c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00187] =  I38e438ab568822a1c40149a2acc5d876['h0030e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00188] =  I38e438ab568822a1c40149a2acc5d876['h00310] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00189] =  I38e438ab568822a1c40149a2acc5d876['h00312] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0018a] =  I38e438ab568822a1c40149a2acc5d876['h00314] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0018b] =  I38e438ab568822a1c40149a2acc5d876['h00316] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0018c] =  I38e438ab568822a1c40149a2acc5d876['h00318] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0018d] =  I38e438ab568822a1c40149a2acc5d876['h0031a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0018e] =  I38e438ab568822a1c40149a2acc5d876['h0031c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0018f] =  I38e438ab568822a1c40149a2acc5d876['h0031e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00190] =  I38e438ab568822a1c40149a2acc5d876['h00320] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00191] =  I38e438ab568822a1c40149a2acc5d876['h00322] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00192] =  I38e438ab568822a1c40149a2acc5d876['h00324] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00193] =  I38e438ab568822a1c40149a2acc5d876['h00326] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00194] =  I38e438ab568822a1c40149a2acc5d876['h00328] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00195] =  I38e438ab568822a1c40149a2acc5d876['h0032a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00196] =  I38e438ab568822a1c40149a2acc5d876['h0032c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00197] =  I38e438ab568822a1c40149a2acc5d876['h0032e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00198] =  I38e438ab568822a1c40149a2acc5d876['h00330] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00199] =  I38e438ab568822a1c40149a2acc5d876['h00332] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0019a] =  I38e438ab568822a1c40149a2acc5d876['h00334] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0019b] =  I38e438ab568822a1c40149a2acc5d876['h00336] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0019c] =  I38e438ab568822a1c40149a2acc5d876['h00338] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0019d] =  I38e438ab568822a1c40149a2acc5d876['h0033a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0019e] =  I38e438ab568822a1c40149a2acc5d876['h0033c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0019f] =  I38e438ab568822a1c40149a2acc5d876['h0033e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001a0] =  I38e438ab568822a1c40149a2acc5d876['h00340] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001a1] =  I38e438ab568822a1c40149a2acc5d876['h00342] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001a2] =  I38e438ab568822a1c40149a2acc5d876['h00344] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001a3] =  I38e438ab568822a1c40149a2acc5d876['h00346] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001a4] =  I38e438ab568822a1c40149a2acc5d876['h00348] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001a5] =  I38e438ab568822a1c40149a2acc5d876['h0034a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001a6] =  I38e438ab568822a1c40149a2acc5d876['h0034c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001a7] =  I38e438ab568822a1c40149a2acc5d876['h0034e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001a8] =  I38e438ab568822a1c40149a2acc5d876['h00350] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001a9] =  I38e438ab568822a1c40149a2acc5d876['h00352] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001aa] =  I38e438ab568822a1c40149a2acc5d876['h00354] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001ab] =  I38e438ab568822a1c40149a2acc5d876['h00356] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001ac] =  I38e438ab568822a1c40149a2acc5d876['h00358] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001ad] =  I38e438ab568822a1c40149a2acc5d876['h0035a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001ae] =  I38e438ab568822a1c40149a2acc5d876['h0035c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001af] =  I38e438ab568822a1c40149a2acc5d876['h0035e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001b0] =  I38e438ab568822a1c40149a2acc5d876['h00360] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001b1] =  I38e438ab568822a1c40149a2acc5d876['h00362] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001b2] =  I38e438ab568822a1c40149a2acc5d876['h00364] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001b3] =  I38e438ab568822a1c40149a2acc5d876['h00366] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001b4] =  I38e438ab568822a1c40149a2acc5d876['h00368] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001b5] =  I38e438ab568822a1c40149a2acc5d876['h0036a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001b6] =  I38e438ab568822a1c40149a2acc5d876['h0036c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001b7] =  I38e438ab568822a1c40149a2acc5d876['h0036e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001b8] =  I38e438ab568822a1c40149a2acc5d876['h00370] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001b9] =  I38e438ab568822a1c40149a2acc5d876['h00372] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001ba] =  I38e438ab568822a1c40149a2acc5d876['h00374] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001bb] =  I38e438ab568822a1c40149a2acc5d876['h00376] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001bc] =  I38e438ab568822a1c40149a2acc5d876['h00378] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001bd] =  I38e438ab568822a1c40149a2acc5d876['h0037a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001be] =  I38e438ab568822a1c40149a2acc5d876['h0037c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001bf] =  I38e438ab568822a1c40149a2acc5d876['h0037e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001c0] =  I38e438ab568822a1c40149a2acc5d876['h00380] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001c1] =  I38e438ab568822a1c40149a2acc5d876['h00382] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001c2] =  I38e438ab568822a1c40149a2acc5d876['h00384] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001c3] =  I38e438ab568822a1c40149a2acc5d876['h00386] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001c4] =  I38e438ab568822a1c40149a2acc5d876['h00388] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001c5] =  I38e438ab568822a1c40149a2acc5d876['h0038a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001c6] =  I38e438ab568822a1c40149a2acc5d876['h0038c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001c7] =  I38e438ab568822a1c40149a2acc5d876['h0038e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001c8] =  I38e438ab568822a1c40149a2acc5d876['h00390] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001c9] =  I38e438ab568822a1c40149a2acc5d876['h00392] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001ca] =  I38e438ab568822a1c40149a2acc5d876['h00394] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001cb] =  I38e438ab568822a1c40149a2acc5d876['h00396] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001cc] =  I38e438ab568822a1c40149a2acc5d876['h00398] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001cd] =  I38e438ab568822a1c40149a2acc5d876['h0039a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001ce] =  I38e438ab568822a1c40149a2acc5d876['h0039c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001cf] =  I38e438ab568822a1c40149a2acc5d876['h0039e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001d0] =  I38e438ab568822a1c40149a2acc5d876['h003a0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001d1] =  I38e438ab568822a1c40149a2acc5d876['h003a2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001d2] =  I38e438ab568822a1c40149a2acc5d876['h003a4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001d3] =  I38e438ab568822a1c40149a2acc5d876['h003a6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001d4] =  I38e438ab568822a1c40149a2acc5d876['h003a8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001d5] =  I38e438ab568822a1c40149a2acc5d876['h003aa] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001d6] =  I38e438ab568822a1c40149a2acc5d876['h003ac] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001d7] =  I38e438ab568822a1c40149a2acc5d876['h003ae] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001d8] =  I38e438ab568822a1c40149a2acc5d876['h003b0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001d9] =  I38e438ab568822a1c40149a2acc5d876['h003b2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001da] =  I38e438ab568822a1c40149a2acc5d876['h003b4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001db] =  I38e438ab568822a1c40149a2acc5d876['h003b6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001dc] =  I38e438ab568822a1c40149a2acc5d876['h003b8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001dd] =  I38e438ab568822a1c40149a2acc5d876['h003ba] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001de] =  I38e438ab568822a1c40149a2acc5d876['h003bc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001df] =  I38e438ab568822a1c40149a2acc5d876['h003be] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001e0] =  I38e438ab568822a1c40149a2acc5d876['h003c0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001e1] =  I38e438ab568822a1c40149a2acc5d876['h003c2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001e2] =  I38e438ab568822a1c40149a2acc5d876['h003c4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001e3] =  I38e438ab568822a1c40149a2acc5d876['h003c6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001e4] =  I38e438ab568822a1c40149a2acc5d876['h003c8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001e5] =  I38e438ab568822a1c40149a2acc5d876['h003ca] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001e6] =  I38e438ab568822a1c40149a2acc5d876['h003cc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001e7] =  I38e438ab568822a1c40149a2acc5d876['h003ce] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001e8] =  I38e438ab568822a1c40149a2acc5d876['h003d0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001e9] =  I38e438ab568822a1c40149a2acc5d876['h003d2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001ea] =  I38e438ab568822a1c40149a2acc5d876['h003d4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001eb] =  I38e438ab568822a1c40149a2acc5d876['h003d6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001ec] =  I38e438ab568822a1c40149a2acc5d876['h003d8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001ed] =  I38e438ab568822a1c40149a2acc5d876['h003da] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001ee] =  I38e438ab568822a1c40149a2acc5d876['h003dc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001ef] =  I38e438ab568822a1c40149a2acc5d876['h003de] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001f0] =  I38e438ab568822a1c40149a2acc5d876['h003e0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001f1] =  I38e438ab568822a1c40149a2acc5d876['h003e2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001f2] =  I38e438ab568822a1c40149a2acc5d876['h003e4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001f3] =  I38e438ab568822a1c40149a2acc5d876['h003e6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001f4] =  I38e438ab568822a1c40149a2acc5d876['h003e8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001f5] =  I38e438ab568822a1c40149a2acc5d876['h003ea] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001f6] =  I38e438ab568822a1c40149a2acc5d876['h003ec] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001f7] =  I38e438ab568822a1c40149a2acc5d876['h003ee] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001f8] =  I38e438ab568822a1c40149a2acc5d876['h003f0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001f9] =  I38e438ab568822a1c40149a2acc5d876['h003f2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001fa] =  I38e438ab568822a1c40149a2acc5d876['h003f4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001fb] =  I38e438ab568822a1c40149a2acc5d876['h003f6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001fc] =  I38e438ab568822a1c40149a2acc5d876['h003f8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001fd] =  I38e438ab568822a1c40149a2acc5d876['h003fa] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001fe] =  I38e438ab568822a1c40149a2acc5d876['h003fc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h001ff] =  I38e438ab568822a1c40149a2acc5d876['h003fe] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00200] =  I38e438ab568822a1c40149a2acc5d876['h00400] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00201] =  I38e438ab568822a1c40149a2acc5d876['h00402] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00202] =  I38e438ab568822a1c40149a2acc5d876['h00404] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00203] =  I38e438ab568822a1c40149a2acc5d876['h00406] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00204] =  I38e438ab568822a1c40149a2acc5d876['h00408] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00205] =  I38e438ab568822a1c40149a2acc5d876['h0040a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00206] =  I38e438ab568822a1c40149a2acc5d876['h0040c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00207] =  I38e438ab568822a1c40149a2acc5d876['h0040e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00208] =  I38e438ab568822a1c40149a2acc5d876['h00410] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00209] =  I38e438ab568822a1c40149a2acc5d876['h00412] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0020a] =  I38e438ab568822a1c40149a2acc5d876['h00414] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0020b] =  I38e438ab568822a1c40149a2acc5d876['h00416] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0020c] =  I38e438ab568822a1c40149a2acc5d876['h00418] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0020d] =  I38e438ab568822a1c40149a2acc5d876['h0041a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0020e] =  I38e438ab568822a1c40149a2acc5d876['h0041c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0020f] =  I38e438ab568822a1c40149a2acc5d876['h0041e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00210] =  I38e438ab568822a1c40149a2acc5d876['h00420] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00211] =  I38e438ab568822a1c40149a2acc5d876['h00422] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00212] =  I38e438ab568822a1c40149a2acc5d876['h00424] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00213] =  I38e438ab568822a1c40149a2acc5d876['h00426] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00214] =  I38e438ab568822a1c40149a2acc5d876['h00428] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00215] =  I38e438ab568822a1c40149a2acc5d876['h0042a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00216] =  I38e438ab568822a1c40149a2acc5d876['h0042c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00217] =  I38e438ab568822a1c40149a2acc5d876['h0042e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00218] =  I38e438ab568822a1c40149a2acc5d876['h00430] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00219] =  I38e438ab568822a1c40149a2acc5d876['h00432] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0021a] =  I38e438ab568822a1c40149a2acc5d876['h00434] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0021b] =  I38e438ab568822a1c40149a2acc5d876['h00436] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0021c] =  I38e438ab568822a1c40149a2acc5d876['h00438] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0021d] =  I38e438ab568822a1c40149a2acc5d876['h0043a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0021e] =  I38e438ab568822a1c40149a2acc5d876['h0043c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0021f] =  I38e438ab568822a1c40149a2acc5d876['h0043e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00220] =  I38e438ab568822a1c40149a2acc5d876['h00440] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00221] =  I38e438ab568822a1c40149a2acc5d876['h00442] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00222] =  I38e438ab568822a1c40149a2acc5d876['h00444] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00223] =  I38e438ab568822a1c40149a2acc5d876['h00446] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00224] =  I38e438ab568822a1c40149a2acc5d876['h00448] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00225] =  I38e438ab568822a1c40149a2acc5d876['h0044a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00226] =  I38e438ab568822a1c40149a2acc5d876['h0044c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00227] =  I38e438ab568822a1c40149a2acc5d876['h0044e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00228] =  I38e438ab568822a1c40149a2acc5d876['h00450] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00229] =  I38e438ab568822a1c40149a2acc5d876['h00452] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0022a] =  I38e438ab568822a1c40149a2acc5d876['h00454] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0022b] =  I38e438ab568822a1c40149a2acc5d876['h00456] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0022c] =  I38e438ab568822a1c40149a2acc5d876['h00458] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0022d] =  I38e438ab568822a1c40149a2acc5d876['h0045a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0022e] =  I38e438ab568822a1c40149a2acc5d876['h0045c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0022f] =  I38e438ab568822a1c40149a2acc5d876['h0045e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00230] =  I38e438ab568822a1c40149a2acc5d876['h00460] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00231] =  I38e438ab568822a1c40149a2acc5d876['h00462] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00232] =  I38e438ab568822a1c40149a2acc5d876['h00464] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00233] =  I38e438ab568822a1c40149a2acc5d876['h00466] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00234] =  I38e438ab568822a1c40149a2acc5d876['h00468] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00235] =  I38e438ab568822a1c40149a2acc5d876['h0046a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00236] =  I38e438ab568822a1c40149a2acc5d876['h0046c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00237] =  I38e438ab568822a1c40149a2acc5d876['h0046e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00238] =  I38e438ab568822a1c40149a2acc5d876['h00470] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00239] =  I38e438ab568822a1c40149a2acc5d876['h00472] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0023a] =  I38e438ab568822a1c40149a2acc5d876['h00474] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0023b] =  I38e438ab568822a1c40149a2acc5d876['h00476] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0023c] =  I38e438ab568822a1c40149a2acc5d876['h00478] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0023d] =  I38e438ab568822a1c40149a2acc5d876['h0047a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0023e] =  I38e438ab568822a1c40149a2acc5d876['h0047c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0023f] =  I38e438ab568822a1c40149a2acc5d876['h0047e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00240] =  I38e438ab568822a1c40149a2acc5d876['h00480] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00241] =  I38e438ab568822a1c40149a2acc5d876['h00482] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00242] =  I38e438ab568822a1c40149a2acc5d876['h00484] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00243] =  I38e438ab568822a1c40149a2acc5d876['h00486] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00244] =  I38e438ab568822a1c40149a2acc5d876['h00488] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00245] =  I38e438ab568822a1c40149a2acc5d876['h0048a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00246] =  I38e438ab568822a1c40149a2acc5d876['h0048c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00247] =  I38e438ab568822a1c40149a2acc5d876['h0048e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00248] =  I38e438ab568822a1c40149a2acc5d876['h00490] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00249] =  I38e438ab568822a1c40149a2acc5d876['h00492] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0024a] =  I38e438ab568822a1c40149a2acc5d876['h00494] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0024b] =  I38e438ab568822a1c40149a2acc5d876['h00496] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0024c] =  I38e438ab568822a1c40149a2acc5d876['h00498] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0024d] =  I38e438ab568822a1c40149a2acc5d876['h0049a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0024e] =  I38e438ab568822a1c40149a2acc5d876['h0049c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0024f] =  I38e438ab568822a1c40149a2acc5d876['h0049e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00250] =  I38e438ab568822a1c40149a2acc5d876['h004a0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00251] =  I38e438ab568822a1c40149a2acc5d876['h004a2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00252] =  I38e438ab568822a1c40149a2acc5d876['h004a4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00253] =  I38e438ab568822a1c40149a2acc5d876['h004a6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00254] =  I38e438ab568822a1c40149a2acc5d876['h004a8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00255] =  I38e438ab568822a1c40149a2acc5d876['h004aa] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00256] =  I38e438ab568822a1c40149a2acc5d876['h004ac] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00257] =  I38e438ab568822a1c40149a2acc5d876['h004ae] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00258] =  I38e438ab568822a1c40149a2acc5d876['h004b0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00259] =  I38e438ab568822a1c40149a2acc5d876['h004b2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0025a] =  I38e438ab568822a1c40149a2acc5d876['h004b4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0025b] =  I38e438ab568822a1c40149a2acc5d876['h004b6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0025c] =  I38e438ab568822a1c40149a2acc5d876['h004b8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0025d] =  I38e438ab568822a1c40149a2acc5d876['h004ba] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0025e] =  I38e438ab568822a1c40149a2acc5d876['h004bc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0025f] =  I38e438ab568822a1c40149a2acc5d876['h004be] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00260] =  I38e438ab568822a1c40149a2acc5d876['h004c0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00261] =  I38e438ab568822a1c40149a2acc5d876['h004c2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00262] =  I38e438ab568822a1c40149a2acc5d876['h004c4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00263] =  I38e438ab568822a1c40149a2acc5d876['h004c6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00264] =  I38e438ab568822a1c40149a2acc5d876['h004c8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00265] =  I38e438ab568822a1c40149a2acc5d876['h004ca] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00266] =  I38e438ab568822a1c40149a2acc5d876['h004cc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00267] =  I38e438ab568822a1c40149a2acc5d876['h004ce] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00268] =  I38e438ab568822a1c40149a2acc5d876['h004d0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00269] =  I38e438ab568822a1c40149a2acc5d876['h004d2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0026a] =  I38e438ab568822a1c40149a2acc5d876['h004d4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0026b] =  I38e438ab568822a1c40149a2acc5d876['h004d6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0026c] =  I38e438ab568822a1c40149a2acc5d876['h004d8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0026d] =  I38e438ab568822a1c40149a2acc5d876['h004da] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0026e] =  I38e438ab568822a1c40149a2acc5d876['h004dc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0026f] =  I38e438ab568822a1c40149a2acc5d876['h004de] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00270] =  I38e438ab568822a1c40149a2acc5d876['h004e0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00271] =  I38e438ab568822a1c40149a2acc5d876['h004e2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00272] =  I38e438ab568822a1c40149a2acc5d876['h004e4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00273] =  I38e438ab568822a1c40149a2acc5d876['h004e6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00274] =  I38e438ab568822a1c40149a2acc5d876['h004e8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00275] =  I38e438ab568822a1c40149a2acc5d876['h004ea] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00276] =  I38e438ab568822a1c40149a2acc5d876['h004ec] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00277] =  I38e438ab568822a1c40149a2acc5d876['h004ee] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00278] =  I38e438ab568822a1c40149a2acc5d876['h004f0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00279] =  I38e438ab568822a1c40149a2acc5d876['h004f2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0027a] =  I38e438ab568822a1c40149a2acc5d876['h004f4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0027b] =  I38e438ab568822a1c40149a2acc5d876['h004f6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0027c] =  I38e438ab568822a1c40149a2acc5d876['h004f8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0027d] =  I38e438ab568822a1c40149a2acc5d876['h004fa] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0027e] =  I38e438ab568822a1c40149a2acc5d876['h004fc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0027f] =  I38e438ab568822a1c40149a2acc5d876['h004fe] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00280] =  I38e438ab568822a1c40149a2acc5d876['h00500] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00281] =  I38e438ab568822a1c40149a2acc5d876['h00502] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00282] =  I38e438ab568822a1c40149a2acc5d876['h00504] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00283] =  I38e438ab568822a1c40149a2acc5d876['h00506] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00284] =  I38e438ab568822a1c40149a2acc5d876['h00508] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00285] =  I38e438ab568822a1c40149a2acc5d876['h0050a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00286] =  I38e438ab568822a1c40149a2acc5d876['h0050c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00287] =  I38e438ab568822a1c40149a2acc5d876['h0050e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00288] =  I38e438ab568822a1c40149a2acc5d876['h00510] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00289] =  I38e438ab568822a1c40149a2acc5d876['h00512] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0028a] =  I38e438ab568822a1c40149a2acc5d876['h00514] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0028b] =  I38e438ab568822a1c40149a2acc5d876['h00516] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0028c] =  I38e438ab568822a1c40149a2acc5d876['h00518] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0028d] =  I38e438ab568822a1c40149a2acc5d876['h0051a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0028e] =  I38e438ab568822a1c40149a2acc5d876['h0051c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0028f] =  I38e438ab568822a1c40149a2acc5d876['h0051e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00290] =  I38e438ab568822a1c40149a2acc5d876['h00520] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00291] =  I38e438ab568822a1c40149a2acc5d876['h00522] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00292] =  I38e438ab568822a1c40149a2acc5d876['h00524] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00293] =  I38e438ab568822a1c40149a2acc5d876['h00526] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00294] =  I38e438ab568822a1c40149a2acc5d876['h00528] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00295] =  I38e438ab568822a1c40149a2acc5d876['h0052a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00296] =  I38e438ab568822a1c40149a2acc5d876['h0052c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00297] =  I38e438ab568822a1c40149a2acc5d876['h0052e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00298] =  I38e438ab568822a1c40149a2acc5d876['h00530] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00299] =  I38e438ab568822a1c40149a2acc5d876['h00532] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0029a] =  I38e438ab568822a1c40149a2acc5d876['h00534] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0029b] =  I38e438ab568822a1c40149a2acc5d876['h00536] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0029c] =  I38e438ab568822a1c40149a2acc5d876['h00538] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0029d] =  I38e438ab568822a1c40149a2acc5d876['h0053a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0029e] =  I38e438ab568822a1c40149a2acc5d876['h0053c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0029f] =  I38e438ab568822a1c40149a2acc5d876['h0053e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002a0] =  I38e438ab568822a1c40149a2acc5d876['h00540] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002a1] =  I38e438ab568822a1c40149a2acc5d876['h00542] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002a2] =  I38e438ab568822a1c40149a2acc5d876['h00544] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002a3] =  I38e438ab568822a1c40149a2acc5d876['h00546] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002a4] =  I38e438ab568822a1c40149a2acc5d876['h00548] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002a5] =  I38e438ab568822a1c40149a2acc5d876['h0054a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002a6] =  I38e438ab568822a1c40149a2acc5d876['h0054c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002a7] =  I38e438ab568822a1c40149a2acc5d876['h0054e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002a8] =  I38e438ab568822a1c40149a2acc5d876['h00550] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002a9] =  I38e438ab568822a1c40149a2acc5d876['h00552] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002aa] =  I38e438ab568822a1c40149a2acc5d876['h00554] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002ab] =  I38e438ab568822a1c40149a2acc5d876['h00556] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002ac] =  I38e438ab568822a1c40149a2acc5d876['h00558] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002ad] =  I38e438ab568822a1c40149a2acc5d876['h0055a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002ae] =  I38e438ab568822a1c40149a2acc5d876['h0055c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002af] =  I38e438ab568822a1c40149a2acc5d876['h0055e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002b0] =  I38e438ab568822a1c40149a2acc5d876['h00560] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002b1] =  I38e438ab568822a1c40149a2acc5d876['h00562] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002b2] =  I38e438ab568822a1c40149a2acc5d876['h00564] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002b3] =  I38e438ab568822a1c40149a2acc5d876['h00566] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002b4] =  I38e438ab568822a1c40149a2acc5d876['h00568] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002b5] =  I38e438ab568822a1c40149a2acc5d876['h0056a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002b6] =  I38e438ab568822a1c40149a2acc5d876['h0056c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002b7] =  I38e438ab568822a1c40149a2acc5d876['h0056e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002b8] =  I38e438ab568822a1c40149a2acc5d876['h00570] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002b9] =  I38e438ab568822a1c40149a2acc5d876['h00572] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002ba] =  I38e438ab568822a1c40149a2acc5d876['h00574] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002bb] =  I38e438ab568822a1c40149a2acc5d876['h00576] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002bc] =  I38e438ab568822a1c40149a2acc5d876['h00578] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002bd] =  I38e438ab568822a1c40149a2acc5d876['h0057a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002be] =  I38e438ab568822a1c40149a2acc5d876['h0057c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002bf] =  I38e438ab568822a1c40149a2acc5d876['h0057e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002c0] =  I38e438ab568822a1c40149a2acc5d876['h00580] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002c1] =  I38e438ab568822a1c40149a2acc5d876['h00582] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002c2] =  I38e438ab568822a1c40149a2acc5d876['h00584] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002c3] =  I38e438ab568822a1c40149a2acc5d876['h00586] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002c4] =  I38e438ab568822a1c40149a2acc5d876['h00588] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002c5] =  I38e438ab568822a1c40149a2acc5d876['h0058a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002c6] =  I38e438ab568822a1c40149a2acc5d876['h0058c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002c7] =  I38e438ab568822a1c40149a2acc5d876['h0058e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002c8] =  I38e438ab568822a1c40149a2acc5d876['h00590] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002c9] =  I38e438ab568822a1c40149a2acc5d876['h00592] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002ca] =  I38e438ab568822a1c40149a2acc5d876['h00594] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002cb] =  I38e438ab568822a1c40149a2acc5d876['h00596] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002cc] =  I38e438ab568822a1c40149a2acc5d876['h00598] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002cd] =  I38e438ab568822a1c40149a2acc5d876['h0059a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002ce] =  I38e438ab568822a1c40149a2acc5d876['h0059c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002cf] =  I38e438ab568822a1c40149a2acc5d876['h0059e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002d0] =  I38e438ab568822a1c40149a2acc5d876['h005a0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002d1] =  I38e438ab568822a1c40149a2acc5d876['h005a2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002d2] =  I38e438ab568822a1c40149a2acc5d876['h005a4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002d3] =  I38e438ab568822a1c40149a2acc5d876['h005a6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002d4] =  I38e438ab568822a1c40149a2acc5d876['h005a8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002d5] =  I38e438ab568822a1c40149a2acc5d876['h005aa] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002d6] =  I38e438ab568822a1c40149a2acc5d876['h005ac] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002d7] =  I38e438ab568822a1c40149a2acc5d876['h005ae] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002d8] =  I38e438ab568822a1c40149a2acc5d876['h005b0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002d9] =  I38e438ab568822a1c40149a2acc5d876['h005b2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002da] =  I38e438ab568822a1c40149a2acc5d876['h005b4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002db] =  I38e438ab568822a1c40149a2acc5d876['h005b6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002dc] =  I38e438ab568822a1c40149a2acc5d876['h005b8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002dd] =  I38e438ab568822a1c40149a2acc5d876['h005ba] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002de] =  I38e438ab568822a1c40149a2acc5d876['h005bc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002df] =  I38e438ab568822a1c40149a2acc5d876['h005be] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002e0] =  I38e438ab568822a1c40149a2acc5d876['h005c0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002e1] =  I38e438ab568822a1c40149a2acc5d876['h005c2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002e2] =  I38e438ab568822a1c40149a2acc5d876['h005c4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002e3] =  I38e438ab568822a1c40149a2acc5d876['h005c6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002e4] =  I38e438ab568822a1c40149a2acc5d876['h005c8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002e5] =  I38e438ab568822a1c40149a2acc5d876['h005ca] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002e6] =  I38e438ab568822a1c40149a2acc5d876['h005cc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002e7] =  I38e438ab568822a1c40149a2acc5d876['h005ce] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002e8] =  I38e438ab568822a1c40149a2acc5d876['h005d0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002e9] =  I38e438ab568822a1c40149a2acc5d876['h005d2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002ea] =  I38e438ab568822a1c40149a2acc5d876['h005d4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002eb] =  I38e438ab568822a1c40149a2acc5d876['h005d6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002ec] =  I38e438ab568822a1c40149a2acc5d876['h005d8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002ed] =  I38e438ab568822a1c40149a2acc5d876['h005da] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002ee] =  I38e438ab568822a1c40149a2acc5d876['h005dc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002ef] =  I38e438ab568822a1c40149a2acc5d876['h005de] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002f0] =  I38e438ab568822a1c40149a2acc5d876['h005e0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002f1] =  I38e438ab568822a1c40149a2acc5d876['h005e2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002f2] =  I38e438ab568822a1c40149a2acc5d876['h005e4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002f3] =  I38e438ab568822a1c40149a2acc5d876['h005e6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002f4] =  I38e438ab568822a1c40149a2acc5d876['h005e8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002f5] =  I38e438ab568822a1c40149a2acc5d876['h005ea] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002f6] =  I38e438ab568822a1c40149a2acc5d876['h005ec] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002f7] =  I38e438ab568822a1c40149a2acc5d876['h005ee] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002f8] =  I38e438ab568822a1c40149a2acc5d876['h005f0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002f9] =  I38e438ab568822a1c40149a2acc5d876['h005f2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002fa] =  I38e438ab568822a1c40149a2acc5d876['h005f4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002fb] =  I38e438ab568822a1c40149a2acc5d876['h005f6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002fc] =  I38e438ab568822a1c40149a2acc5d876['h005f8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002fd] =  I38e438ab568822a1c40149a2acc5d876['h005fa] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002fe] =  I38e438ab568822a1c40149a2acc5d876['h005fc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h002ff] =  I38e438ab568822a1c40149a2acc5d876['h005fe] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00300] =  I38e438ab568822a1c40149a2acc5d876['h00600] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00301] =  I38e438ab568822a1c40149a2acc5d876['h00602] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00302] =  I38e438ab568822a1c40149a2acc5d876['h00604] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00303] =  I38e438ab568822a1c40149a2acc5d876['h00606] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00304] =  I38e438ab568822a1c40149a2acc5d876['h00608] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00305] =  I38e438ab568822a1c40149a2acc5d876['h0060a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00306] =  I38e438ab568822a1c40149a2acc5d876['h0060c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00307] =  I38e438ab568822a1c40149a2acc5d876['h0060e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00308] =  I38e438ab568822a1c40149a2acc5d876['h00610] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00309] =  I38e438ab568822a1c40149a2acc5d876['h00612] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0030a] =  I38e438ab568822a1c40149a2acc5d876['h00614] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0030b] =  I38e438ab568822a1c40149a2acc5d876['h00616] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0030c] =  I38e438ab568822a1c40149a2acc5d876['h00618] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0030d] =  I38e438ab568822a1c40149a2acc5d876['h0061a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0030e] =  I38e438ab568822a1c40149a2acc5d876['h0061c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0030f] =  I38e438ab568822a1c40149a2acc5d876['h0061e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00310] =  I38e438ab568822a1c40149a2acc5d876['h00620] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00311] =  I38e438ab568822a1c40149a2acc5d876['h00622] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00312] =  I38e438ab568822a1c40149a2acc5d876['h00624] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00313] =  I38e438ab568822a1c40149a2acc5d876['h00626] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00314] =  I38e438ab568822a1c40149a2acc5d876['h00628] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00315] =  I38e438ab568822a1c40149a2acc5d876['h0062a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00316] =  I38e438ab568822a1c40149a2acc5d876['h0062c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00317] =  I38e438ab568822a1c40149a2acc5d876['h0062e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00318] =  I38e438ab568822a1c40149a2acc5d876['h00630] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00319] =  I38e438ab568822a1c40149a2acc5d876['h00632] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0031a] =  I38e438ab568822a1c40149a2acc5d876['h00634] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0031b] =  I38e438ab568822a1c40149a2acc5d876['h00636] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0031c] =  I38e438ab568822a1c40149a2acc5d876['h00638] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0031d] =  I38e438ab568822a1c40149a2acc5d876['h0063a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0031e] =  I38e438ab568822a1c40149a2acc5d876['h0063c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0031f] =  I38e438ab568822a1c40149a2acc5d876['h0063e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00320] =  I38e438ab568822a1c40149a2acc5d876['h00640] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00321] =  I38e438ab568822a1c40149a2acc5d876['h00642] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00322] =  I38e438ab568822a1c40149a2acc5d876['h00644] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00323] =  I38e438ab568822a1c40149a2acc5d876['h00646] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00324] =  I38e438ab568822a1c40149a2acc5d876['h00648] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00325] =  I38e438ab568822a1c40149a2acc5d876['h0064a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00326] =  I38e438ab568822a1c40149a2acc5d876['h0064c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00327] =  I38e438ab568822a1c40149a2acc5d876['h0064e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00328] =  I38e438ab568822a1c40149a2acc5d876['h00650] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00329] =  I38e438ab568822a1c40149a2acc5d876['h00652] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0032a] =  I38e438ab568822a1c40149a2acc5d876['h00654] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0032b] =  I38e438ab568822a1c40149a2acc5d876['h00656] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0032c] =  I38e438ab568822a1c40149a2acc5d876['h00658] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0032d] =  I38e438ab568822a1c40149a2acc5d876['h0065a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0032e] =  I38e438ab568822a1c40149a2acc5d876['h0065c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0032f] =  I38e438ab568822a1c40149a2acc5d876['h0065e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00330] =  I38e438ab568822a1c40149a2acc5d876['h00660] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00331] =  I38e438ab568822a1c40149a2acc5d876['h00662] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00332] =  I38e438ab568822a1c40149a2acc5d876['h00664] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00333] =  I38e438ab568822a1c40149a2acc5d876['h00666] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00334] =  I38e438ab568822a1c40149a2acc5d876['h00668] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00335] =  I38e438ab568822a1c40149a2acc5d876['h0066a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00336] =  I38e438ab568822a1c40149a2acc5d876['h0066c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00337] =  I38e438ab568822a1c40149a2acc5d876['h0066e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00338] =  I38e438ab568822a1c40149a2acc5d876['h00670] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00339] =  I38e438ab568822a1c40149a2acc5d876['h00672] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0033a] =  I38e438ab568822a1c40149a2acc5d876['h00674] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0033b] =  I38e438ab568822a1c40149a2acc5d876['h00676] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0033c] =  I38e438ab568822a1c40149a2acc5d876['h00678] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0033d] =  I38e438ab568822a1c40149a2acc5d876['h0067a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0033e] =  I38e438ab568822a1c40149a2acc5d876['h0067c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0033f] =  I38e438ab568822a1c40149a2acc5d876['h0067e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00340] =  I38e438ab568822a1c40149a2acc5d876['h00680] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00341] =  I38e438ab568822a1c40149a2acc5d876['h00682] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00342] =  I38e438ab568822a1c40149a2acc5d876['h00684] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00343] =  I38e438ab568822a1c40149a2acc5d876['h00686] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00344] =  I38e438ab568822a1c40149a2acc5d876['h00688] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00345] =  I38e438ab568822a1c40149a2acc5d876['h0068a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00346] =  I38e438ab568822a1c40149a2acc5d876['h0068c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00347] =  I38e438ab568822a1c40149a2acc5d876['h0068e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00348] =  I38e438ab568822a1c40149a2acc5d876['h00690] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00349] =  I38e438ab568822a1c40149a2acc5d876['h00692] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0034a] =  I38e438ab568822a1c40149a2acc5d876['h00694] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0034b] =  I38e438ab568822a1c40149a2acc5d876['h00696] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0034c] =  I38e438ab568822a1c40149a2acc5d876['h00698] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0034d] =  I38e438ab568822a1c40149a2acc5d876['h0069a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0034e] =  I38e438ab568822a1c40149a2acc5d876['h0069c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0034f] =  I38e438ab568822a1c40149a2acc5d876['h0069e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00350] =  I38e438ab568822a1c40149a2acc5d876['h006a0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00351] =  I38e438ab568822a1c40149a2acc5d876['h006a2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00352] =  I38e438ab568822a1c40149a2acc5d876['h006a4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00353] =  I38e438ab568822a1c40149a2acc5d876['h006a6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00354] =  I38e438ab568822a1c40149a2acc5d876['h006a8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00355] =  I38e438ab568822a1c40149a2acc5d876['h006aa] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00356] =  I38e438ab568822a1c40149a2acc5d876['h006ac] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00357] =  I38e438ab568822a1c40149a2acc5d876['h006ae] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00358] =  I38e438ab568822a1c40149a2acc5d876['h006b0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00359] =  I38e438ab568822a1c40149a2acc5d876['h006b2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0035a] =  I38e438ab568822a1c40149a2acc5d876['h006b4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0035b] =  I38e438ab568822a1c40149a2acc5d876['h006b6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0035c] =  I38e438ab568822a1c40149a2acc5d876['h006b8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0035d] =  I38e438ab568822a1c40149a2acc5d876['h006ba] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0035e] =  I38e438ab568822a1c40149a2acc5d876['h006bc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0035f] =  I38e438ab568822a1c40149a2acc5d876['h006be] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00360] =  I38e438ab568822a1c40149a2acc5d876['h006c0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00361] =  I38e438ab568822a1c40149a2acc5d876['h006c2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00362] =  I38e438ab568822a1c40149a2acc5d876['h006c4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00363] =  I38e438ab568822a1c40149a2acc5d876['h006c6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00364] =  I38e438ab568822a1c40149a2acc5d876['h006c8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00365] =  I38e438ab568822a1c40149a2acc5d876['h006ca] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00366] =  I38e438ab568822a1c40149a2acc5d876['h006cc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00367] =  I38e438ab568822a1c40149a2acc5d876['h006ce] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00368] =  I38e438ab568822a1c40149a2acc5d876['h006d0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00369] =  I38e438ab568822a1c40149a2acc5d876['h006d2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0036a] =  I38e438ab568822a1c40149a2acc5d876['h006d4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0036b] =  I38e438ab568822a1c40149a2acc5d876['h006d6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0036c] =  I38e438ab568822a1c40149a2acc5d876['h006d8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0036d] =  I38e438ab568822a1c40149a2acc5d876['h006da] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0036e] =  I38e438ab568822a1c40149a2acc5d876['h006dc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0036f] =  I38e438ab568822a1c40149a2acc5d876['h006de] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00370] =  I38e438ab568822a1c40149a2acc5d876['h006e0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00371] =  I38e438ab568822a1c40149a2acc5d876['h006e2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00372] =  I38e438ab568822a1c40149a2acc5d876['h006e4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00373] =  I38e438ab568822a1c40149a2acc5d876['h006e6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00374] =  I38e438ab568822a1c40149a2acc5d876['h006e8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00375] =  I38e438ab568822a1c40149a2acc5d876['h006ea] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00376] =  I38e438ab568822a1c40149a2acc5d876['h006ec] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00377] =  I38e438ab568822a1c40149a2acc5d876['h006ee] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00378] =  I38e438ab568822a1c40149a2acc5d876['h006f0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00379] =  I38e438ab568822a1c40149a2acc5d876['h006f2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0037a] =  I38e438ab568822a1c40149a2acc5d876['h006f4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0037b] =  I38e438ab568822a1c40149a2acc5d876['h006f6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0037c] =  I38e438ab568822a1c40149a2acc5d876['h006f8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0037d] =  I38e438ab568822a1c40149a2acc5d876['h006fa] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0037e] =  I38e438ab568822a1c40149a2acc5d876['h006fc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0037f] =  I38e438ab568822a1c40149a2acc5d876['h006fe] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00380] =  I38e438ab568822a1c40149a2acc5d876['h00700] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00381] =  I38e438ab568822a1c40149a2acc5d876['h00702] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00382] =  I38e438ab568822a1c40149a2acc5d876['h00704] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00383] =  I38e438ab568822a1c40149a2acc5d876['h00706] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00384] =  I38e438ab568822a1c40149a2acc5d876['h00708] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00385] =  I38e438ab568822a1c40149a2acc5d876['h0070a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00386] =  I38e438ab568822a1c40149a2acc5d876['h0070c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00387] =  I38e438ab568822a1c40149a2acc5d876['h0070e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00388] =  I38e438ab568822a1c40149a2acc5d876['h00710] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00389] =  I38e438ab568822a1c40149a2acc5d876['h00712] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0038a] =  I38e438ab568822a1c40149a2acc5d876['h00714] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0038b] =  I38e438ab568822a1c40149a2acc5d876['h00716] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0038c] =  I38e438ab568822a1c40149a2acc5d876['h00718] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0038d] =  I38e438ab568822a1c40149a2acc5d876['h0071a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0038e] =  I38e438ab568822a1c40149a2acc5d876['h0071c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0038f] =  I38e438ab568822a1c40149a2acc5d876['h0071e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00390] =  I38e438ab568822a1c40149a2acc5d876['h00720] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00391] =  I38e438ab568822a1c40149a2acc5d876['h00722] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00392] =  I38e438ab568822a1c40149a2acc5d876['h00724] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00393] =  I38e438ab568822a1c40149a2acc5d876['h00726] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00394] =  I38e438ab568822a1c40149a2acc5d876['h00728] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00395] =  I38e438ab568822a1c40149a2acc5d876['h0072a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00396] =  I38e438ab568822a1c40149a2acc5d876['h0072c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00397] =  I38e438ab568822a1c40149a2acc5d876['h0072e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00398] =  I38e438ab568822a1c40149a2acc5d876['h00730] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h00399] =  I38e438ab568822a1c40149a2acc5d876['h00732] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0039a] =  I38e438ab568822a1c40149a2acc5d876['h00734] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0039b] =  I38e438ab568822a1c40149a2acc5d876['h00736] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0039c] =  I38e438ab568822a1c40149a2acc5d876['h00738] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0039d] =  I38e438ab568822a1c40149a2acc5d876['h0073a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0039e] =  I38e438ab568822a1c40149a2acc5d876['h0073c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h0039f] =  I38e438ab568822a1c40149a2acc5d876['h0073e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003a0] =  I38e438ab568822a1c40149a2acc5d876['h00740] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003a1] =  I38e438ab568822a1c40149a2acc5d876['h00742] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003a2] =  I38e438ab568822a1c40149a2acc5d876['h00744] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003a3] =  I38e438ab568822a1c40149a2acc5d876['h00746] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003a4] =  I38e438ab568822a1c40149a2acc5d876['h00748] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003a5] =  I38e438ab568822a1c40149a2acc5d876['h0074a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003a6] =  I38e438ab568822a1c40149a2acc5d876['h0074c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003a7] =  I38e438ab568822a1c40149a2acc5d876['h0074e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003a8] =  I38e438ab568822a1c40149a2acc5d876['h00750] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003a9] =  I38e438ab568822a1c40149a2acc5d876['h00752] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003aa] =  I38e438ab568822a1c40149a2acc5d876['h00754] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003ab] =  I38e438ab568822a1c40149a2acc5d876['h00756] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003ac] =  I38e438ab568822a1c40149a2acc5d876['h00758] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003ad] =  I38e438ab568822a1c40149a2acc5d876['h0075a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003ae] =  I38e438ab568822a1c40149a2acc5d876['h0075c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003af] =  I38e438ab568822a1c40149a2acc5d876['h0075e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003b0] =  I38e438ab568822a1c40149a2acc5d876['h00760] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003b1] =  I38e438ab568822a1c40149a2acc5d876['h00762] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003b2] =  I38e438ab568822a1c40149a2acc5d876['h00764] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003b3] =  I38e438ab568822a1c40149a2acc5d876['h00766] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003b4] =  I38e438ab568822a1c40149a2acc5d876['h00768] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003b5] =  I38e438ab568822a1c40149a2acc5d876['h0076a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003b6] =  I38e438ab568822a1c40149a2acc5d876['h0076c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003b7] =  I38e438ab568822a1c40149a2acc5d876['h0076e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003b8] =  I38e438ab568822a1c40149a2acc5d876['h00770] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003b9] =  I38e438ab568822a1c40149a2acc5d876['h00772] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003ba] =  I38e438ab568822a1c40149a2acc5d876['h00774] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003bb] =  I38e438ab568822a1c40149a2acc5d876['h00776] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003bc] =  I38e438ab568822a1c40149a2acc5d876['h00778] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003bd] =  I38e438ab568822a1c40149a2acc5d876['h0077a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003be] =  I38e438ab568822a1c40149a2acc5d876['h0077c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003bf] =  I38e438ab568822a1c40149a2acc5d876['h0077e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003c0] =  I38e438ab568822a1c40149a2acc5d876['h00780] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003c1] =  I38e438ab568822a1c40149a2acc5d876['h00782] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003c2] =  I38e438ab568822a1c40149a2acc5d876['h00784] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003c3] =  I38e438ab568822a1c40149a2acc5d876['h00786] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003c4] =  I38e438ab568822a1c40149a2acc5d876['h00788] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003c5] =  I38e438ab568822a1c40149a2acc5d876['h0078a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003c6] =  I38e438ab568822a1c40149a2acc5d876['h0078c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003c7] =  I38e438ab568822a1c40149a2acc5d876['h0078e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003c8] =  I38e438ab568822a1c40149a2acc5d876['h00790] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003c9] =  I38e438ab568822a1c40149a2acc5d876['h00792] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003ca] =  I38e438ab568822a1c40149a2acc5d876['h00794] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003cb] =  I38e438ab568822a1c40149a2acc5d876['h00796] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003cc] =  I38e438ab568822a1c40149a2acc5d876['h00798] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003cd] =  I38e438ab568822a1c40149a2acc5d876['h0079a] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003ce] =  I38e438ab568822a1c40149a2acc5d876['h0079c] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003cf] =  I38e438ab568822a1c40149a2acc5d876['h0079e] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003d0] =  I38e438ab568822a1c40149a2acc5d876['h007a0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003d1] =  I38e438ab568822a1c40149a2acc5d876['h007a2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003d2] =  I38e438ab568822a1c40149a2acc5d876['h007a4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003d3] =  I38e438ab568822a1c40149a2acc5d876['h007a6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003d4] =  I38e438ab568822a1c40149a2acc5d876['h007a8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003d5] =  I38e438ab568822a1c40149a2acc5d876['h007aa] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003d6] =  I38e438ab568822a1c40149a2acc5d876['h007ac] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003d7] =  I38e438ab568822a1c40149a2acc5d876['h007ae] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003d8] =  I38e438ab568822a1c40149a2acc5d876['h007b0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003d9] =  I38e438ab568822a1c40149a2acc5d876['h007b2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003da] =  I38e438ab568822a1c40149a2acc5d876['h007b4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003db] =  I38e438ab568822a1c40149a2acc5d876['h007b6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003dc] =  I38e438ab568822a1c40149a2acc5d876['h007b8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003dd] =  I38e438ab568822a1c40149a2acc5d876['h007ba] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003de] =  I38e438ab568822a1c40149a2acc5d876['h007bc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003df] =  I38e438ab568822a1c40149a2acc5d876['h007be] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003e0] =  I38e438ab568822a1c40149a2acc5d876['h007c0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003e1] =  I38e438ab568822a1c40149a2acc5d876['h007c2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003e2] =  I38e438ab568822a1c40149a2acc5d876['h007c4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003e3] =  I38e438ab568822a1c40149a2acc5d876['h007c6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003e4] =  I38e438ab568822a1c40149a2acc5d876['h007c8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003e5] =  I38e438ab568822a1c40149a2acc5d876['h007ca] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003e6] =  I38e438ab568822a1c40149a2acc5d876['h007cc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003e7] =  I38e438ab568822a1c40149a2acc5d876['h007ce] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003e8] =  I38e438ab568822a1c40149a2acc5d876['h007d0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003e9] =  I38e438ab568822a1c40149a2acc5d876['h007d2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003ea] =  I38e438ab568822a1c40149a2acc5d876['h007d4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003eb] =  I38e438ab568822a1c40149a2acc5d876['h007d6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003ec] =  I38e438ab568822a1c40149a2acc5d876['h007d8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003ed] =  I38e438ab568822a1c40149a2acc5d876['h007da] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003ee] =  I38e438ab568822a1c40149a2acc5d876['h007dc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003ef] =  I38e438ab568822a1c40149a2acc5d876['h007de] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003f0] =  I38e438ab568822a1c40149a2acc5d876['h007e0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003f1] =  I38e438ab568822a1c40149a2acc5d876['h007e2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003f2] =  I38e438ab568822a1c40149a2acc5d876['h007e4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003f3] =  I38e438ab568822a1c40149a2acc5d876['h007e6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003f4] =  I38e438ab568822a1c40149a2acc5d876['h007e8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003f5] =  I38e438ab568822a1c40149a2acc5d876['h007ea] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003f6] =  I38e438ab568822a1c40149a2acc5d876['h007ec] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003f7] =  I38e438ab568822a1c40149a2acc5d876['h007ee] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003f8] =  I38e438ab568822a1c40149a2acc5d876['h007f0] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003f9] =  I38e438ab568822a1c40149a2acc5d876['h007f2] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003fa] =  I38e438ab568822a1c40149a2acc5d876['h007f4] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003fb] =  I38e438ab568822a1c40149a2acc5d876['h007f6] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003fc] =  I38e438ab568822a1c40149a2acc5d876['h007f8] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003fd] =  I38e438ab568822a1c40149a2acc5d876['h007fa] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003fe] =  I38e438ab568822a1c40149a2acc5d876['h007fc] ;
//end
//always_comb begin // 
               I810764ca41a2b12d686e115c79b0578f['h003ff] =  I38e438ab568822a1c40149a2acc5d876['h007fe] ;
//end
