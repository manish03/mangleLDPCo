//`include "GF2_LDPC_flogtanh_0x0000c_assign_inc.sv"
//always_comb begin
              I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00000] = 
          (!flogtanh_sel['h0000c]) ? 
                       I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00000] : //%
                       I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00001] ;
//end
//always_comb begin
              I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00001] = 
          (!flogtanh_sel['h0000c]) ? 
                       I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00002] : //%
                       I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00003] ;
//end
//always_comb begin
              I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00002] = 
          (!flogtanh_sel['h0000c]) ? 
                       I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00004] : //%
                       I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00005] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00003] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00006] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00004] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00008] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00005] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0000a] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00006] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0000c] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00007] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0000e] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00008] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00010] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00009] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00012] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0000a] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00014] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0000b] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00016] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0000c] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00018] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0000d] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0001a] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0000e] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0001c] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0000f] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0001e] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00010] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00020] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00011] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00022] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00012] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00024] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00013] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00026] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00014] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00028] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00015] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0002a] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00016] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0002c] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00017] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0002e] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00018] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00030] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00019] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00032] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0001a] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00034] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0001b] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00036] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0001c] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00038] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0001d] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0003a] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0001e] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0003c] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0001f] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0003e] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00020] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00040] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00021] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00042] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00022] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00044] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00023] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00046] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00024] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00048] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00025] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0004a] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00026] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0004c] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00027] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0004e] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00028] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00050] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00029] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00052] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0002a] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00054] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0002b] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00056] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0002c] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00058] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0002d] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0005a] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0002e] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0005c] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0002f] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0005e] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00030] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00060] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00031] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00062] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00032] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00064] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00033] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00066] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00034] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00068] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00035] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0006a] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00036] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0006c] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00037] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0006e] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00038] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00070] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00039] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00072] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0003a] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00074] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0003b] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00076] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0003c] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00078] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0003d] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0007a] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0003e] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0007c] ;
//end
//always_comb begin // 
               I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0003f] =  I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0007e] ;
//end
