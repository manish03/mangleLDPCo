 reg  ['h1ff:0] [$clog2('h7000+1)-1:0] I986ccea2f9226242e2772b9c3af42d87 ;
