reg [fgallag_WDTH -1:0] Ic95a3f9bce1f573855ca615170882870, I999768f7a0479b93e065e98bb8d71bb7;
reg [fgallag_WDTH -1:0] I7b13a2539c028f1b1704554ec14280f5, I6668f7bb8dc077f0ff1cac6d088185c3;
reg [fgallag_WDTH -1:0] I9b426da62c1159dd95754d51e3d8b4e8, I99ce11aaea6da1dfb5d0567597b95ef4;
reg [fgallag_WDTH -1:0] I77a77a7a6a437c395358b6f0beafd9f2, I75b52e5dd015a0e0cfc2f7d453857ccd;
reg [fgallag_WDTH -1:0] I1efd99d9686a0c7e1187d852a3572023, If01ebfc5e8f0038e0fd309e8b69f89e4;
reg [fgallag_WDTH -1:0] Ia0c03de62b7bfb76e6fea17bd0e8d003, Id265f18fa76b685483b0694a5bb7ed43;
reg Ic5f8ad0b8b66b30eaaee70ac52ea6465 ;
always @(posedge clk or negedge rstn)
if (!rstn) begin
 I999768f7a0479b93e065e98bb8d71bb7 <= 'h0;
 I6668f7bb8dc077f0ff1cac6d088185c3 <= 'h0;
 I99ce11aaea6da1dfb5d0567597b95ef4 <= 'h0;
 I75b52e5dd015a0e0cfc2f7d453857ccd <= 'h0;
 If01ebfc5e8f0038e0fd309e8b69f89e4 <= 'h0;
 Id265f18fa76b685483b0694a5bb7ed43 <= 'h0;
 Ic5f8ad0b8b66b30eaaee70ac52ea6465 <= 'h0;
end
else
begin
 I999768f7a0479b93e065e98bb8d71bb7 <=  Ic95a3f9bce1f573855ca615170882870;
 I6668f7bb8dc077f0ff1cac6d088185c3 <=  I7b13a2539c028f1b1704554ec14280f5;
 I99ce11aaea6da1dfb5d0567597b95ef4 <=  I9b426da62c1159dd95754d51e3d8b4e8;
 I75b52e5dd015a0e0cfc2f7d453857ccd <=  I77a77a7a6a437c395358b6f0beafd9f2;
 If01ebfc5e8f0038e0fd309e8b69f89e4 <=  I1efd99d9686a0c7e1187d852a3572023;
 Id265f18fa76b685483b0694a5bb7ed43 <=  Ia0c03de62b7bfb76e6fea17bd0e8d003;
 Ic5f8ad0b8b66b30eaaee70ac52ea6465 <=  If677b4bb108ef735b4ad076cbbfd3094;
end
