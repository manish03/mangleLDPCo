 reg  ['hfff:0] [$clog2('h7000+1)-1:0] Ic8a4ab93493bd6cdd4939054e46d2247 ;
