//`include "GF2_LDPC_flogtanh_0x0000b_assign_inc.sv"
//always_comb begin
              I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00000] = 
          (!flogtanh_sel['h0000b]) ? 
                       I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00000] : //%
                       I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00001] ;
//end
//always_comb begin
              I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00001] = 
          (!flogtanh_sel['h0000b]) ? 
                       I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00002] : //%
                       I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00003] ;
//end
//always_comb begin
              I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00002] = 
          (!flogtanh_sel['h0000b]) ? 
                       I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00004] : //%
                       I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00005] ;
//end
//always_comb begin
              I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00003] = 
          (!flogtanh_sel['h0000b]) ? 
                       I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00006] : //%
                       I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00007] ;
//end
//always_comb begin
              I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00004] = 
          (!flogtanh_sel['h0000b]) ? 
                       I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00008] : //%
                       I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00009] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00005] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0000a] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00006] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0000c] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00007] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0000e] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00008] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00010] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00009] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00012] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0000a] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00014] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0000b] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00016] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0000c] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00018] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0000d] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0001a] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0000e] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0001c] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0000f] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0001e] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00010] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00020] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00011] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00022] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00012] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00024] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00013] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00026] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00014] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00028] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00015] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0002a] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00016] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0002c] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00017] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0002e] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00018] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00030] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00019] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00032] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0001a] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00034] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0001b] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00036] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0001c] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00038] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0001d] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0003a] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0001e] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0003c] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0001f] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0003e] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00020] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00040] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00021] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00042] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00022] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00044] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00023] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00046] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00024] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00048] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00025] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0004a] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00026] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0004c] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00027] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0004e] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00028] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00050] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00029] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00052] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0002a] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00054] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0002b] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00056] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0002c] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00058] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0002d] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0005a] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0002e] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0005c] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0002f] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0005e] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00030] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00060] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00031] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00062] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00032] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00064] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00033] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00066] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00034] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00068] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00035] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0006a] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00036] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0006c] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00037] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0006e] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00038] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00070] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00039] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00072] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0003a] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00074] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0003b] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00076] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0003c] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00078] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0003d] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0007a] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0003e] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0007c] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0003f] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0007e] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00040] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00080] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00041] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00082] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00042] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00084] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00043] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00086] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00044] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00088] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00045] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0008a] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00046] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0008c] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00047] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0008e] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00048] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00090] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00049] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00092] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0004a] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00094] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0004b] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00096] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0004c] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00098] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0004d] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0009a] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0004e] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0009c] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0004f] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0009e] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00050] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000a0] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00051] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000a2] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00052] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000a4] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00053] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000a6] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00054] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000a8] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00055] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000aa] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00056] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000ac] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00057] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000ae] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00058] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000b0] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00059] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000b2] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0005a] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000b4] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0005b] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000b6] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0005c] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000b8] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0005d] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000ba] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0005e] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000bc] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0005f] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000be] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00060] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000c0] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00061] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000c2] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00062] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000c4] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00063] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000c6] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00064] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000c8] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00065] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000ca] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00066] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000cc] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00067] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000ce] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00068] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000d0] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00069] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000d2] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0006a] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000d4] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0006b] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000d6] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0006c] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000d8] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0006d] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000da] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0006e] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000dc] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0006f] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000de] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00070] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000e0] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00071] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000e2] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00072] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000e4] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00073] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000e6] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00074] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000e8] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00075] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000ea] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00076] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000ec] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00077] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000ee] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00078] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000f0] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h00079] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000f2] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0007a] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000f4] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0007b] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000f6] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0007c] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000f8] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0007d] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000fa] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0007e] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000fc] ;
//end
//always_comb begin // 
               I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211['h0007f] =  I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000fe] ;
//end
