 reg  ['h1fff:0] [$clog2('h7000+1)-1:0] I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2 ;
