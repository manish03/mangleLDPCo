 reg  ['h3f:0] [$clog2('h7000+1)-1:0] Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6 ;
