reg [flogtanh_WDTH -1:0] Ib2aa0dad949a7608d49dfdec8811fead, I12635a66e3fe4dd930e858a0a7580cea;
reg [flogtanh_WDTH -1:0] Ia6b922271dbe47dd60eb4d0492fd5739, I71130fa5b933e0e26dbab66f37fb8925;
reg [flogtanh_WDTH -1:0] Idf881bd96e29e48e7efacbb467ff7c5c, I9371a6ffdba2a5bd6c4ac3fb38010117;
reg [flogtanh_WDTH -1:0] I20717481aece4914e0f7222ae35d1456, I4001f1ca6d56d63aca19160a999b23de;
reg [flogtanh_WDTH -1:0] Ifcfb5c6c620ff437f7830d0c6d939e62, Icf4458bcd36b49edb3c99d94980b2fcf;
reg [flogtanh_WDTH -1:0] I286aa151ea1dba5e7e6c4639e80b8cf2, Ia336a15ef64f48975747202ff0586f96;
reg [flogtanh_WDTH -1:0] Ia14165ce5e9de831dcd289ac0495e42e, I0ab4d4499b838b988c31c5d2162b0aa2;
reg [flogtanh_WDTH -1:0] Iad283604bd9143b0729e1d7d1f49dfbb, I8cc0695ebf79a9943050729478d73c9c;
reg [flogtanh_WDTH -1:0] If14b995d06822c80d9d714d4bbbcda58, I1207b10797bccdad5ee7e32abbfc9531;
reg [flogtanh_WDTH -1:0] Iece268d0f9e7bdda5bcf50208cf24762, Ie37f7a4132d9db8e6589e4818da8f71e;
reg [flogtanh_WDTH -1:0] I087bd6d6037f7ee9e82663387ac0f820, Ief67dacff61c30f4f07a8b9426499320;
reg [flogtanh_WDTH -1:0] I0c2fb3d39b747d63854302c08ec8b1c2, I64c9510573d0b631cd08f41a30b4bf94;
reg [flogtanh_WDTH -1:0] Id3d9536b013c4766333f6d23066ead54, I496d08bbbe57943dde0a060794dd44f2;
reg [flogtanh_WDTH -1:0] Ibc1ee835e7e2d5432583440c90304c56, I6ea770088be3718bb9cbbf4015d7a698;
reg [flogtanh_WDTH -1:0] I594ca16757d13f9bd17dae2114615a80, I96e8e53f5e2fe546281cb33632075218;
reg [flogtanh_WDTH -1:0] Id7f43a01fda8433c8b72871f35ef7bdc, Iad67f635fc879ccccb83e4e8090e851f;
reg [flogtanh_WDTH -1:0] Id850fafd66d7cd6901821100a3290a23, Ic4eeb8715a3ab8d9da059d43c2f73e31;
reg [flogtanh_WDTH -1:0] I9a0a13f48f3e52b33be36fe03a9f2da3, I06d19f878da9b67396ff63c2b0ac8a1e;
reg [flogtanh_WDTH -1:0] I77ad3e9b4bafb0b2a4e86f453c9c59a0, Ied5797945822a58d6850b3d5472b6657;
reg [flogtanh_WDTH -1:0] Ic3b0467ebe638a2bd44437784b22329e, I79706d7caf960d3eee136724e1474c14;
reg [flogtanh_WDTH -1:0] Id57e199202dd2b2fd585b7cbde5f2ad3, Ic43fc3a05372e660dd974dd41d61966d;
reg [flogtanh_WDTH -1:0] I03ea04be646c4834304d4f82d3171243, Id05004336c93a8f315406a56d1ea9401;
reg [flogtanh_WDTH -1:0] I8ac44624c0749e8e870c9dde42ffb8dd, I4257f21c0512ab632f6d8e3e49b6bc86;
reg [flogtanh_WDTH -1:0] I7852770263dd0c5503c75135d38058c4, I38e64d8c0bfe85f483b46ad9d510bbf1;
reg [flogtanh_WDTH -1:0] Icf8a31b29e9f8918802c3bf5baa48fa5, If9f0572284b7c7b6fe299fb8f45c57d5;
reg [flogtanh_WDTH -1:0] I94a9a947dc58e38c7c3e13bf1bab6f51, I248384903432b0ea141bdb0ba98bd3a3;
reg [flogtanh_WDTH -1:0] Ic92921fa31c014ee1c49384973b33176, I81f42775b2a3e4badcc3910838808691;
reg [flogtanh_WDTH -1:0] Iabedd360b191a5862ad534eea51ab52e, Iec5241a1c42d080412dff5e9494851e9;
reg [flogtanh_WDTH -1:0] I4659f7245c85f3db58d6be3f97cb3cf0, I1f10ad5fe2f55ebdb372cc672d8dd978;
reg [flogtanh_WDTH -1:0] I164cbb304f4db6a716bd788036086266, I1ca0505131c6887eaf1e7e80473e3add;
reg [flogtanh_WDTH -1:0] I8775c4f7dd528188506d94cc13862f93, Ib49ad95d66dc9b1f5b9b225aa8124010;
reg [flogtanh_WDTH -1:0] Ibb600c26f9f0972df669d2d04a96c7f6, I1d942dd2be55359b99052dc72e795590;
reg [flogtanh_WDTH -1:0] Ied0b82caf207f1992f7ec334a9fb423c, Id414b502a923f77f986b3c2f223798c4;
reg [flogtanh_WDTH -1:0] I235cbb8f044d1ac3bf4f53c932b5a34b, I0b6ec8b66cdd200b2eb618e53a9a3bc1;
reg [flogtanh_WDTH -1:0] I1d25723c499c68dea49c4d762d80bcc3, I1178b66ba1832d0acdf2683631bcebcc;
reg [flogtanh_WDTH -1:0] I6309f136f930378ab3b8cf5a29cfafdf, I361d0be38e55d517342ea4b081c0fc23;
reg [flogtanh_WDTH -1:0] I4d5d1e9c151f5e4e18596916c57b891d, I11ea42222da256fa229e3f7f74a29fd1;
reg [flogtanh_WDTH -1:0] I134c07a35862ad54f8852c17a8bab5de, I2ac252803e9dee4dde03c09629f6a8dc;
reg [flogtanh_WDTH -1:0] I5b663cc1d7cc3069f33b63799aa34796, I7714bd5031cea3a279cf989b22b30579;
reg [flogtanh_WDTH -1:0] Ia2ed52a8130a197b3a198aa454d980b0, Ifed18851e47a0fe3da23dee1e77aa07b;
reg [flogtanh_WDTH -1:0] I13acb2c915e11641c53157310e44892b, Ic1ffa3d6c9037998cdf86b17c269216b;
reg [flogtanh_WDTH -1:0] I6a5212af01917f8e71e3e83bd9e8caf2, Ieceeefbdcb9554432f7568493e4b532f;
reg [flogtanh_WDTH -1:0] I3fe2af1aa64d019af984fa86c1292ad9, I7780a0f25847a4e699619e564751c9a2;
reg [flogtanh_WDTH -1:0] Ic09f027112d6b05b07873fda8e85bea2, I8a966b7a6353ba171cc98fb541e80623;
reg [flogtanh_WDTH -1:0] If35467fdae216528f1dd248b2c19feba, I64e434f7354d5b36a40f23792bed6616;
reg [flogtanh_WDTH -1:0] I6681491d836b3bf63f771b708625f7b6, Iae66d17c285d26bc13a560a3c46768ca;
reg Id11ca9ab1b4b30c21f7314a04c9c7fae ;
always @(posedge clk or negedge rstn)
if (!rstn) begin
 I12635a66e3fe4dd930e858a0a7580cea <= 'h0;
 I71130fa5b933e0e26dbab66f37fb8925 <= 'h0;
 I9371a6ffdba2a5bd6c4ac3fb38010117 <= 'h0;
 I4001f1ca6d56d63aca19160a999b23de <= 'h0;
 Icf4458bcd36b49edb3c99d94980b2fcf <= 'h0;
 Ia336a15ef64f48975747202ff0586f96 <= 'h0;
 I0ab4d4499b838b988c31c5d2162b0aa2 <= 'h0;
 I8cc0695ebf79a9943050729478d73c9c <= 'h0;
 I1207b10797bccdad5ee7e32abbfc9531 <= 'h0;
 Ie37f7a4132d9db8e6589e4818da8f71e <= 'h0;
 Ief67dacff61c30f4f07a8b9426499320 <= 'h0;
 I64c9510573d0b631cd08f41a30b4bf94 <= 'h0;
 I496d08bbbe57943dde0a060794dd44f2 <= 'h0;
 I6ea770088be3718bb9cbbf4015d7a698 <= 'h0;
 I96e8e53f5e2fe546281cb33632075218 <= 'h0;
 Iad67f635fc879ccccb83e4e8090e851f <= 'h0;
 Ic4eeb8715a3ab8d9da059d43c2f73e31 <= 'h0;
 I06d19f878da9b67396ff63c2b0ac8a1e <= 'h0;
 Ied5797945822a58d6850b3d5472b6657 <= 'h0;
 I79706d7caf960d3eee136724e1474c14 <= 'h0;
 Ic43fc3a05372e660dd974dd41d61966d <= 'h0;
 Id05004336c93a8f315406a56d1ea9401 <= 'h0;
 I4257f21c0512ab632f6d8e3e49b6bc86 <= 'h0;
 I38e64d8c0bfe85f483b46ad9d510bbf1 <= 'h0;
 If9f0572284b7c7b6fe299fb8f45c57d5 <= 'h0;
 I248384903432b0ea141bdb0ba98bd3a3 <= 'h0;
 I81f42775b2a3e4badcc3910838808691 <= 'h0;
 Iec5241a1c42d080412dff5e9494851e9 <= 'h0;
 I1f10ad5fe2f55ebdb372cc672d8dd978 <= 'h0;
 I1ca0505131c6887eaf1e7e80473e3add <= 'h0;
 Ib49ad95d66dc9b1f5b9b225aa8124010 <= 'h0;
 I1d942dd2be55359b99052dc72e795590 <= 'h0;
 Id414b502a923f77f986b3c2f223798c4 <= 'h0;
 I0b6ec8b66cdd200b2eb618e53a9a3bc1 <= 'h0;
 I1178b66ba1832d0acdf2683631bcebcc <= 'h0;
 I361d0be38e55d517342ea4b081c0fc23 <= 'h0;
 I11ea42222da256fa229e3f7f74a29fd1 <= 'h0;
 I2ac252803e9dee4dde03c09629f6a8dc <= 'h0;
 I7714bd5031cea3a279cf989b22b30579 <= 'h0;
 Ifed18851e47a0fe3da23dee1e77aa07b <= 'h0;
 Ic1ffa3d6c9037998cdf86b17c269216b <= 'h0;
 Ieceeefbdcb9554432f7568493e4b532f <= 'h0;
 I7780a0f25847a4e699619e564751c9a2 <= 'h0;
 I8a966b7a6353ba171cc98fb541e80623 <= 'h0;
 I64e434f7354d5b36a40f23792bed6616 <= 'h0;
 Iae66d17c285d26bc13a560a3c46768ca <= 'h0;
 Id11ca9ab1b4b30c21f7314a04c9c7fae <= 'h0;
end
else
begin
 I12635a66e3fe4dd930e858a0a7580cea <=  Ib2aa0dad949a7608d49dfdec8811fead;
 I71130fa5b933e0e26dbab66f37fb8925 <=  Ia6b922271dbe47dd60eb4d0492fd5739;
 I9371a6ffdba2a5bd6c4ac3fb38010117 <=  Idf881bd96e29e48e7efacbb467ff7c5c;
 I4001f1ca6d56d63aca19160a999b23de <=  I20717481aece4914e0f7222ae35d1456;
 Icf4458bcd36b49edb3c99d94980b2fcf <=  Ifcfb5c6c620ff437f7830d0c6d939e62;
 Ia336a15ef64f48975747202ff0586f96 <=  I286aa151ea1dba5e7e6c4639e80b8cf2;
 I0ab4d4499b838b988c31c5d2162b0aa2 <=  Ia14165ce5e9de831dcd289ac0495e42e;
 I8cc0695ebf79a9943050729478d73c9c <=  Iad283604bd9143b0729e1d7d1f49dfbb;
 I1207b10797bccdad5ee7e32abbfc9531 <=  If14b995d06822c80d9d714d4bbbcda58;
 Ie37f7a4132d9db8e6589e4818da8f71e <=  Iece268d0f9e7bdda5bcf50208cf24762;
 Ief67dacff61c30f4f07a8b9426499320 <=  I087bd6d6037f7ee9e82663387ac0f820;
 I64c9510573d0b631cd08f41a30b4bf94 <=  I0c2fb3d39b747d63854302c08ec8b1c2;
 I496d08bbbe57943dde0a060794dd44f2 <=  Id3d9536b013c4766333f6d23066ead54;
 I6ea770088be3718bb9cbbf4015d7a698 <=  Ibc1ee835e7e2d5432583440c90304c56;
 I96e8e53f5e2fe546281cb33632075218 <=  I594ca16757d13f9bd17dae2114615a80;
 Iad67f635fc879ccccb83e4e8090e851f <=  Id7f43a01fda8433c8b72871f35ef7bdc;
 Ic4eeb8715a3ab8d9da059d43c2f73e31 <=  Id850fafd66d7cd6901821100a3290a23;
 I06d19f878da9b67396ff63c2b0ac8a1e <=  I9a0a13f48f3e52b33be36fe03a9f2da3;
 Ied5797945822a58d6850b3d5472b6657 <=  I77ad3e9b4bafb0b2a4e86f453c9c59a0;
 I79706d7caf960d3eee136724e1474c14 <=  Ic3b0467ebe638a2bd44437784b22329e;
 Ic43fc3a05372e660dd974dd41d61966d <=  Id57e199202dd2b2fd585b7cbde5f2ad3;
 Id05004336c93a8f315406a56d1ea9401 <=  I03ea04be646c4834304d4f82d3171243;
 I4257f21c0512ab632f6d8e3e49b6bc86 <=  I8ac44624c0749e8e870c9dde42ffb8dd;
 I38e64d8c0bfe85f483b46ad9d510bbf1 <=  I7852770263dd0c5503c75135d38058c4;
 If9f0572284b7c7b6fe299fb8f45c57d5 <=  Icf8a31b29e9f8918802c3bf5baa48fa5;
 I248384903432b0ea141bdb0ba98bd3a3 <=  I94a9a947dc58e38c7c3e13bf1bab6f51;
 I81f42775b2a3e4badcc3910838808691 <=  Ic92921fa31c014ee1c49384973b33176;
 Iec5241a1c42d080412dff5e9494851e9 <=  Iabedd360b191a5862ad534eea51ab52e;
 I1f10ad5fe2f55ebdb372cc672d8dd978 <=  I4659f7245c85f3db58d6be3f97cb3cf0;
 I1ca0505131c6887eaf1e7e80473e3add <=  I164cbb304f4db6a716bd788036086266;
 Ib49ad95d66dc9b1f5b9b225aa8124010 <=  I8775c4f7dd528188506d94cc13862f93;
 I1d942dd2be55359b99052dc72e795590 <=  Ibb600c26f9f0972df669d2d04a96c7f6;
 Id414b502a923f77f986b3c2f223798c4 <=  Ied0b82caf207f1992f7ec334a9fb423c;
 I0b6ec8b66cdd200b2eb618e53a9a3bc1 <=  I235cbb8f044d1ac3bf4f53c932b5a34b;
 I1178b66ba1832d0acdf2683631bcebcc <=  I1d25723c499c68dea49c4d762d80bcc3;
 I361d0be38e55d517342ea4b081c0fc23 <=  I6309f136f930378ab3b8cf5a29cfafdf;
 I11ea42222da256fa229e3f7f74a29fd1 <=  I4d5d1e9c151f5e4e18596916c57b891d;
 I2ac252803e9dee4dde03c09629f6a8dc <=  I134c07a35862ad54f8852c17a8bab5de;
 I7714bd5031cea3a279cf989b22b30579 <=  I5b663cc1d7cc3069f33b63799aa34796;
 Ifed18851e47a0fe3da23dee1e77aa07b <=  Ia2ed52a8130a197b3a198aa454d980b0;
 Ic1ffa3d6c9037998cdf86b17c269216b <=  I13acb2c915e11641c53157310e44892b;
 Ieceeefbdcb9554432f7568493e4b532f <=  I6a5212af01917f8e71e3e83bd9e8caf2;
 I7780a0f25847a4e699619e564751c9a2 <=  I3fe2af1aa64d019af984fa86c1292ad9;
 I8a966b7a6353ba171cc98fb541e80623 <=  Ic09f027112d6b05b07873fda8e85bea2;
 I64e434f7354d5b36a40f23792bed6616 <=  If35467fdae216528f1dd248b2c19feba;
 Iae66d17c285d26bc13a560a3c46768ca <=  I6681491d836b3bf63f771b708625f7b6;
 Id11ca9ab1b4b30c21f7314a04c9c7fae <=  If6d744ed5db03bac562b8bea5fd72479;
end
