 reg  ['h3f:0] [$clog2('h7000+1)-1:0] Ie4acdb20b1de9050267f708a13a337e0 ;
