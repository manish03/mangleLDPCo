 reg  ['h7ff:0] [$clog2('h7000+1)-1:0] I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed ;
