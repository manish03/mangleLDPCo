//`include "GF2_LDPC_fgallag_0x0000a_assign_inc.sv"
//always_comb begin
              Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00000] = 
          (!fgallag_sel['h0000a]) ? 
                       Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00000] : //%
                       Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00001] ;
//end
//always_comb begin
              Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00001] = 
          (!fgallag_sel['h0000a]) ? 
                       Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00002] : //%
                       Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00003] ;
//end
//always_comb begin
              Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00002] = 
          (!fgallag_sel['h0000a]) ? 
                       Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00004] : //%
                       Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00005] ;
//end
//always_comb begin
              Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00003] = 
          (!fgallag_sel['h0000a]) ? 
                       Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00006] : //%
                       Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00007] ;
//end
//always_comb begin
              Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00004] = 
          (!fgallag_sel['h0000a]) ? 
                       Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00008] : //%
                       Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00009] ;
//end
//always_comb begin
              Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00005] = 
          (!fgallag_sel['h0000a]) ? 
                       Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0000a] : //%
                       Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0000b] ;
//end
//always_comb begin
              Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00006] = 
          (!fgallag_sel['h0000a]) ? 
                       Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0000c] : //%
                       Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0000d] ;
//end
//always_comb begin
              Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00007] = 
          (!fgallag_sel['h0000a]) ? 
                       Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0000e] : //%
                       Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0000f] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00008] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00010] ;
//end
//always_comb begin
              Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00009] = 
          (!fgallag_sel['h0000a]) ? 
                       Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00012] : //%
                       Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00013] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0000a] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00014] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0000b] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00016] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0000c] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00018] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0000d] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0001a] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0000e] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0001c] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0000f] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0001e] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00010] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00020] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00011] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00022] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00012] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00024] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00013] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00026] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00014] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00028] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00015] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0002a] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00016] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0002c] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00017] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0002e] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00018] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00030] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00019] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00032] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0001a] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00034] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0001b] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00036] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0001c] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00038] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0001d] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0003a] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0001e] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0003c] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0001f] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0003e] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00020] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00040] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00021] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00042] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00022] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00044] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00023] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00046] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00024] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00048] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00025] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0004a] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00026] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0004c] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00027] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0004e] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00028] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00050] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00029] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00052] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0002a] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00054] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0002b] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00056] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0002c] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00058] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0002d] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0005a] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0002e] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0005c] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0002f] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0005e] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00030] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00060] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00031] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00062] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00032] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00064] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00033] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00066] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00034] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00068] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00035] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0006a] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00036] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0006c] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00037] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0006e] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00038] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00070] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00039] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00072] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0003a] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00074] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0003b] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00076] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0003c] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00078] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0003d] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0007a] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0003e] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0007c] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0003f] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0007e] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00040] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00080] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00041] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00082] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00042] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00084] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00043] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00086] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00044] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00088] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00045] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0008a] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00046] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0008c] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00047] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0008e] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00048] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00090] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00049] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00092] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0004a] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00094] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0004b] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00096] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0004c] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00098] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0004d] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0009a] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0004e] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0009c] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0004f] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0009e] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00050] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000a0] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00051] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000a2] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00052] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000a4] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00053] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000a6] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00054] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000a8] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00055] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000aa] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00056] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000ac] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00057] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000ae] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00058] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000b0] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00059] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000b2] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0005a] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000b4] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0005b] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000b6] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0005c] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000b8] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0005d] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000ba] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0005e] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000bc] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0005f] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000be] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00060] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000c0] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00061] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000c2] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00062] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000c4] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00063] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000c6] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00064] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000c8] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00065] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000ca] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00066] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000cc] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00067] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000ce] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00068] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000d0] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00069] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000d2] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0006a] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000d4] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0006b] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000d6] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0006c] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000d8] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0006d] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000da] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0006e] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000dc] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0006f] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000de] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00070] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000e0] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00071] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000e2] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00072] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000e4] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00073] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000e6] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00074] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000e8] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00075] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000ea] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00076] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000ec] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00077] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000ee] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00078] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000f0] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00079] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000f2] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0007a] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000f4] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0007b] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000f6] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0007c] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000f8] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0007d] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000fa] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0007e] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000fc] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0007f] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000fe] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00080] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00100] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00081] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00102] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00082] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00104] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00083] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00106] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00084] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00108] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00085] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0010a] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00086] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0010c] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00087] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0010e] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00088] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00110] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00089] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00112] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0008a] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00114] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0008b] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00116] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0008c] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00118] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0008d] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0011a] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0008e] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0011c] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0008f] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0011e] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00090] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00120] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00091] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00122] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00092] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00124] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00093] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00126] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00094] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00128] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00095] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0012a] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00096] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0012c] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00097] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0012e] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00098] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00130] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00099] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00132] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0009a] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00134] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0009b] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00136] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0009c] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00138] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0009d] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0013a] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0009e] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0013c] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0009f] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0013e] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000a0] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00140] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000a1] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00142] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000a2] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00144] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000a3] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00146] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000a4] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00148] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000a5] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0014a] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000a6] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0014c] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000a7] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0014e] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000a8] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00150] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000a9] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00152] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000aa] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00154] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000ab] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00156] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000ac] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00158] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000ad] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0015a] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000ae] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0015c] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000af] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0015e] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000b0] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00160] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000b1] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00162] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000b2] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00164] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000b3] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00166] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000b4] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00168] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000b5] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0016a] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000b6] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0016c] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000b7] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0016e] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000b8] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00170] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000b9] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00172] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000ba] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00174] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000bb] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00176] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000bc] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00178] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000bd] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0017a] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000be] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0017c] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000bf] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0017e] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000c0] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00180] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000c1] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00182] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000c2] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00184] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000c3] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00186] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000c4] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00188] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000c5] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0018a] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000c6] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0018c] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000c7] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0018e] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000c8] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00190] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000c9] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00192] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000ca] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00194] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000cb] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00196] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000cc] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00198] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000cd] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0019a] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000ce] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0019c] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000cf] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0019e] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000d0] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001a0] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000d1] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001a2] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000d2] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001a4] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000d3] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001a6] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000d4] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001a8] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000d5] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001aa] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000d6] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001ac] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000d7] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001ae] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000d8] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001b0] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000d9] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001b2] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000da] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001b4] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000db] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001b6] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000dc] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001b8] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000dd] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001ba] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000de] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001bc] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000df] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001be] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000e0] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001c0] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000e1] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001c2] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000e2] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001c4] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000e3] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001c6] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000e4] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001c8] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000e5] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001ca] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000e6] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001cc] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000e7] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001ce] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000e8] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001d0] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000e9] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001d2] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000ea] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001d4] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000eb] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001d6] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000ec] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001d8] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000ed] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001da] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000ee] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001dc] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000ef] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001de] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000f0] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001e0] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000f1] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001e2] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000f2] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001e4] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000f3] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001e6] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000f4] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001e8] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000f5] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001ea] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000f6] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001ec] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000f7] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001ee] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000f8] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001f0] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000f9] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001f2] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000fa] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001f4] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000fb] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001f6] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000fc] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001f8] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000fd] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001fa] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000fe] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001fc] ;
//end
//always_comb begin // 
               Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000ff] =  Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001fe] ;
//end
