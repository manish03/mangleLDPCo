 reg  ['hf:0] [$clog2('h7000+1)-1:0] I333510d8572134ddfb62c52fc8869a236241ec893f038dd668e3222609245de0 ;
