//`include "GF2_LDPC_fgallag_0x00009_assign_inc.sv"
//always_comb begin
              Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00000] = 
          (!fgallag_sel['h00009]) ? 
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00000] : //%
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00001] ;
//end
//always_comb begin
              Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00001] = 
          (!fgallag_sel['h00009]) ? 
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00002] : //%
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00003] ;
//end
//always_comb begin
              Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00002] = 
          (!fgallag_sel['h00009]) ? 
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00004] : //%
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00005] ;
//end
//always_comb begin
              Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00003] = 
          (!fgallag_sel['h00009]) ? 
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00006] : //%
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00007] ;
//end
//always_comb begin
              Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00004] = 
          (!fgallag_sel['h00009]) ? 
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00008] : //%
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00009] ;
//end
//always_comb begin
              Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00005] = 
          (!fgallag_sel['h00009]) ? 
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0000a] : //%
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0000b] ;
//end
//always_comb begin
              Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00006] = 
          (!fgallag_sel['h00009]) ? 
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0000c] : //%
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0000d] ;
//end
//always_comb begin
              Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00007] = 
          (!fgallag_sel['h00009]) ? 
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0000e] : //%
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0000f] ;
//end
//always_comb begin
              Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00008] = 
          (!fgallag_sel['h00009]) ? 
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00010] : //%
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00011] ;
//end
//always_comb begin
              Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00009] = 
          (!fgallag_sel['h00009]) ? 
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00012] : //%
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00013] ;
//end
//always_comb begin
              Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0000a] = 
          (!fgallag_sel['h00009]) ? 
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00014] : //%
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00015] ;
//end
//always_comb begin
              Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0000b] = 
          (!fgallag_sel['h00009]) ? 
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00016] : //%
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00017] ;
//end
//always_comb begin
              Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0000c] = 
          (!fgallag_sel['h00009]) ? 
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00018] : //%
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00019] ;
//end
//always_comb begin
              Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0000d] = 
          (!fgallag_sel['h00009]) ? 
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0001a] : //%
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0001b] ;
//end
//always_comb begin
              Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0000e] = 
          (!fgallag_sel['h00009]) ? 
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0001c] : //%
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0001d] ;
//end
//always_comb begin
              Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0000f] = 
          (!fgallag_sel['h00009]) ? 
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0001e] : //%
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0001f] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00010] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00020] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00011] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00022] ;
//end
//always_comb begin
              Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00012] = 
          (!fgallag_sel['h00009]) ? 
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00024] : //%
                       I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00025] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00013] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00026] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00014] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00028] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00015] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0002a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00016] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0002c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00017] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0002e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00018] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00030] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00019] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00032] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0001a] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00034] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0001b] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00036] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0001c] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00038] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0001d] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0003a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0001e] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0003c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0001f] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0003e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00020] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00040] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00021] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00042] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00022] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00044] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00023] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00046] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00024] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00048] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00025] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0004a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00026] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0004c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00027] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0004e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00028] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00050] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00029] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00052] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0002a] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00054] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0002b] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00056] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0002c] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00058] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0002d] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0005a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0002e] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0005c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0002f] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0005e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00030] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00060] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00031] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00062] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00032] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00064] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00033] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00066] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00034] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00068] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00035] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0006a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00036] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0006c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00037] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0006e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00038] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00070] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00039] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00072] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0003a] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00074] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0003b] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00076] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0003c] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00078] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0003d] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0007a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0003e] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0007c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0003f] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0007e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00040] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00080] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00041] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00082] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00042] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00084] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00043] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00086] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00044] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00088] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00045] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0008a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00046] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0008c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00047] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0008e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00048] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00090] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00049] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00092] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0004a] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00094] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0004b] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00096] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0004c] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00098] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0004d] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0009a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0004e] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0009c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0004f] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0009e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00050] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000a0] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00051] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000a2] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00052] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000a4] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00053] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000a6] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00054] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000a8] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00055] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000aa] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00056] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000ac] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00057] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000ae] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00058] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000b0] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00059] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000b2] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0005a] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000b4] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0005b] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000b6] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0005c] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000b8] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0005d] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000ba] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0005e] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000bc] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0005f] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000be] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00060] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000c0] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00061] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000c2] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00062] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000c4] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00063] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000c6] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00064] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000c8] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00065] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000ca] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00066] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000cc] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00067] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000ce] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00068] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000d0] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00069] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000d2] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0006a] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000d4] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0006b] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000d6] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0006c] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000d8] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0006d] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000da] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0006e] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000dc] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0006f] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000de] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00070] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000e0] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00071] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000e2] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00072] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000e4] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00073] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000e6] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00074] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000e8] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00075] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000ea] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00076] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000ec] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00077] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000ee] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00078] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000f0] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00079] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000f2] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0007a] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000f4] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0007b] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000f6] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0007c] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000f8] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0007d] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000fa] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0007e] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000fc] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0007f] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000fe] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00080] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00100] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00081] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00102] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00082] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00104] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00083] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00106] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00084] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00108] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00085] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0010a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00086] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0010c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00087] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0010e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00088] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00110] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00089] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00112] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0008a] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00114] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0008b] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00116] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0008c] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00118] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0008d] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0011a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0008e] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0011c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0008f] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0011e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00090] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00120] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00091] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00122] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00092] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00124] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00093] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00126] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00094] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00128] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00095] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0012a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00096] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0012c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00097] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0012e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00098] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00130] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00099] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00132] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0009a] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00134] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0009b] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00136] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0009c] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00138] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0009d] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0013a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0009e] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0013c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0009f] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0013e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000a0] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00140] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000a1] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00142] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000a2] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00144] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000a3] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00146] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000a4] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00148] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000a5] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0014a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000a6] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0014c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000a7] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0014e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000a8] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00150] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000a9] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00152] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000aa] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00154] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000ab] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00156] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000ac] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00158] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000ad] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0015a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000ae] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0015c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000af] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0015e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000b0] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00160] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000b1] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00162] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000b2] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00164] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000b3] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00166] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000b4] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00168] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000b5] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0016a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000b6] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0016c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000b7] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0016e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000b8] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00170] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000b9] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00172] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000ba] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00174] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000bb] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00176] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000bc] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00178] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000bd] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0017a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000be] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0017c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000bf] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0017e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000c0] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00180] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000c1] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00182] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000c2] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00184] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000c3] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00186] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000c4] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00188] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000c5] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0018a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000c6] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0018c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000c7] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0018e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000c8] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00190] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000c9] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00192] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000ca] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00194] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000cb] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00196] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000cc] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00198] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000cd] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0019a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000ce] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0019c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000cf] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0019e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000d0] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001a0] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000d1] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001a2] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000d2] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001a4] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000d3] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001a6] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000d4] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001a8] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000d5] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001aa] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000d6] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001ac] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000d7] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001ae] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000d8] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001b0] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000d9] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001b2] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000da] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001b4] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000db] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001b6] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000dc] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001b8] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000dd] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001ba] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000de] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001bc] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000df] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001be] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000e0] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001c0] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000e1] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001c2] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000e2] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001c4] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000e3] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001c6] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000e4] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001c8] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000e5] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001ca] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000e6] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001cc] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000e7] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001ce] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000e8] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001d0] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000e9] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001d2] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000ea] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001d4] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000eb] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001d6] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000ec] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001d8] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000ed] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001da] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000ee] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001dc] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000ef] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001de] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000f0] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001e0] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000f1] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001e2] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000f2] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001e4] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000f3] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001e6] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000f4] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001e8] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000f5] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001ea] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000f6] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001ec] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000f7] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001ee] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000f8] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001f0] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000f9] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001f2] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000fa] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001f4] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000fb] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001f6] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000fc] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001f8] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000fd] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001fa] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000fe] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001fc] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h000ff] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001fe] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00100] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00200] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00101] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00202] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00102] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00204] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00103] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00206] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00104] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00208] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00105] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0020a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00106] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0020c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00107] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0020e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00108] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00210] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00109] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00212] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0010a] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00214] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0010b] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00216] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0010c] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00218] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0010d] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0021a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0010e] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0021c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0010f] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0021e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00110] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00220] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00111] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00222] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00112] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00224] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00113] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00226] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00114] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00228] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00115] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0022a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00116] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0022c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00117] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0022e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00118] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00230] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00119] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00232] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0011a] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00234] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0011b] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00236] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0011c] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00238] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0011d] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0023a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0011e] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0023c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0011f] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0023e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00120] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00240] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00121] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00242] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00122] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00244] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00123] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00246] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00124] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00248] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00125] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0024a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00126] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0024c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00127] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0024e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00128] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00250] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00129] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00252] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0012a] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00254] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0012b] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00256] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0012c] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00258] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0012d] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0025a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0012e] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0025c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0012f] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0025e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00130] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00260] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00131] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00262] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00132] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00264] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00133] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00266] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00134] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00268] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00135] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0026a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00136] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0026c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00137] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0026e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00138] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00270] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00139] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00272] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0013a] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00274] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0013b] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00276] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0013c] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00278] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0013d] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0027a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0013e] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0027c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0013f] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0027e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00140] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00280] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00141] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00282] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00142] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00284] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00143] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00286] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00144] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00288] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00145] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0028a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00146] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0028c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00147] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0028e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00148] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00290] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00149] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00292] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0014a] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00294] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0014b] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00296] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0014c] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00298] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0014d] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0029a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0014e] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0029c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0014f] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0029e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00150] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002a0] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00151] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002a2] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00152] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002a4] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00153] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002a6] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00154] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002a8] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00155] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002aa] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00156] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002ac] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00157] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002ae] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00158] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002b0] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00159] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002b2] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0015a] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002b4] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0015b] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002b6] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0015c] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002b8] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0015d] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002ba] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0015e] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002bc] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0015f] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002be] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00160] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002c0] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00161] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002c2] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00162] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002c4] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00163] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002c6] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00164] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002c8] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00165] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002ca] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00166] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002cc] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00167] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002ce] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00168] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002d0] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00169] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002d2] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0016a] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002d4] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0016b] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002d6] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0016c] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002d8] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0016d] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002da] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0016e] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002dc] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0016f] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002de] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00170] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002e0] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00171] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002e2] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00172] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002e4] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00173] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002e6] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00174] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002e8] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00175] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002ea] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00176] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002ec] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00177] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002ee] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00178] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002f0] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00179] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002f2] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0017a] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002f4] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0017b] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002f6] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0017c] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002f8] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0017d] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002fa] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0017e] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002fc] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0017f] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002fe] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00180] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00300] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00181] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00302] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00182] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00304] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00183] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00306] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00184] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00308] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00185] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0030a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00186] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0030c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00187] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0030e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00188] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00310] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00189] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00312] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0018a] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00314] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0018b] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00316] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0018c] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00318] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0018d] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0031a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0018e] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0031c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0018f] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0031e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00190] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00320] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00191] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00322] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00192] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00324] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00193] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00326] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00194] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00328] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00195] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0032a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00196] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0032c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00197] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0032e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00198] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00330] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h00199] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00332] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0019a] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00334] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0019b] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00336] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0019c] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00338] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0019d] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0033a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0019e] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0033c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h0019f] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0033e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001a0] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00340] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001a1] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00342] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001a2] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00344] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001a3] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00346] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001a4] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00348] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001a5] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0034a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001a6] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0034c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001a7] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0034e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001a8] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00350] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001a9] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00352] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001aa] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00354] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001ab] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00356] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001ac] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00358] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001ad] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0035a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001ae] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0035c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001af] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0035e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001b0] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00360] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001b1] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00362] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001b2] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00364] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001b3] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00366] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001b4] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00368] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001b5] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0036a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001b6] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0036c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001b7] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0036e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001b8] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00370] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001b9] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00372] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001ba] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00374] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001bb] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00376] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001bc] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00378] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001bd] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0037a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001be] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0037c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001bf] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0037e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001c0] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00380] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001c1] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00382] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001c2] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00384] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001c3] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00386] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001c4] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00388] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001c5] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0038a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001c6] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0038c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001c7] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0038e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001c8] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00390] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001c9] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00392] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001ca] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00394] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001cb] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00396] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001cc] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00398] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001cd] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0039a] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001ce] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0039c] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001cf] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0039e] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001d0] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003a0] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001d1] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003a2] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001d2] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003a4] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001d3] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003a6] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001d4] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003a8] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001d5] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003aa] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001d6] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003ac] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001d7] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003ae] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001d8] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003b0] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001d9] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003b2] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001da] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003b4] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001db] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003b6] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001dc] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003b8] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001dd] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003ba] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001de] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003bc] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001df] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003be] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001e0] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003c0] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001e1] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003c2] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001e2] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003c4] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001e3] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003c6] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001e4] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003c8] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001e5] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003ca] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001e6] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003cc] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001e7] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003ce] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001e8] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003d0] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001e9] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003d2] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001ea] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003d4] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001eb] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003d6] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001ec] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003d8] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001ed] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003da] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001ee] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003dc] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001ef] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003de] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001f0] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003e0] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001f1] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003e2] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001f2] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003e4] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001f3] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003e6] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001f4] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003e8] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001f5] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003ea] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001f6] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003ec] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001f7] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003ee] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001f8] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003f0] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001f9] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003f2] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001fa] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003f4] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001fb] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003f6] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001fc] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003f8] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001fd] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003fa] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001fe] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003fc] ;
//end
//always_comb begin // 
               Ie40ac59fa3e2a4c35c71502fa3c82ebd96cb04e8e20dc3de3a4a223110fe38bd['h001ff] =  I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003fe] ;
//end
