 reg  ['h1ffff:0] [$clog2('h7000+1)-1:0] I3ce4b5a9d489daf4ff3697c7985730e1691281c16db6c67d16744b8a169a7716 ;
