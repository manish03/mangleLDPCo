 reg  ['h1ffff:0] [$clog2('h7000+1)-1:0] I9b16ca74bf83f6ffcaec2715f08644d43b958e8a67a64ef1326a2e3f8ba9a8a3 ;
