reg [flogtanh_WDTH -1:0] I9752ae2367e1a6c6f7352ea46ab95440, I6ceb8a53497c625c878b1bd0b10147d1;
reg [flogtanh_WDTH -1:0] I798dac490a694c8373633de0ebc4a72f, Iebd6f893703430ccce739c17a091180a;
reg [flogtanh_WDTH -1:0] I071022266cc4a3e5b31bfa3e084079d7, I87206f7a8f80c6791355b9e35fa789d4;
reg [flogtanh_WDTH -1:0] Ie1307d4ee93e9125654b49ccf5ead6b1, Ibeedd439ada9e1204f23f8b4c59d160e;
reg [flogtanh_WDTH -1:0] I880d7d200dbb730929b87b4936abb6b7, I722b96e8bbdedcbbf709b7ff75a343f2;
reg [flogtanh_WDTH -1:0] Ib692b0f0a9bd1601ef72ea3f12452a6a, Id82ca4ddd6bd7bd3eba9321f61fc83b1;
reg [flogtanh_WDTH -1:0] I697f7ccafe006697dd1aa6298a1cd9b7, I2cf927aba0ba024e37641e82687e3134;
reg [flogtanh_WDTH -1:0] I81006820f7f068a2ea7f42564c53345a, I0495eb40055242fe8d9886724a00437b;
reg [flogtanh_WDTH -1:0] Ic2dcdead9d2a2f6575fdec1ba1a2833c, Iaabf9a9cb8e18da9c94d145c54613499;
reg [flogtanh_WDTH -1:0] I88648891ecdf43525247de0259c99cb6, I9de00fb5f405754b7af66ab5206ee12c;
reg [flogtanh_WDTH -1:0] Ic4cfab074168cc1d247169480fdd03f6, I8f63c4af862af47948080677b089cc32;
reg [flogtanh_WDTH -1:0] I49b23654497581d82ca47a35e429a6ed, Iec915d0edfe90c0a3889228715277570;
reg [flogtanh_WDTH -1:0] I8f05a4f32582e13de9003ea0651b5e9f, I79f6ccccd78a7701f6302aab4293286c;
reg [flogtanh_WDTH -1:0] I317fe175f4bc5b04ed6b72d871974ef9, I90fe152dd5144845dd3b473f4cafb74e;
reg [flogtanh_WDTH -1:0] If84908bb6f231e3fad7d0f4cbab882de, I0bab994e09bb74cd97afe36943a98690;
reg [flogtanh_WDTH -1:0] I4f761cecb0e8b5c1bdab0e913cf3a798, Ic806ded37e428ee89a5725a3f0c69632;
reg [flogtanh_WDTH -1:0] Iaf08740a169f6f62bddfde35939f0e54, I1bb8a779c4c359bfc508d95a8d99c676;
reg [flogtanh_WDTH -1:0] I6577387fa85776dd6899c8b6fe15d202, Ic7037aee76219d7437fb16a34cd0575b;
reg [flogtanh_WDTH -1:0] Ib6958647f2dd08482fe95961b7f8dd09, I31653f719f0514a1e8b4dc749fa89eab;
reg [flogtanh_WDTH -1:0] I9ae8ddd960f78a4b6fcf14c9247a8ae5, Iee53e3dc893e03efc0d4f8b9e165a5df;
reg [flogtanh_WDTH -1:0] I7cef29b33735fd849743c3f06a82cba9, I12f3e3785de1cf141ea2c3efa11b6323;
reg [flogtanh_WDTH -1:0] I0cc3d5d926f4c45056afe4e02d652768, I415f363f69a1088c765e22738019ec87;
reg [flogtanh_WDTH -1:0] I1660f9dcac2e19e275df76b02173f49e, I3e72d56a69d40deafd501605f0257ac0;
reg [flogtanh_WDTH -1:0] I5c3b87e1908cc3d152b01573f7a87f2e, I6529b2ba884c7977f550cf3410db444d;
reg [flogtanh_WDTH -1:0] I302648ef72470338675f108cfc2936b0, If14fba2b2f70d2602b88ff0e739e113e;
reg [flogtanh_WDTH -1:0] I6e11ba6fced3ffc0d8f8003bf04bdfbf, I0685af82b58f41fa65efe1125fdaabeb;
reg [flogtanh_WDTH -1:0] Ia73537a3f8f0321742cdd459d952f4af, I1ad44f9d9abb2121b183a93dd1af4fa5;
reg [flogtanh_WDTH -1:0] I297ad7a97cf35acb5bfd1d0612044c49, I0f9dbc9aa169f7d63cc5789cb75c3a2d;
reg [flogtanh_WDTH -1:0] I712af4b1f576a39d2d96aff81da4863a, I5e458356e7698884ee785b2d5f1c368a;
reg [flogtanh_WDTH -1:0] I4a7d547601279634b9aaa30a51fbf741, I9b0f07f47267e3b0e0c545f44f5dd9f9;
reg [flogtanh_WDTH -1:0] Icec463cb0767bf054a74408bc41536b8, I3a4dd73e8b3f48746a991573531315dd;
reg [flogtanh_WDTH -1:0] I1ac433e960367e2ca78597357deb20a5, If727e9507d63727b0d597e9a5fee202a;
reg [flogtanh_WDTH -1:0] I7ca1e2fa8fc3e66fb6e747f2e0808e00, I9253bbcea2dc3a74433955d5f5aff705;
reg [flogtanh_WDTH -1:0] Id8930a77f5475a80411dfae4698cdfd8, Ibbabd657d00fc10d293b680d89593ca7;
reg [flogtanh_WDTH -1:0] Ifc5cdac396efc12756b713195f9fd57a, I79b7daae3f9f65acd3f79d579d2af25a;
reg [flogtanh_WDTH -1:0] I504e5446ead186c601225c6664e047c8, I74a4a1e449670380db8fbedbcf2aec04;
reg [flogtanh_WDTH -1:0] I8d9b55049a74bde1fdf26004008679a6, I9f7da2708edf4c941682b24f3999b159;
reg [flogtanh_WDTH -1:0] I155a7cee8b9f8b4d03f59ecde58fde8a, Id5d585b0c590354af34d02ba320f80d9;
reg [flogtanh_WDTH -1:0] I9cd50d02d3f7a189b5e70907ec8d1e73, Idab5b4bb4ed70dfe122f645eaf32852c;
reg [flogtanh_WDTH -1:0] I04a06a7a7af3891b0d53b95f24954344, Ic1793b6e075a12f6c1dda7e9fddc8b6e;
reg [flogtanh_WDTH -1:0] I21ea05b8f1be5a38bf4a4251644c370c, I168c51768b35b16f0033808f0b915e8c;
reg [flogtanh_WDTH -1:0] I89b558f53cd3391108aaee100bb68698, Ia7fa2fefde3f2ad6a0bee771a131219b;
reg [flogtanh_WDTH -1:0] I0b5cdc03696628bcb061aa2113444e50, I22d2ffb044bf579a2cccd3fcc70dae45;
reg [flogtanh_WDTH -1:0] I4293b2867a22e5f63df2ee4c19c88f79, Ib4b3cd8d5376f6ddb653c8cf72dceabf;
reg [flogtanh_WDTH -1:0] I966aa14cea82d7fd5872c135f0bbab70, I2c0b6e7a1fbcd97b6b78e65bf6d61213;
reg [flogtanh_WDTH -1:0] Id87f3e498747081eddc52a1fb671838d, Ifabbe9c31875e40eb81a87f0b19134e5;
reg [flogtanh_WDTH -1:0] Iabb62eea1f75ca64312cbb047714b9ca, Ic20259ce7eabae2029ca2ce312c6bfed;
reg [flogtanh_WDTH -1:0] Ie231dafa87260c19f1ac9c33085b94f4, Icaf0213b02a3cad251718b9ff86c108b;
reg [flogtanh_WDTH -1:0] Ief8246918e80c45898a4c38d0d5c3cbb, If71ff543c013f0111318a06039267570;
reg [flogtanh_WDTH -1:0] I574b308a0fd88d3f211b2acd576a3efb, I7871649505392bea882ad24b821c953c;
reg [flogtanh_WDTH -1:0] I8b32db6febf453df9d355666241b9a80, I5c4bcb5584cd15cbbec2709f29e15f36;
reg [flogtanh_WDTH -1:0] I7066424a4d00d757a4a0af28b0d95166, I73b98efd2185919a61b91a641fd6bdd7;
reg [flogtanh_WDTH -1:0] Ifc4d0343efb2e2f499cc6d8e37591f48, Ic2519d8c4e9b2c6f2126407a7a39fefe;
reg [flogtanh_WDTH -1:0] I1600115eb31dadcd5e87696ca1a34fbd, Ia806cdd7fbd6b44a8256aee7250ddd8b;
reg [flogtanh_WDTH -1:0] I5dce546007aab5da05bbd33b54ee3dba, I9badff60aa84397c6a408b846feceb91;
reg [flogtanh_WDTH -1:0] I6a5b90479676374b60fa668a358b852c, I885c54956c3ff7dfcd971f9d7ddf2db1;
reg [flogtanh_WDTH -1:0] Ieb0c46dc3852312024e2bf158d159f20, Ie3ae98a6abd28a3c39863a981e88e63f;
reg [flogtanh_WDTH -1:0] I56080da8b243334ef8414a095477c286, Ia1fed14f941d2ef3e78c490f81a5bd04;
reg [flogtanh_WDTH -1:0] I661a66590947450472c1cc6b8dc9239b, I714c5a8ac1480b08aa2859680ae40660;
reg [flogtanh_WDTH -1:0] Ie56fe9b766c784f90771d1335e397e99, I11d5e654536cd6b6e9b91487d76facb6;
reg [flogtanh_WDTH -1:0] Icaa6152af5f6bed3d595d51767c9ec49, I32f53cb8d864ff40c8d0ef95e9bdde54;
reg [flogtanh_WDTH -1:0] I99bddf2f101ab41147b2849d22bd8e0c, I0c3874311a119530873f475b01006dd4;
reg [flogtanh_WDTH -1:0] I5ef97e1962a901d1e6557c0dfcae036e, I585684cf3ba45f359e0f0752e9e88819;
reg [flogtanh_WDTH -1:0] I3e1118befba3c769deb7bbf9d1875d00, I998f8a35c7ec923067dc75c76c9df713;
reg [flogtanh_WDTH -1:0] I435152993799746e1f967343ce1b106f, I4e8f27bdc42f1e3f4024b020d5821dff;
reg [flogtanh_WDTH -1:0] I9e10d71db16be96b3087a3a584a5b55b, I93f0932897b358b6c4e3386609cffa36;
reg [flogtanh_WDTH -1:0] Ic943175727986874531ace57f5697df3, I9ae8e176f8f34220d2cac97abe1fd32a;
reg [flogtanh_WDTH -1:0] I18d1d32d1e58254b964c670e0d83c119, I7fdc9543e6c7c0324293936b1c2c8f2d;
reg [flogtanh_WDTH -1:0] I96b27127bbc15301b57d83982260853b, Ic9bc7816fcb1f128d833fde39ad8cf1d;
reg [flogtanh_WDTH -1:0] I12d97a28ef39f26eb4996aa2f1d9eafb, Ifd16243bd087b16c5bfa2bfbb8239ee1;
reg [flogtanh_WDTH -1:0] Iddafd4529ad594eda9835e76efa116bb, I3479e7931017ab45aa4e99ca34b8b5cb;
reg [flogtanh_WDTH -1:0] Ice9aeaff41b923556b30553d8b42da47, I7cf57ee976846690c3286f08ef932683;
reg [flogtanh_WDTH -1:0] I33e7dfa55b2d2ac83a8f57797fcd68db, I32769b7f105065785745633dfef8a4c5;
reg [flogtanh_WDTH -1:0] I5c3dedd601ffa33d7b649b2c08df54e6, I47e2d27cbd69c85106a4aa3ac2784eb0;
reg [flogtanh_WDTH -1:0] I1660ea57c727ecd6e71a4e9c4c288b45, Ibd0efa281371fa3b94eed5e021c73642;
reg [flogtanh_WDTH -1:0] I1c9e513f7524f52e24e7e80807a18ac6, I82aaeb65a83948cd75521499d2719001;
reg [flogtanh_WDTH -1:0] I3d1372ff9b830f5eeb50c4e47d322cf7, If9854de536b8ba1392ba0328ef7cebba;
reg [flogtanh_WDTH -1:0] I69460735237cd5bd0f26254f6f32e357, I731416642a03748ca4698a73e094c500;
reg [flogtanh_WDTH -1:0] Iac63249f3101e957234cb4efee5f6771, I23c90590a514d430c9828af570ebf16a;
reg [flogtanh_WDTH -1:0] I769cf83f4404ee0d85e6c13b7d0c737b, I2d07aa91cf23a7789428c96e4f73109e;
reg [flogtanh_WDTH -1:0] Ieff66b38feb970b4ab3006fb31e5cce3, I89fc8a2a491dcc20f2556e7042d22384;
reg [flogtanh_WDTH -1:0] Ifbef84b3392347c7e0e52e232d26f9bd, I0f76a71ea70551bbf89f01a689811954;
reg [flogtanh_WDTH -1:0] I13989f78ab3eab13b7f0619fb0386e3d, I0b6ce8e59afb2e48df79fefd5450971e;
reg [flogtanh_WDTH -1:0] I61af8fbc53b6f763a8b77012fb56be23, I35a8c09862db36ffde26d27b74baa8ba;
reg [flogtanh_WDTH -1:0] Id0969f699976b1041d15d62912a04b5f, I920593851f5860485fd105f8d4c1b8c9;
reg [flogtanh_WDTH -1:0] I3be47f6dae15615b1b6b0cb52bb8cd5a, I51dcc6894ba28567c3077ea409871161;
reg [flogtanh_WDTH -1:0] Iabe728226ae671218667d92139083a4c, I79489994f40f88e0b5a8a8be6322f3ec;
reg [flogtanh_WDTH -1:0] I49d60f1269fcc5a98196ac391823ca1a, I6503341e5d6ced0d71bd29bbc622020b;
reg [flogtanh_WDTH -1:0] Ic88cdb92bf89df187d801b480c7c2770, I178d103fabf53395ce88cdbfc14917ce;
reg [flogtanh_WDTH -1:0] I60a972d5f2465dd5f9c3665eee4cffc2, I3a8d57af0e6ed1437d572534742a9f2f;
reg [flogtanh_WDTH -1:0] Iaafcf98c2c079884e32f2bd70972e5b3, I4602a0caf02e37e360e5cf9de1003cd2;
reg [flogtanh_WDTH -1:0] I3c4a90a70e7cfe814427262cae88e2a6, I245a6df9f9d730338cd52169a3f466d3;
reg [flogtanh_WDTH -1:0] I7eb2363c8fe8f49f839b59df19165aab, Ia7a8ebe681523a490c83dcb84ac82a2a;
reg [flogtanh_WDTH -1:0] I60bf9f27a86ec731795d79b656e2229c, I7caf04f8880b455d92307bf521540c38;
reg [flogtanh_WDTH -1:0] I8d4fa08cc0155e81bb2ce4ab9a39df4a, I401eb53331986f8474c861acb2b2a445;
reg [flogtanh_WDTH -1:0] Ie21b4ae619493ef57536508645aa29bb, If3e4f18a03ca4b7b1d89ef842c68e96d;
reg [flogtanh_WDTH -1:0] I854fac49e7921a59773ab612181b9569, I0d6bc03eddef33a7d70ac2cc27049107;
reg [flogtanh_WDTH -1:0] I20a9b10f04d9eeca6058889d5c930294, I2214bdaf7568fd3c20109ead1daf861d;
reg [flogtanh_WDTH -1:0] I122fde74534a82953b1a5a476e2e8151, I6138bf9b2a35f3b08f216eeaf3c0ebee;
reg [flogtanh_WDTH -1:0] Ia535aa71b5100fd37cb15ba1612d2d52, Ibd3927f27dbf4a60128f60f31b5a32e6;
reg [flogtanh_WDTH -1:0] I8b588d7b4605f968fd007ed894b4ee68, I26faa75fc5dd15baf23481311b220832;
reg [flogtanh_WDTH -1:0] I88d97aa0544a09e2a0df10ec0a57ea54, I373328eb3cc59c5d3d7a5102535c5410;
reg [flogtanh_WDTH -1:0] I81cb66f14210612d88911543c3517731, I1bb3c77cdfd0b229bbdf7b33fd4a613c;
reg [flogtanh_WDTH -1:0] Ibd10299291ec40ff247b816be64f07ec, Ia1c8178574520829f24c8cc08e15e8f1;
reg [flogtanh_WDTH -1:0] I3e4ecb5c8164f70ca4b16eb004cb276c, Ib911176056f3c0378dfa8a77e0c5b69a;
reg [flogtanh_WDTH -1:0] Id5e6fca7b1cebfd4f2caf7465fb678fa, If9afa8946804ce9c74ef43d3ca669849;
reg [flogtanh_WDTH -1:0] I58a570689c10954778a3e3ded8d4f9b4, I6bb576223350a8373e430d185efe7fd9;
reg [flogtanh_WDTH -1:0] I0a8dea5e3f82d6954d294cf3c3c858d2, Id7008a8f0d70f1e23a073745ed4a57c0;
reg [flogtanh_WDTH -1:0] I9aea2a89a8d17d14da2fccad570cfc7d, I87e0bcba46bcc28ad02b7e0af773d82a;
reg [flogtanh_WDTH -1:0] I8b661503122504ce012fe534dad9c394, I3bb6f388db8c8dc2b6c963749ef48096;
reg [flogtanh_WDTH -1:0] Ib9a8e5b5096d6c5ed5cc315a5899b8d5, Iea2bbf25e38901d15434dfc83d65ada4;
reg [flogtanh_WDTH -1:0] Iebf5cd787ff1d73dfbe4e52cfbaffc14, Ie5e331564633cd16934cd0714b2953cb;
reg [flogtanh_WDTH -1:0] I4096de17c18f5e0af8d288bc6887c6cb, Ibcc6c8744ee9a2ad9766c0f9fa196036;
reg [flogtanh_WDTH -1:0] I949e53f68343283236a519295c606cc2, Ic425c518a69f3f85e219b1f15baa5d36;
reg [flogtanh_WDTH -1:0] Id9fc0dbdd3cd0709ef28238589312443, I78ba7a5627868f3c0b75555131470aa4;
reg [flogtanh_WDTH -1:0] Idf5ff15e65f46f3b569ef0d634cd5819, I3b5bd630c8d2bdb455b6f75a6a8a4a53;
reg [flogtanh_WDTH -1:0] I3d70051f81db3db896a8455dda9f0022, I4274a587dd459b29ecee1ff1554a12f7;
reg [flogtanh_WDTH -1:0] I737715c7b75b324dca40210b708166ac, I9728cc3e93018b67d2c2e94f9d90f433;
reg [flogtanh_WDTH -1:0] I3deb95e95d3308de220901f8fe6d2ee4, If77d0921ff0a38d2b3fcd28c5be4a131;
reg [flogtanh_WDTH -1:0] I5e7775e3bc484bed7a57f04b0cd7ccca, I29046786efe54344e3cffb3e5e913667;
reg [flogtanh_WDTH -1:0] Ic557aa69aa946711cc39627fe6133f87, I6fbdabe9ecefa8648c4ca4ec51e251a4;
reg [flogtanh_WDTH -1:0] I004142a2c8e12e72c3ac4a439b281fcc, Ia456c9d3e431416da7685ea0c42371f9;
reg [flogtanh_WDTH -1:0] Ia112b4cab1631793a8cc6291027c616c, Ib68b82bab62a694692b3fd2191b5f29c;
reg [flogtanh_WDTH -1:0] I3d3a0cda05e77a00523ea3f4aae38d82, Iacfc43c384ab56bf924d5ae09a59fb17;
reg [flogtanh_WDTH -1:0] I723f34fa0b35af4e77fbecc65d2ca88b, Id5c5e697446d9974b383880138f73778;
reg [flogtanh_WDTH -1:0] I460bbb250271f3fa5414de2e68474fbc, I441c5f07ae7d849600f2d02cc5753d5a;
reg [flogtanh_WDTH -1:0] I1e29e4b5d18509694df3a0e7b7cd2a7d, Ic117c98ae21f7640aa5a68539ec03821;
reg [flogtanh_WDTH -1:0] Ie25c961fe6b06030e848c7b9eb751909, I4c3f1b807cae7d5a4a5dcd3c8180c0fe;
reg [flogtanh_WDTH -1:0] I16c56d8b22dd23fbb09ebf4f36107cc9, Idc31f916f132a0c203eb03a7d1de62bb;
reg [flogtanh_WDTH -1:0] I1e10a4b5844d25334b74e1088e2d3deb, I68ae757abeedcaee5336b7d45a29b8c7;
reg [flogtanh_WDTH -1:0] Ic524b9ac09a3499b67313edee303c53f, I5e4276800e079f48c3953f01869bcfa0;
reg [flogtanh_WDTH -1:0] Ie332a236ba72fed22c9d7670390dc3d1, I30254925c90cc28a13afa22e983854bb;
reg [flogtanh_WDTH -1:0] Ia04ae82f80fd35c0eb30fd17ec9f74a2, I5955344e0f04e1ddf15eecf2eede2346;
reg [flogtanh_WDTH -1:0] I009b2657f941367412da0645c61a6161, I82b8db69079237f10477ebd39a13bc16;
reg [flogtanh_WDTH -1:0] If84fc94571af2905f59753301bfb7fec, I83df9b9b4dc9b0eeaf05f25e513d1603;
reg [flogtanh_WDTH -1:0] I782050339f5fcecb44819e7cb6dac5d6, I54e2da03e41cfdd43ca24929ef467819;
reg [flogtanh_WDTH -1:0] I5ce602af9806ed123e70480c643be643, I5b3e2ec3e81cfbb4cff4a55faf1779ce;
reg [flogtanh_WDTH -1:0] Id2450e8bc8cad7c46f1d47372a344f12, Ib5d40f3069e5a3e1da68013a7f5e640d;
reg [flogtanh_WDTH -1:0] Id074a700da35c1548c27b5d1c7e9eea0, Iecc3e2589b1a21ad89360386cbc59203;
reg [flogtanh_WDTH -1:0] I689e819fcdc296cb4b537538012615f6, Ia4d367afebe196ee6debdda4251771b6;
reg [flogtanh_WDTH -1:0] Ic2824f1963f1158e7ad33e9c81bc7d08, Ibce5b55e9f3477e8cac134660f3e056d;
reg [flogtanh_WDTH -1:0] Id0ae33a482904b109068ad943d76d758, I5f2c9622ecb56c3385f986e11cda6344;
reg [flogtanh_WDTH -1:0] I7b7386e46768f03c912485c3c80065dc, Ic95be5fcb699a68e0e796dc0408fd5f3;
reg [flogtanh_WDTH -1:0] Ib0e71935bab4a9ebf00d9b2d170b571a, I01c4e6856aaa370540e370d30223a3e9;
reg [flogtanh_WDTH -1:0] I4613dca4c7c67e9dffb22110f62d93a1, I693343088a46766b65b21833e8c93424;
reg [flogtanh_WDTH -1:0] Ifc0a83912f31329972ce02109fe40df0, I363bfe5c6d747f1b0bf3b3795973cc1a;
reg [flogtanh_WDTH -1:0] I021270a1b11bc14783313a27684e1a08, Ibcd20a65390727b99272e778f6b5cd48;
reg [flogtanh_WDTH -1:0] I0f8f6a239a05dba04dd3b845c9e8ac9b, I824e45de28b3352d3189623ca276ceb4;
reg [flogtanh_WDTH -1:0] I99d616bf2017cd8e4f019fa9356a4c9f, Iee99e323224f79b59ff094ca4e0b730f;
reg [flogtanh_WDTH -1:0] I48c538d54789fc85a7349065dc33b20d, Id6c903e77c0ae87fc00b0a19926eac0d;
reg [flogtanh_WDTH -1:0] Idf3ebc5f6ef593255d94f70583e028ba, Icf2d8147505a677d965332527efd32e5;
reg [flogtanh_WDTH -1:0] I5ec053664237ddc305a831b20239a5b3, I10edceddaabd0b5704cfe32642099bfc;
reg [flogtanh_WDTH -1:0] I2150bffc35644044c52346accf50c6a6, I7af4f3f04f52198149fab343b09a7c33;
reg [flogtanh_WDTH -1:0] I9a16fe81b2e09494fb280b564b2d8447, I5b772125b565150758a1dd9173661a69;
reg [flogtanh_WDTH -1:0] I3a78158e0bcd94e117696bd698f00e43, I8d3688317aaf1a973e53e7d82c07aff5;
reg [flogtanh_WDTH -1:0] Ia674fb4751c28067672ed365648d4046, Id1bd6b209ebbc1dc87ef765e8311d13d;
reg [flogtanh_WDTH -1:0] I7c2f789de92dcd3106cd534d547ff653, I2145db99a9f07a8dcca7bb21537c3c6b;
reg [flogtanh_WDTH -1:0] I42484fc96375ed4f28054b45a7a573a4, I0578f5f40c3743a4c0184768a6842378;
reg [flogtanh_WDTH -1:0] Ife0e6d58f356f10d7f769f225de5a7cc, Ia36d890f9c568613260b96683ad1442e;
reg [flogtanh_WDTH -1:0] Id958719d49aab2d0b082a6d24fe4c3ed, Idd923fa51da8d881654d1a0b2939bf45;
reg [flogtanh_WDTH -1:0] I6f030649ec413f3a8b1b2818f11fdeb9, I83e8203369eabb1165454d054fc6368a;
reg [flogtanh_WDTH -1:0] I1b4cbdf5cfa3d8c53d2000918dab9d92, I811bb1c2a735a7b3b494db92a6e09bc1;
reg [flogtanh_WDTH -1:0] Id48425985a33f1512c0dd32361ceb85e, I2cf7c8df11a71a3952a5c11fce1ab746;
reg [flogtanh_WDTH -1:0] I37d45d42016be2e2bc96ae6fd4287f97, Ic219b4e5b38cf27b7c30f1b1455db7c1;
reg [flogtanh_WDTH -1:0] I6715c7f4ac584103721a33ead7ed395b, I964950b31cf4117e79e46a2282faf273;
reg [flogtanh_WDTH -1:0] Ia8e9d2fd6a51de4383c16a35737a1831, Ic4ddd59bdd32e1c8481e7d39707d2628;
reg [flogtanh_WDTH -1:0] I3efa217d3d93a9a2f15bdcd906a2a230, I754ed93d8e7f3ed1b9bbf1aa0a780631;
reg [flogtanh_WDTH -1:0] I016707bf26cc19976929a8b14f535455, Ieb469f605aef6bb6cc19088b0a8d191e;
reg [flogtanh_WDTH -1:0] I698072a5328a85b0b22ec7bc94b8372e, I0be6033ae52cefc976cf28e9c6972b2c;
reg [flogtanh_WDTH -1:0] I70a428ae2a62212ed93be37b860e8231, I913ad4107114014e726ae5a684208f1f;
reg [flogtanh_WDTH -1:0] I5193a317b4c9d2bf1992ca5cf9936681, I332be99f2c509a0ad9ce2003f3894900;
reg [flogtanh_WDTH -1:0] I9cb0c1a404a77903890379f0f658c70a, If615b5edf5772640f5e7db1b7c2b827e;
reg [flogtanh_WDTH -1:0] I861bb6fa26ecdc43776d01811abe7bc3, Ic98c3c04426af7540b59e85693f8c85e;
reg [flogtanh_WDTH -1:0] I92ad6f4d3a62fbd3e86cda7457115093, Ia8b37c51a90549caefe7c587af95efcf;
reg [flogtanh_WDTH -1:0] I17f6c0345023a3824d5e40506e4c1919, Ie34547c669ac94c6b215f01c235086e4;
reg [flogtanh_WDTH -1:0] Ic309d272e0e79647de87c07aae1e798c, Ibed1e35fd09ac08952020a915b52aae9;
reg [flogtanh_WDTH -1:0] I24a4c216e917b9b9ad744c7bfa4a7d24, I27def56001fb56e6a85c9c61ba8d55bd;
reg [flogtanh_WDTH -1:0] I7112d906a2a8245dd62b7ef26d7e54ee, I6540e74c5f9178782a17fe7460aaf4ee;
reg Icf92b5275d264e1b6d832272a0d01a66 ;
always @(posedge clk or negedge rstn)
if (!rstn) begin
 I6ceb8a53497c625c878b1bd0b10147d1 <= 'h0;
 Iebd6f893703430ccce739c17a091180a <= 'h0;
 I87206f7a8f80c6791355b9e35fa789d4 <= 'h0;
 Ibeedd439ada9e1204f23f8b4c59d160e <= 'h0;
 I722b96e8bbdedcbbf709b7ff75a343f2 <= 'h0;
 Id82ca4ddd6bd7bd3eba9321f61fc83b1 <= 'h0;
 I2cf927aba0ba024e37641e82687e3134 <= 'h0;
 I0495eb40055242fe8d9886724a00437b <= 'h0;
 Iaabf9a9cb8e18da9c94d145c54613499 <= 'h0;
 I9de00fb5f405754b7af66ab5206ee12c <= 'h0;
 I8f63c4af862af47948080677b089cc32 <= 'h0;
 Iec915d0edfe90c0a3889228715277570 <= 'h0;
 I79f6ccccd78a7701f6302aab4293286c <= 'h0;
 I90fe152dd5144845dd3b473f4cafb74e <= 'h0;
 I0bab994e09bb74cd97afe36943a98690 <= 'h0;
 Ic806ded37e428ee89a5725a3f0c69632 <= 'h0;
 I1bb8a779c4c359bfc508d95a8d99c676 <= 'h0;
 Ic7037aee76219d7437fb16a34cd0575b <= 'h0;
 I31653f719f0514a1e8b4dc749fa89eab <= 'h0;
 Iee53e3dc893e03efc0d4f8b9e165a5df <= 'h0;
 I12f3e3785de1cf141ea2c3efa11b6323 <= 'h0;
 I415f363f69a1088c765e22738019ec87 <= 'h0;
 I3e72d56a69d40deafd501605f0257ac0 <= 'h0;
 I6529b2ba884c7977f550cf3410db444d <= 'h0;
 If14fba2b2f70d2602b88ff0e739e113e <= 'h0;
 I0685af82b58f41fa65efe1125fdaabeb <= 'h0;
 I1ad44f9d9abb2121b183a93dd1af4fa5 <= 'h0;
 I0f9dbc9aa169f7d63cc5789cb75c3a2d <= 'h0;
 I5e458356e7698884ee785b2d5f1c368a <= 'h0;
 I9b0f07f47267e3b0e0c545f44f5dd9f9 <= 'h0;
 I3a4dd73e8b3f48746a991573531315dd <= 'h0;
 If727e9507d63727b0d597e9a5fee202a <= 'h0;
 I9253bbcea2dc3a74433955d5f5aff705 <= 'h0;
 Ibbabd657d00fc10d293b680d89593ca7 <= 'h0;
 I79b7daae3f9f65acd3f79d579d2af25a <= 'h0;
 I74a4a1e449670380db8fbedbcf2aec04 <= 'h0;
 I9f7da2708edf4c941682b24f3999b159 <= 'h0;
 Id5d585b0c590354af34d02ba320f80d9 <= 'h0;
 Idab5b4bb4ed70dfe122f645eaf32852c <= 'h0;
 Ic1793b6e075a12f6c1dda7e9fddc8b6e <= 'h0;
 I168c51768b35b16f0033808f0b915e8c <= 'h0;
 Ia7fa2fefde3f2ad6a0bee771a131219b <= 'h0;
 I22d2ffb044bf579a2cccd3fcc70dae45 <= 'h0;
 Ib4b3cd8d5376f6ddb653c8cf72dceabf <= 'h0;
 I2c0b6e7a1fbcd97b6b78e65bf6d61213 <= 'h0;
 Ifabbe9c31875e40eb81a87f0b19134e5 <= 'h0;
 Ic20259ce7eabae2029ca2ce312c6bfed <= 'h0;
 Icaf0213b02a3cad251718b9ff86c108b <= 'h0;
 If71ff543c013f0111318a06039267570 <= 'h0;
 I7871649505392bea882ad24b821c953c <= 'h0;
 I5c4bcb5584cd15cbbec2709f29e15f36 <= 'h0;
 I73b98efd2185919a61b91a641fd6bdd7 <= 'h0;
 Ic2519d8c4e9b2c6f2126407a7a39fefe <= 'h0;
 Ia806cdd7fbd6b44a8256aee7250ddd8b <= 'h0;
 I9badff60aa84397c6a408b846feceb91 <= 'h0;
 I885c54956c3ff7dfcd971f9d7ddf2db1 <= 'h0;
 Ie3ae98a6abd28a3c39863a981e88e63f <= 'h0;
 Ia1fed14f941d2ef3e78c490f81a5bd04 <= 'h0;
 I714c5a8ac1480b08aa2859680ae40660 <= 'h0;
 I11d5e654536cd6b6e9b91487d76facb6 <= 'h0;
 I32f53cb8d864ff40c8d0ef95e9bdde54 <= 'h0;
 I0c3874311a119530873f475b01006dd4 <= 'h0;
 I585684cf3ba45f359e0f0752e9e88819 <= 'h0;
 I998f8a35c7ec923067dc75c76c9df713 <= 'h0;
 I4e8f27bdc42f1e3f4024b020d5821dff <= 'h0;
 I93f0932897b358b6c4e3386609cffa36 <= 'h0;
 I9ae8e176f8f34220d2cac97abe1fd32a <= 'h0;
 I7fdc9543e6c7c0324293936b1c2c8f2d <= 'h0;
 Ic9bc7816fcb1f128d833fde39ad8cf1d <= 'h0;
 Ifd16243bd087b16c5bfa2bfbb8239ee1 <= 'h0;
 I3479e7931017ab45aa4e99ca34b8b5cb <= 'h0;
 I7cf57ee976846690c3286f08ef932683 <= 'h0;
 I32769b7f105065785745633dfef8a4c5 <= 'h0;
 I47e2d27cbd69c85106a4aa3ac2784eb0 <= 'h0;
 Ibd0efa281371fa3b94eed5e021c73642 <= 'h0;
 I82aaeb65a83948cd75521499d2719001 <= 'h0;
 If9854de536b8ba1392ba0328ef7cebba <= 'h0;
 I731416642a03748ca4698a73e094c500 <= 'h0;
 I23c90590a514d430c9828af570ebf16a <= 'h0;
 I2d07aa91cf23a7789428c96e4f73109e <= 'h0;
 I89fc8a2a491dcc20f2556e7042d22384 <= 'h0;
 I0f76a71ea70551bbf89f01a689811954 <= 'h0;
 I0b6ce8e59afb2e48df79fefd5450971e <= 'h0;
 I35a8c09862db36ffde26d27b74baa8ba <= 'h0;
 I920593851f5860485fd105f8d4c1b8c9 <= 'h0;
 I51dcc6894ba28567c3077ea409871161 <= 'h0;
 I79489994f40f88e0b5a8a8be6322f3ec <= 'h0;
 I6503341e5d6ced0d71bd29bbc622020b <= 'h0;
 I178d103fabf53395ce88cdbfc14917ce <= 'h0;
 I3a8d57af0e6ed1437d572534742a9f2f <= 'h0;
 I4602a0caf02e37e360e5cf9de1003cd2 <= 'h0;
 I245a6df9f9d730338cd52169a3f466d3 <= 'h0;
 Ia7a8ebe681523a490c83dcb84ac82a2a <= 'h0;
 I7caf04f8880b455d92307bf521540c38 <= 'h0;
 I401eb53331986f8474c861acb2b2a445 <= 'h0;
 If3e4f18a03ca4b7b1d89ef842c68e96d <= 'h0;
 I0d6bc03eddef33a7d70ac2cc27049107 <= 'h0;
 I2214bdaf7568fd3c20109ead1daf861d <= 'h0;
 I6138bf9b2a35f3b08f216eeaf3c0ebee <= 'h0;
 Ibd3927f27dbf4a60128f60f31b5a32e6 <= 'h0;
 I26faa75fc5dd15baf23481311b220832 <= 'h0;
 I373328eb3cc59c5d3d7a5102535c5410 <= 'h0;
 I1bb3c77cdfd0b229bbdf7b33fd4a613c <= 'h0;
 Ia1c8178574520829f24c8cc08e15e8f1 <= 'h0;
 Ib911176056f3c0378dfa8a77e0c5b69a <= 'h0;
 If9afa8946804ce9c74ef43d3ca669849 <= 'h0;
 I6bb576223350a8373e430d185efe7fd9 <= 'h0;
 Id7008a8f0d70f1e23a073745ed4a57c0 <= 'h0;
 I87e0bcba46bcc28ad02b7e0af773d82a <= 'h0;
 I3bb6f388db8c8dc2b6c963749ef48096 <= 'h0;
 Iea2bbf25e38901d15434dfc83d65ada4 <= 'h0;
 Ie5e331564633cd16934cd0714b2953cb <= 'h0;
 Ibcc6c8744ee9a2ad9766c0f9fa196036 <= 'h0;
 Ic425c518a69f3f85e219b1f15baa5d36 <= 'h0;
 I78ba7a5627868f3c0b75555131470aa4 <= 'h0;
 I3b5bd630c8d2bdb455b6f75a6a8a4a53 <= 'h0;
 I4274a587dd459b29ecee1ff1554a12f7 <= 'h0;
 I9728cc3e93018b67d2c2e94f9d90f433 <= 'h0;
 If77d0921ff0a38d2b3fcd28c5be4a131 <= 'h0;
 I29046786efe54344e3cffb3e5e913667 <= 'h0;
 I6fbdabe9ecefa8648c4ca4ec51e251a4 <= 'h0;
 Ia456c9d3e431416da7685ea0c42371f9 <= 'h0;
 Ib68b82bab62a694692b3fd2191b5f29c <= 'h0;
 Iacfc43c384ab56bf924d5ae09a59fb17 <= 'h0;
 Id5c5e697446d9974b383880138f73778 <= 'h0;
 I441c5f07ae7d849600f2d02cc5753d5a <= 'h0;
 Ic117c98ae21f7640aa5a68539ec03821 <= 'h0;
 I4c3f1b807cae7d5a4a5dcd3c8180c0fe <= 'h0;
 Idc31f916f132a0c203eb03a7d1de62bb <= 'h0;
 I68ae757abeedcaee5336b7d45a29b8c7 <= 'h0;
 I5e4276800e079f48c3953f01869bcfa0 <= 'h0;
 I30254925c90cc28a13afa22e983854bb <= 'h0;
 I5955344e0f04e1ddf15eecf2eede2346 <= 'h0;
 I82b8db69079237f10477ebd39a13bc16 <= 'h0;
 I83df9b9b4dc9b0eeaf05f25e513d1603 <= 'h0;
 I54e2da03e41cfdd43ca24929ef467819 <= 'h0;
 I5b3e2ec3e81cfbb4cff4a55faf1779ce <= 'h0;
 Ib5d40f3069e5a3e1da68013a7f5e640d <= 'h0;
 Iecc3e2589b1a21ad89360386cbc59203 <= 'h0;
 Ia4d367afebe196ee6debdda4251771b6 <= 'h0;
 Ibce5b55e9f3477e8cac134660f3e056d <= 'h0;
 I5f2c9622ecb56c3385f986e11cda6344 <= 'h0;
 Ic95be5fcb699a68e0e796dc0408fd5f3 <= 'h0;
 I01c4e6856aaa370540e370d30223a3e9 <= 'h0;
 I693343088a46766b65b21833e8c93424 <= 'h0;
 I363bfe5c6d747f1b0bf3b3795973cc1a <= 'h0;
 Ibcd20a65390727b99272e778f6b5cd48 <= 'h0;
 I824e45de28b3352d3189623ca276ceb4 <= 'h0;
 Iee99e323224f79b59ff094ca4e0b730f <= 'h0;
 Id6c903e77c0ae87fc00b0a19926eac0d <= 'h0;
 Icf2d8147505a677d965332527efd32e5 <= 'h0;
 I10edceddaabd0b5704cfe32642099bfc <= 'h0;
 I7af4f3f04f52198149fab343b09a7c33 <= 'h0;
 I5b772125b565150758a1dd9173661a69 <= 'h0;
 I8d3688317aaf1a973e53e7d82c07aff5 <= 'h0;
 Id1bd6b209ebbc1dc87ef765e8311d13d <= 'h0;
 I2145db99a9f07a8dcca7bb21537c3c6b <= 'h0;
 I0578f5f40c3743a4c0184768a6842378 <= 'h0;
 Ia36d890f9c568613260b96683ad1442e <= 'h0;
 Idd923fa51da8d881654d1a0b2939bf45 <= 'h0;
 I83e8203369eabb1165454d054fc6368a <= 'h0;
 I811bb1c2a735a7b3b494db92a6e09bc1 <= 'h0;
 I2cf7c8df11a71a3952a5c11fce1ab746 <= 'h0;
 Ic219b4e5b38cf27b7c30f1b1455db7c1 <= 'h0;
 I964950b31cf4117e79e46a2282faf273 <= 'h0;
 Ic4ddd59bdd32e1c8481e7d39707d2628 <= 'h0;
 I754ed93d8e7f3ed1b9bbf1aa0a780631 <= 'h0;
 Ieb469f605aef6bb6cc19088b0a8d191e <= 'h0;
 I0be6033ae52cefc976cf28e9c6972b2c <= 'h0;
 I913ad4107114014e726ae5a684208f1f <= 'h0;
 I332be99f2c509a0ad9ce2003f3894900 <= 'h0;
 If615b5edf5772640f5e7db1b7c2b827e <= 'h0;
 Ic98c3c04426af7540b59e85693f8c85e <= 'h0;
 Ia8b37c51a90549caefe7c587af95efcf <= 'h0;
 Ie34547c669ac94c6b215f01c235086e4 <= 'h0;
 Ibed1e35fd09ac08952020a915b52aae9 <= 'h0;
 I27def56001fb56e6a85c9c61ba8d55bd <= 'h0;
 I6540e74c5f9178782a17fe7460aaf4ee <= 'h0;
 Icf92b5275d264e1b6d832272a0d01a66 <= 'h0;
end
else
begin
 I6ceb8a53497c625c878b1bd0b10147d1 <=  I9752ae2367e1a6c6f7352ea46ab95440;
 Iebd6f893703430ccce739c17a091180a <=  I798dac490a694c8373633de0ebc4a72f;
 I87206f7a8f80c6791355b9e35fa789d4 <=  I071022266cc4a3e5b31bfa3e084079d7;
 Ibeedd439ada9e1204f23f8b4c59d160e <=  Ie1307d4ee93e9125654b49ccf5ead6b1;
 I722b96e8bbdedcbbf709b7ff75a343f2 <=  I880d7d200dbb730929b87b4936abb6b7;
 Id82ca4ddd6bd7bd3eba9321f61fc83b1 <=  Ib692b0f0a9bd1601ef72ea3f12452a6a;
 I2cf927aba0ba024e37641e82687e3134 <=  I697f7ccafe006697dd1aa6298a1cd9b7;
 I0495eb40055242fe8d9886724a00437b <=  I81006820f7f068a2ea7f42564c53345a;
 Iaabf9a9cb8e18da9c94d145c54613499 <=  Ic2dcdead9d2a2f6575fdec1ba1a2833c;
 I9de00fb5f405754b7af66ab5206ee12c <=  I88648891ecdf43525247de0259c99cb6;
 I8f63c4af862af47948080677b089cc32 <=  Ic4cfab074168cc1d247169480fdd03f6;
 Iec915d0edfe90c0a3889228715277570 <=  I49b23654497581d82ca47a35e429a6ed;
 I79f6ccccd78a7701f6302aab4293286c <=  I8f05a4f32582e13de9003ea0651b5e9f;
 I90fe152dd5144845dd3b473f4cafb74e <=  I317fe175f4bc5b04ed6b72d871974ef9;
 I0bab994e09bb74cd97afe36943a98690 <=  If84908bb6f231e3fad7d0f4cbab882de;
 Ic806ded37e428ee89a5725a3f0c69632 <=  I4f761cecb0e8b5c1bdab0e913cf3a798;
 I1bb8a779c4c359bfc508d95a8d99c676 <=  Iaf08740a169f6f62bddfde35939f0e54;
 Ic7037aee76219d7437fb16a34cd0575b <=  I6577387fa85776dd6899c8b6fe15d202;
 I31653f719f0514a1e8b4dc749fa89eab <=  Ib6958647f2dd08482fe95961b7f8dd09;
 Iee53e3dc893e03efc0d4f8b9e165a5df <=  I9ae8ddd960f78a4b6fcf14c9247a8ae5;
 I12f3e3785de1cf141ea2c3efa11b6323 <=  I7cef29b33735fd849743c3f06a82cba9;
 I415f363f69a1088c765e22738019ec87 <=  I0cc3d5d926f4c45056afe4e02d652768;
 I3e72d56a69d40deafd501605f0257ac0 <=  I1660f9dcac2e19e275df76b02173f49e;
 I6529b2ba884c7977f550cf3410db444d <=  I5c3b87e1908cc3d152b01573f7a87f2e;
 If14fba2b2f70d2602b88ff0e739e113e <=  I302648ef72470338675f108cfc2936b0;
 I0685af82b58f41fa65efe1125fdaabeb <=  I6e11ba6fced3ffc0d8f8003bf04bdfbf;
 I1ad44f9d9abb2121b183a93dd1af4fa5 <=  Ia73537a3f8f0321742cdd459d952f4af;
 I0f9dbc9aa169f7d63cc5789cb75c3a2d <=  I297ad7a97cf35acb5bfd1d0612044c49;
 I5e458356e7698884ee785b2d5f1c368a <=  I712af4b1f576a39d2d96aff81da4863a;
 I9b0f07f47267e3b0e0c545f44f5dd9f9 <=  I4a7d547601279634b9aaa30a51fbf741;
 I3a4dd73e8b3f48746a991573531315dd <=  Icec463cb0767bf054a74408bc41536b8;
 If727e9507d63727b0d597e9a5fee202a <=  I1ac433e960367e2ca78597357deb20a5;
 I9253bbcea2dc3a74433955d5f5aff705 <=  I7ca1e2fa8fc3e66fb6e747f2e0808e00;
 Ibbabd657d00fc10d293b680d89593ca7 <=  Id8930a77f5475a80411dfae4698cdfd8;
 I79b7daae3f9f65acd3f79d579d2af25a <=  Ifc5cdac396efc12756b713195f9fd57a;
 I74a4a1e449670380db8fbedbcf2aec04 <=  I504e5446ead186c601225c6664e047c8;
 I9f7da2708edf4c941682b24f3999b159 <=  I8d9b55049a74bde1fdf26004008679a6;
 Id5d585b0c590354af34d02ba320f80d9 <=  I155a7cee8b9f8b4d03f59ecde58fde8a;
 Idab5b4bb4ed70dfe122f645eaf32852c <=  I9cd50d02d3f7a189b5e70907ec8d1e73;
 Ic1793b6e075a12f6c1dda7e9fddc8b6e <=  I04a06a7a7af3891b0d53b95f24954344;
 I168c51768b35b16f0033808f0b915e8c <=  I21ea05b8f1be5a38bf4a4251644c370c;
 Ia7fa2fefde3f2ad6a0bee771a131219b <=  I89b558f53cd3391108aaee100bb68698;
 I22d2ffb044bf579a2cccd3fcc70dae45 <=  I0b5cdc03696628bcb061aa2113444e50;
 Ib4b3cd8d5376f6ddb653c8cf72dceabf <=  I4293b2867a22e5f63df2ee4c19c88f79;
 I2c0b6e7a1fbcd97b6b78e65bf6d61213 <=  I966aa14cea82d7fd5872c135f0bbab70;
 Ifabbe9c31875e40eb81a87f0b19134e5 <=  Id87f3e498747081eddc52a1fb671838d;
 Ic20259ce7eabae2029ca2ce312c6bfed <=  Iabb62eea1f75ca64312cbb047714b9ca;
 Icaf0213b02a3cad251718b9ff86c108b <=  Ie231dafa87260c19f1ac9c33085b94f4;
 If71ff543c013f0111318a06039267570 <=  Ief8246918e80c45898a4c38d0d5c3cbb;
 I7871649505392bea882ad24b821c953c <=  I574b308a0fd88d3f211b2acd576a3efb;
 I5c4bcb5584cd15cbbec2709f29e15f36 <=  I8b32db6febf453df9d355666241b9a80;
 I73b98efd2185919a61b91a641fd6bdd7 <=  I7066424a4d00d757a4a0af28b0d95166;
 Ic2519d8c4e9b2c6f2126407a7a39fefe <=  Ifc4d0343efb2e2f499cc6d8e37591f48;
 Ia806cdd7fbd6b44a8256aee7250ddd8b <=  I1600115eb31dadcd5e87696ca1a34fbd;
 I9badff60aa84397c6a408b846feceb91 <=  I5dce546007aab5da05bbd33b54ee3dba;
 I885c54956c3ff7dfcd971f9d7ddf2db1 <=  I6a5b90479676374b60fa668a358b852c;
 Ie3ae98a6abd28a3c39863a981e88e63f <=  Ieb0c46dc3852312024e2bf158d159f20;
 Ia1fed14f941d2ef3e78c490f81a5bd04 <=  I56080da8b243334ef8414a095477c286;
 I714c5a8ac1480b08aa2859680ae40660 <=  I661a66590947450472c1cc6b8dc9239b;
 I11d5e654536cd6b6e9b91487d76facb6 <=  Ie56fe9b766c784f90771d1335e397e99;
 I32f53cb8d864ff40c8d0ef95e9bdde54 <=  Icaa6152af5f6bed3d595d51767c9ec49;
 I0c3874311a119530873f475b01006dd4 <=  I99bddf2f101ab41147b2849d22bd8e0c;
 I585684cf3ba45f359e0f0752e9e88819 <=  I5ef97e1962a901d1e6557c0dfcae036e;
 I998f8a35c7ec923067dc75c76c9df713 <=  I3e1118befba3c769deb7bbf9d1875d00;
 I4e8f27bdc42f1e3f4024b020d5821dff <=  I435152993799746e1f967343ce1b106f;
 I93f0932897b358b6c4e3386609cffa36 <=  I9e10d71db16be96b3087a3a584a5b55b;
 I9ae8e176f8f34220d2cac97abe1fd32a <=  Ic943175727986874531ace57f5697df3;
 I7fdc9543e6c7c0324293936b1c2c8f2d <=  I18d1d32d1e58254b964c670e0d83c119;
 Ic9bc7816fcb1f128d833fde39ad8cf1d <=  I96b27127bbc15301b57d83982260853b;
 Ifd16243bd087b16c5bfa2bfbb8239ee1 <=  I12d97a28ef39f26eb4996aa2f1d9eafb;
 I3479e7931017ab45aa4e99ca34b8b5cb <=  Iddafd4529ad594eda9835e76efa116bb;
 I7cf57ee976846690c3286f08ef932683 <=  Ice9aeaff41b923556b30553d8b42da47;
 I32769b7f105065785745633dfef8a4c5 <=  I33e7dfa55b2d2ac83a8f57797fcd68db;
 I47e2d27cbd69c85106a4aa3ac2784eb0 <=  I5c3dedd601ffa33d7b649b2c08df54e6;
 Ibd0efa281371fa3b94eed5e021c73642 <=  I1660ea57c727ecd6e71a4e9c4c288b45;
 I82aaeb65a83948cd75521499d2719001 <=  I1c9e513f7524f52e24e7e80807a18ac6;
 If9854de536b8ba1392ba0328ef7cebba <=  I3d1372ff9b830f5eeb50c4e47d322cf7;
 I731416642a03748ca4698a73e094c500 <=  I69460735237cd5bd0f26254f6f32e357;
 I23c90590a514d430c9828af570ebf16a <=  Iac63249f3101e957234cb4efee5f6771;
 I2d07aa91cf23a7789428c96e4f73109e <=  I769cf83f4404ee0d85e6c13b7d0c737b;
 I89fc8a2a491dcc20f2556e7042d22384 <=  Ieff66b38feb970b4ab3006fb31e5cce3;
 I0f76a71ea70551bbf89f01a689811954 <=  Ifbef84b3392347c7e0e52e232d26f9bd;
 I0b6ce8e59afb2e48df79fefd5450971e <=  I13989f78ab3eab13b7f0619fb0386e3d;
 I35a8c09862db36ffde26d27b74baa8ba <=  I61af8fbc53b6f763a8b77012fb56be23;
 I920593851f5860485fd105f8d4c1b8c9 <=  Id0969f699976b1041d15d62912a04b5f;
 I51dcc6894ba28567c3077ea409871161 <=  I3be47f6dae15615b1b6b0cb52bb8cd5a;
 I79489994f40f88e0b5a8a8be6322f3ec <=  Iabe728226ae671218667d92139083a4c;
 I6503341e5d6ced0d71bd29bbc622020b <=  I49d60f1269fcc5a98196ac391823ca1a;
 I178d103fabf53395ce88cdbfc14917ce <=  Ic88cdb92bf89df187d801b480c7c2770;
 I3a8d57af0e6ed1437d572534742a9f2f <=  I60a972d5f2465dd5f9c3665eee4cffc2;
 I4602a0caf02e37e360e5cf9de1003cd2 <=  Iaafcf98c2c079884e32f2bd70972e5b3;
 I245a6df9f9d730338cd52169a3f466d3 <=  I3c4a90a70e7cfe814427262cae88e2a6;
 Ia7a8ebe681523a490c83dcb84ac82a2a <=  I7eb2363c8fe8f49f839b59df19165aab;
 I7caf04f8880b455d92307bf521540c38 <=  I60bf9f27a86ec731795d79b656e2229c;
 I401eb53331986f8474c861acb2b2a445 <=  I8d4fa08cc0155e81bb2ce4ab9a39df4a;
 If3e4f18a03ca4b7b1d89ef842c68e96d <=  Ie21b4ae619493ef57536508645aa29bb;
 I0d6bc03eddef33a7d70ac2cc27049107 <=  I854fac49e7921a59773ab612181b9569;
 I2214bdaf7568fd3c20109ead1daf861d <=  I20a9b10f04d9eeca6058889d5c930294;
 I6138bf9b2a35f3b08f216eeaf3c0ebee <=  I122fde74534a82953b1a5a476e2e8151;
 Ibd3927f27dbf4a60128f60f31b5a32e6 <=  Ia535aa71b5100fd37cb15ba1612d2d52;
 I26faa75fc5dd15baf23481311b220832 <=  I8b588d7b4605f968fd007ed894b4ee68;
 I373328eb3cc59c5d3d7a5102535c5410 <=  I88d97aa0544a09e2a0df10ec0a57ea54;
 I1bb3c77cdfd0b229bbdf7b33fd4a613c <=  I81cb66f14210612d88911543c3517731;
 Ia1c8178574520829f24c8cc08e15e8f1 <=  Ibd10299291ec40ff247b816be64f07ec;
 Ib911176056f3c0378dfa8a77e0c5b69a <=  I3e4ecb5c8164f70ca4b16eb004cb276c;
 If9afa8946804ce9c74ef43d3ca669849 <=  Id5e6fca7b1cebfd4f2caf7465fb678fa;
 I6bb576223350a8373e430d185efe7fd9 <=  I58a570689c10954778a3e3ded8d4f9b4;
 Id7008a8f0d70f1e23a073745ed4a57c0 <=  I0a8dea5e3f82d6954d294cf3c3c858d2;
 I87e0bcba46bcc28ad02b7e0af773d82a <=  I9aea2a89a8d17d14da2fccad570cfc7d;
 I3bb6f388db8c8dc2b6c963749ef48096 <=  I8b661503122504ce012fe534dad9c394;
 Iea2bbf25e38901d15434dfc83d65ada4 <=  Ib9a8e5b5096d6c5ed5cc315a5899b8d5;
 Ie5e331564633cd16934cd0714b2953cb <=  Iebf5cd787ff1d73dfbe4e52cfbaffc14;
 Ibcc6c8744ee9a2ad9766c0f9fa196036 <=  I4096de17c18f5e0af8d288bc6887c6cb;
 Ic425c518a69f3f85e219b1f15baa5d36 <=  I949e53f68343283236a519295c606cc2;
 I78ba7a5627868f3c0b75555131470aa4 <=  Id9fc0dbdd3cd0709ef28238589312443;
 I3b5bd630c8d2bdb455b6f75a6a8a4a53 <=  Idf5ff15e65f46f3b569ef0d634cd5819;
 I4274a587dd459b29ecee1ff1554a12f7 <=  I3d70051f81db3db896a8455dda9f0022;
 I9728cc3e93018b67d2c2e94f9d90f433 <=  I737715c7b75b324dca40210b708166ac;
 If77d0921ff0a38d2b3fcd28c5be4a131 <=  I3deb95e95d3308de220901f8fe6d2ee4;
 I29046786efe54344e3cffb3e5e913667 <=  I5e7775e3bc484bed7a57f04b0cd7ccca;
 I6fbdabe9ecefa8648c4ca4ec51e251a4 <=  Ic557aa69aa946711cc39627fe6133f87;
 Ia456c9d3e431416da7685ea0c42371f9 <=  I004142a2c8e12e72c3ac4a439b281fcc;
 Ib68b82bab62a694692b3fd2191b5f29c <=  Ia112b4cab1631793a8cc6291027c616c;
 Iacfc43c384ab56bf924d5ae09a59fb17 <=  I3d3a0cda05e77a00523ea3f4aae38d82;
 Id5c5e697446d9974b383880138f73778 <=  I723f34fa0b35af4e77fbecc65d2ca88b;
 I441c5f07ae7d849600f2d02cc5753d5a <=  I460bbb250271f3fa5414de2e68474fbc;
 Ic117c98ae21f7640aa5a68539ec03821 <=  I1e29e4b5d18509694df3a0e7b7cd2a7d;
 I4c3f1b807cae7d5a4a5dcd3c8180c0fe <=  Ie25c961fe6b06030e848c7b9eb751909;
 Idc31f916f132a0c203eb03a7d1de62bb <=  I16c56d8b22dd23fbb09ebf4f36107cc9;
 I68ae757abeedcaee5336b7d45a29b8c7 <=  I1e10a4b5844d25334b74e1088e2d3deb;
 I5e4276800e079f48c3953f01869bcfa0 <=  Ic524b9ac09a3499b67313edee303c53f;
 I30254925c90cc28a13afa22e983854bb <=  Ie332a236ba72fed22c9d7670390dc3d1;
 I5955344e0f04e1ddf15eecf2eede2346 <=  Ia04ae82f80fd35c0eb30fd17ec9f74a2;
 I82b8db69079237f10477ebd39a13bc16 <=  I009b2657f941367412da0645c61a6161;
 I83df9b9b4dc9b0eeaf05f25e513d1603 <=  If84fc94571af2905f59753301bfb7fec;
 I54e2da03e41cfdd43ca24929ef467819 <=  I782050339f5fcecb44819e7cb6dac5d6;
 I5b3e2ec3e81cfbb4cff4a55faf1779ce <=  I5ce602af9806ed123e70480c643be643;
 Ib5d40f3069e5a3e1da68013a7f5e640d <=  Id2450e8bc8cad7c46f1d47372a344f12;
 Iecc3e2589b1a21ad89360386cbc59203 <=  Id074a700da35c1548c27b5d1c7e9eea0;
 Ia4d367afebe196ee6debdda4251771b6 <=  I689e819fcdc296cb4b537538012615f6;
 Ibce5b55e9f3477e8cac134660f3e056d <=  Ic2824f1963f1158e7ad33e9c81bc7d08;
 I5f2c9622ecb56c3385f986e11cda6344 <=  Id0ae33a482904b109068ad943d76d758;
 Ic95be5fcb699a68e0e796dc0408fd5f3 <=  I7b7386e46768f03c912485c3c80065dc;
 I01c4e6856aaa370540e370d30223a3e9 <=  Ib0e71935bab4a9ebf00d9b2d170b571a;
 I693343088a46766b65b21833e8c93424 <=  I4613dca4c7c67e9dffb22110f62d93a1;
 I363bfe5c6d747f1b0bf3b3795973cc1a <=  Ifc0a83912f31329972ce02109fe40df0;
 Ibcd20a65390727b99272e778f6b5cd48 <=  I021270a1b11bc14783313a27684e1a08;
 I824e45de28b3352d3189623ca276ceb4 <=  I0f8f6a239a05dba04dd3b845c9e8ac9b;
 Iee99e323224f79b59ff094ca4e0b730f <=  I99d616bf2017cd8e4f019fa9356a4c9f;
 Id6c903e77c0ae87fc00b0a19926eac0d <=  I48c538d54789fc85a7349065dc33b20d;
 Icf2d8147505a677d965332527efd32e5 <=  Idf3ebc5f6ef593255d94f70583e028ba;
 I10edceddaabd0b5704cfe32642099bfc <=  I5ec053664237ddc305a831b20239a5b3;
 I7af4f3f04f52198149fab343b09a7c33 <=  I2150bffc35644044c52346accf50c6a6;
 I5b772125b565150758a1dd9173661a69 <=  I9a16fe81b2e09494fb280b564b2d8447;
 I8d3688317aaf1a973e53e7d82c07aff5 <=  I3a78158e0bcd94e117696bd698f00e43;
 Id1bd6b209ebbc1dc87ef765e8311d13d <=  Ia674fb4751c28067672ed365648d4046;
 I2145db99a9f07a8dcca7bb21537c3c6b <=  I7c2f789de92dcd3106cd534d547ff653;
 I0578f5f40c3743a4c0184768a6842378 <=  I42484fc96375ed4f28054b45a7a573a4;
 Ia36d890f9c568613260b96683ad1442e <=  Ife0e6d58f356f10d7f769f225de5a7cc;
 Idd923fa51da8d881654d1a0b2939bf45 <=  Id958719d49aab2d0b082a6d24fe4c3ed;
 I83e8203369eabb1165454d054fc6368a <=  I6f030649ec413f3a8b1b2818f11fdeb9;
 I811bb1c2a735a7b3b494db92a6e09bc1 <=  I1b4cbdf5cfa3d8c53d2000918dab9d92;
 I2cf7c8df11a71a3952a5c11fce1ab746 <=  Id48425985a33f1512c0dd32361ceb85e;
 Ic219b4e5b38cf27b7c30f1b1455db7c1 <=  I37d45d42016be2e2bc96ae6fd4287f97;
 I964950b31cf4117e79e46a2282faf273 <=  I6715c7f4ac584103721a33ead7ed395b;
 Ic4ddd59bdd32e1c8481e7d39707d2628 <=  Ia8e9d2fd6a51de4383c16a35737a1831;
 I754ed93d8e7f3ed1b9bbf1aa0a780631 <=  I3efa217d3d93a9a2f15bdcd906a2a230;
 Ieb469f605aef6bb6cc19088b0a8d191e <=  I016707bf26cc19976929a8b14f535455;
 I0be6033ae52cefc976cf28e9c6972b2c <=  I698072a5328a85b0b22ec7bc94b8372e;
 I913ad4107114014e726ae5a684208f1f <=  I70a428ae2a62212ed93be37b860e8231;
 I332be99f2c509a0ad9ce2003f3894900 <=  I5193a317b4c9d2bf1992ca5cf9936681;
 If615b5edf5772640f5e7db1b7c2b827e <=  I9cb0c1a404a77903890379f0f658c70a;
 Ic98c3c04426af7540b59e85693f8c85e <=  I861bb6fa26ecdc43776d01811abe7bc3;
 Ia8b37c51a90549caefe7c587af95efcf <=  I92ad6f4d3a62fbd3e86cda7457115093;
 Ie34547c669ac94c6b215f01c235086e4 <=  I17f6c0345023a3824d5e40506e4c1919;
 Ibed1e35fd09ac08952020a915b52aae9 <=  Ic309d272e0e79647de87c07aae1e798c;
 I27def56001fb56e6a85c9c61ba8d55bd <=  I24a4c216e917b9b9ad744c7bfa4a7d24;
 I6540e74c5f9178782a17fe7460aaf4ee <=  I7112d906a2a8245dd62b7ef26d7e54ee;
 Icf92b5275d264e1b6d832272a0d01a66 <=  I2590acd159fd90fe367126ce432e39e8;
end
