 reg  ['h7f:0] [$clog2('h7000+1)-1:0] I111cd97f7c5c13e18b528ffe1d1a871f ;
